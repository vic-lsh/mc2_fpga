// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
xFgZOM9lLzP+r/egZDQV9jTcfvonTybJi03wHXdtY8faXiGEXU1iCwlBxrNx
oAOMyzP/b7/S4OiUspIcxEI9VHmJPBuav/Ch2n3Ze2lYdPhTQeiUV4tBGniz
wPUElO/Jl4CJmox1vgCp1nwjvCulxtGpMbwjPBpknv6EXN0Gqa9UU0hlcnX/
BInwEITPoANCmmzaE0Jb65cY5SkE8caNRnaMyotKfmIdEblmcWav8TcdIVZc
2JA0IMl+nV55CqNW/DbjQDccvlS7jLnPjjlM621IoPcJgMybVOxEDqWDr++E
EIsc45TomFjHZjydlhOOKOnENrmxvYf/80zbBVOTJw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HJjhaowhQD+tPKdvq0pbK/mcXPRWzNB+II0IsQSa35/2vffUWFxve2jEtuz0
4++cZZyJknO3ra3HaNX1ppzdoTD5uDmFsNvpB+j65NxMhdmVzxu0Bf5faH40
AIURJqutB+60z0vL8y+nYP3TtfGAlBQgGu1lrEnTVEhLZVYPegqBFHevafzq
VKgT9jgFkFjM/et1j2nzrKqMV/Nxp2lTc4UpNNtLGL1XepKK7e13Zc5YvENX
J4zbEQsOT8T4I8iSLfG2X9G+CpEHmJLdt4BugEc95yraO4xfGqSqXXRmKzuC
kjbU+hzZWf2yjwZlvNXFIA+GUhzdQvv2QyK7BkAMnA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
O47jJ6SRYzUIrgc/cT17iZiWnwMC+bbKkjf77ZzYyLwZFlIR7f3F82/6fANZ
mdQNuzTnRkTj8ZjBxdV8PCpYz7iLX2x6zvZgci5jkTgAGFezha2xICg0Fnzj
7wzoTc65Wobuv7S1vza0xLHzpef4Mdu2F9c+QPaEAKeTCLvaL/nShvSviFSF
6v0xyB2AMPQc1VDDkwnW1L8eAuxrTak4ZAh2meioYqjrQJcytfb0kp3YcvKs
irSdx77CPSRr04NkDh8AIyqRNoMCk4FGIl4SRtOOitH96fvbEGRFDD0+s4nk
7AF6Hd1kUEyERQsMQLpLZs6CxBm2bwtfzFGBeqkN/g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
A4KV+VsOs3DlgLU/4fQQGj2wXyhSXkg4zau5IguRKNdkVVflx7nKb6epZt3C
y4DT/DIHS2eRzkgwTkWHpuD9oWI/QcfwaDmR+ZPlLDOhqBd+8u4J4KgpAy+Z
psHpLoBbvDtA1RXtlFwJ2lArn4AmCPaHHj8IFVpjHgH8iVddNzwZW9zRmv8S
8EBs2FJETRawtqLyRQ1BxBYJsvjdpYXq/gUkNFl2Gt+vSpDMmyqPz00CuKZZ
wUEWbfiU2L9aKP/OrE4vHnJ6VoqxyPPHTyEEECkAH877Tp7ytym5d7JeWuky
9paw+lMsC0ACj97fGQ0Dl5dj+Nah7YAuWzqZriS8lA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lc2aORHesmIbL6iHX6pe2cH0c4ndEI5hNzsY3N8o5ybw7rpKuiUK8YssfRwO
pLyFG/JlcSTgdOLhmrPvJ7/g2QIwqBg25ScgSLvbDFEPCNjDzmxEstl25tOt
U2X5OgrDIuIXYqDfDXD2+/UpfXtbD59OC18FAwOJq8Oe86Zd3FQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
bP2abv8xcI0sD41i1UUmzlF6up5A1MoeRwtBROcX6fmeDmW5SXdQDOexZmVC
4Qm5FtBoosGoQZyVWkgtUhxkblHA8Nspv43PptB7RawgmSiVloC3q6XQUMis
affpfoV9om18tDuJVcENm6rhZNVTsWB9TgGB6y976x9EWn1NPCW082cG3w91
kJrUc8qd1sHJhBlLFLegkb6w1tyZHcVMtgH6khBbNQJS/AicQWF5QZXXUQDH
EeyD4vlRtg7kM9KouCyUMFE+5PQXxL8PX1s+1v3rzqfYYUBH9X1CX3uxJIQ0
/EcLTVTspd2AsJhiaWmF0BE3vlV06zLjTVhkMjVvEx7x0BrAMHjubTBSxDlI
Grsk7EdGIw++ZAbtaUwUGLWjkF+KG/7LPqVJ+gLasozVgvHBACkwOjBVU4PH
P2D8L6FpFXe0sELAq0qRAEpIH/cTwuNIojCepauAneIvHJoHns4bhvGs8yqK
wkRZp7wX95KpvmzcpTelzSlKluYWGnfM


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KLvG2jePSPhdl9OtY9IAa/GAFSU9Z9d4s3U9GFm/EEfM06qbahbq1WNItbrT
3osj92Yt1BdmECzjEiPbGRiccmbwRF13o71AtnAejQHqUeSpsSuwLc3nRcvU
Stc6U0+A/odZVYqEjl1o1DQbvspJ7W6ZukoZv8NshpYE/CyxNVw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
H0jlqCZ3M2kz9RfjyIu6euUXMcFHeWXwFircsG5LBR6dfN9HqoG9WCi72sYB
y3Hpn6FWq4hCjptGUq1s4yGEVaDg07CiPPwP6r+29CvXDsJoL7wMXEjtZZ+b
9bpHOV56y+dBizUgxebqcY2+CWBGlWSFH7Auyfufp8QWsZmIcXA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 38912)
`pragma protect data_block
AWR3ny/r0yPQEymonPvKY1pQHYPZkOFnAtw8B2ny05JaNGQANbAbnAngiaD5
wFau8vG0NHBmY3B0aMu8zOY6H+3uv3r1vyyzH7dwDbAlxeX4NE6QDMhznrI+
3hnvoPKCKb3AU7697KwDK9050RAoXpHq8FhLz327n2td7wMQ9K2iV/Z5iqqv
iBSvubtkpkcO82h5QXxMX8j5NaMxdYVF1dISS4suSyNglyb2Vcv0WmDobmIb
lAdD+uFjk5KA+e9Q98q/CzXCX1HU1VqaLbNmS1Tze+JfwnMjqJ8oHmPE5dIE
V1bffXmTn49LVypy2aTDw6Y4RkXtWPqXbW3PNgt0D3raYTTNwZesfoUoAjTs
kGIRTzfSF+AbupYgReLh21TKIFJRgY9Lg+iy60i43boKzCWjys5nQz9phW+U
aFlTBb8ouOpQEOKzfCLtTP4im8pZ5op3RfiOROqxnJNroGao82vs+7Zs1w6j
taYRW4aK0hQolnshrl9+i8tTlBqserJ9kLWO1UvwexMykxT6FM6vJDRhoQqE
cwfSHz01Ah/+F7a6tCp3BubRR7lx8IR4mA2vcVgpTBkgGWkS7Mpzfk8WAQUw
XB5U07AO+Lz9jMWXdFQJmD7an/AyX4bLs7twbtOEjPc5hkx9QZeR24BAkZF1
mO7DHAwcMLgJp4ZSOqULju8yQAf4cEppPiaWUqKhtAw3VyWZUCXUfyIVtiAV
+SosCE+oeKAlEGS3DrJ0wiySJNIPC9uIBt8BOFZjr/zobCOJPGmKnOOl8Gch
E4mVK+hISXVSBM/SgQih4O+CMY1kSsiSArBtUE4+mPT46m1fj2w6QBtP+s3a
rJgkYMyZjAKSKg8gEx2NR2kz6Up4Z2wVmaCR7RpnU13wLjhO48CracAL6xgA
2TpOZoYKBF8RZwuI4rK53SwfFvxqN0+rnTt7tFRTcvdF85DEhjp05/48zGGf
kq61Zq7sXxKF3rB0Ler0v4KUAfyIBESFeb6wNvl0IoDawjenyZ1dJT1SAfMQ
/N2pQ+Gjs8Xu7ghbFJdL6uSA1nCnoas3N/W8Pf34M+KBBl00HibbH6ojWb+O
jWM8mEj7zSx8iAvf9LF6jKrXu+k3Zc5ZLxWnPVAQXpp+j+Xnv5HfH+qq62sL
1n03TJjdkN6uTBjLNbsxfuRGStBhw05pFoE34HSrtL/L7o0+z+++87j4VRIB
fyLmi4J2pKPrXo4G9usCU79r4M/NrsuHHZVARvpeFVe1twUG5nOFSwXXLbIR
fH71h9oCWlo5ur63tnw8qINmHy991UYGjsxAWxXOS7KhHALypkK12VXnKOw2
o7C7KLpcA/eiee2mg41sr3nskYkHpHD8AQW1Gu7TY6WsdoYccjUggUbeAgZV
tu+JnMB12W8zAYOxI6d99VXLNTX0HFOctiGqcREWS9U6QYHIrDwV3Jyg6zPY
NXgty3zVP2LS9itnjmJrbMCGzVG5bs375Dst8AYZpbhMpbeh9F75xZVy87AC
vuCuZnwRD1TetBqJlkmRkF9PeS5EJaTHkhsEHspyavfQVTO3Vs49i3+9OMbJ
JI5FANm+34m87+cQg2gudJE8jn0qZ+Xb2tD0H6H81is6IjwboljJ3lpkGbrn
W7OVKU1YqUVyFtoYC2Zg29LrtZD5zZuodQJiYOAtcQAO0NzIE6LDSC4Aht6k
Ht4jKPAnOH8p+P4HTnWsIlLrP4oS6+9PeELo5moZiNzjA6LpFCpBWY9A4/3h
1Pk73tRsofOSznrRFAn4bcaUwJplrT4hVdAzDFrPXpSmwrW+6+su3q3DhUzB
tJgMb4c66C8NPwqF9v+8dfWgGGToReocRDYAwzmjbz4TrUkW0YUvIqC5hWNn
6pQZGLKAZmeNaHgPF45CdntT5FTfapGnAXrBKkcD8C65SxiyTmEcplPg4GxC
RbI36rBa1XVayKaN4oGRxsq0826f/HeFJJrgP4+gx0DQlJ0VcekGxt1pwXIO
Indnc7NFX2yTyhuwetgys/0zstC5pX3Ccv3MO4R6P3lBHb2eiDW3XBX8tBch
k7YRKIHyoYLPRHba5SNrlFufz535vpccZl37vqkX9pbRKcZ6/6uiAV3DUkJf
l+BKNh2e9Z2ZjWvBlullgx9Di7rFhzZpjMmv7O2GNOqMsQ9uhqLS8Ke2gMWl
32FQ3EZ1NE63fzJIY0qdGuPelQSOUHnvevvXq9L/ZfwiBWPTDcQeWI3yYgPm
zFsIHKyAshZjfTQIN0o5MR89R+xilr3JrLjFEwYEo6wmrzURyzUBU0F10WMl
l+bOcj7OAU+NNKYKYr/ieTe6QlFErLzyqcZ02VTmk7iO2ZWajE3fYNvRJXgN
KE2tgfCFiSDIIs0iuhAEtOm8vuQVmrWMbmtBabOg72G/FDkTUnL8UnVoDmaS
kb/3XwhK7ADFIpVUpXybnVSj5VtdBZvhJv5vR9ze1YmCBabwq0gld73g0als
LEPv/Z/OSj6IIFdr3xodFrRbj12fQrgyoptpUiAN7Kp00p03JKnigYqhJxPy
S3bQH6xRSHmm71hEyekxmfNKRNtt9dv/M2niVRqS/PRzC3qjAfmXF1lblwnI
rkDjl9oLlLkL4ML9ZUQB0Aex6xeC1vUzyoqw9TnBKL5Qd0FtPiXgDZT8oe6W
+pSraI+ycsPHYLoR6gMgBSAeA+DZ19iPpLlr2qr0t5sOBIRCTHF8jL/LXPsV
u+Br9Qr68yrgkorI7VWkw7/3qDYw/KULCeFldtRHjKJJ1Wi3l0hmF3wjmBjG
VKUrPRKlmcohwOB/7D5v1OnlmTNdl8miLszd2OOmSdlA7cW4aMIdbkMn89Cw
w1F1n/ATp4IFXQRWJxjS2JlPri7CUWrU4Ibk5mK0g5PaUaRCPSYQatRdWaOO
3tLn0Yr0Km5uoknssCTcZKSfaC1vdo8i5JK8yqYM32ZEQW+cjcsERxW+dDu7
v9yMXBCXDHAnSGNr2pm5xud668sibjyTvY3HpWJCwiTpaakZhofyEBgtnEfG
WA26vcprkX+fGVdcJx7j/wNJxk44G13WJEdt2mRYxcCFPpbxN2Y3z+rQjT8/
aehcmLiXqEcmobiWZ3vSMqOEHBHtMZfh/OCept4Jdgpfr586H+5eA9nx92mz
XDWRs2aN9WJ36LxnS13JKihVepOdIVqslJMFN3xOEz5/SdyKVU6uS2zcQ9UZ
8D1VGIrk3PZ3kD3Bz7/JV51Q/ZggMEIiqTfLyG/5bPKRTD4GNN9jlItp6Jc3
udgWkyGFzoPWhbgy4FsmtNZCAaWaM4bwxK/kxfoIxF3TkdugqJz2wgRgU8l4
dOm2hmkqZ6wRTJgRrZTmFStdMgIeDA7hAqUgM7ui69nyEs7bwit9aQp7HrF3
LyYsPo23WPou8sl4woOPt6pzuU/ByCHlsP9gWLCuPI+xzjj/793QZS5kWgLZ
ABgBvcsaq5e4DWBQdwJ5g7tTxLjdbmCAF/jSU/2JofmoHWAOiF8/Pd17TUia
hK7WgiDk3GPU4X3rqrt0ZydJPLR9o3hWNkcsIt3hNM/SlgyB1ePb6a8qy4fl
uOSJqgZp4kdZx7kTwXyfxfjolz03sa95uP5/mtgaMCvjdtbNMkGTLoab/DVJ
075VoYdKvJz3chCELEq3kwe894r/fqUJuodpx9VhVd6VMgag20jSISL03rgO
eOUqr9Jy4FBD6OXFMOb2D+vSXzINlLUOtVljk0dv/NSs06mcbGB4EbRWVwaZ
qLP2Bu1rAKDPeFaSCHhN3nAZhxdRuwy/fyBeb+M7GKEnbzULqyUVfp40rOQr
mDCjexB3yYbczqtBTBTY4hIvceP3qbIn81M6F8TXaivLE1ejTW/wnPdm78z8
Ujz5ZNqPNFl67AGbNVK1f8RazOXtRasW/9MNAKrmNVPakSww79uZtozdRVAu
pJBkUeanOMA00Kzw8r+lgAFyhbbZnyCVtnYbwl7lFwRQp9TC/Av0uWdsFL26
OPWs/17MdoVJugtiwalyc3YrzbDWLLli21Yq12v3F75ZsYLKY2LAoo+zvSfH
qXPcKVYCogP4+A1DV4b85IJ+yCNnhu9cSU7ZMKgqUAq7kxK4hPCZJY6cZm+F
HPR5owVozd0QuX3NxycfRuA1MUNQvc21TbER56gXEoclxVi4oPLsiXMrD2bZ
qMZFPzk29/SllZdjSSnXP1iMTk5whs5Gz/dbvFpmN0G9JDl5y8f/p9yag1Eh
hG0Xbx6v5BtXyyGYsoG0J26C4p1rxVfKm1Qo1rSZWUukB3ySIY2vpqyGcwK4
gaVMH1607BiqbiyrHcLDbsaRRIOTvlCeL8/VhnfdXGUf0kUA/ThljHD17B8e
LnpA/6vD+nUMymmaK2Y9p9c8FQaAqGx47ySVtDJdQpzrEUVIkpOw0YZKE6Z5
2GRrv0oaXzHkYjSrIg/YuAoIJZzebX0CYF0ilqwYd2IrX5SiclpHDDpXG0Mj
vyIf05sIiCf9GXy2BzVHNqnblych443MppbLy+TFOW2pFX+a3FLG2ghJJ3NM
pvSsv/0hDJ7juBwo+unf+Fot7ld1hztRnZYVyRok9ehk98ycj632EYhD56k1
YFeT7lULXJ29blbQkE581b0e4/K1la8NiuvtsnFHXdS/ZY5udZEW/C+HwK0I
+oBdbMZx9hyWWk7aFELUp0hTjIdcoSo97pXFYpO1SodsDmIi1XTZHIaMOTt5
gc3r7DnZbGXxrfa4633MT73yPOQ1YalGessZTWDjPoW3Eblc1CZ9Q7mYnUpq
GDk701rdxXmW7pGhukHbuo2EnpV0LTyNMt37/b0Io6clWulad1s0cv5DkAYf
NWkKQgNKXJF5SGfh9ZF7O91PetAmx/N6RsSWsFAoaymoWit0IoTSrfiAifJp
v3leSMqlC4YCXSU6Zbx+IoP/3gHcC4a1wa5i1EpI4IlYteRwjygzwn7fOGMk
F97DzD283qfArZG+TWuI1ShaSp/R1RnPi1xqzJl+mDTKTiUysaJMsgntGocW
HOCDG2uewB/f15P8ywzXM7bYx7C3TQrgfASAurNOnqVS5WcEj1g10R1F4XED
FFU9z+T5IuCCC7ykTUIttKrM0m7NtBAh2ywQFOfjJV4wCOdM4otJ5B+VD4wH
FiXkpd9Bx34cVLpAWsWfFEex/0UdGPW+Wo4GzwYEvx15vsNxB2pvXkozhdHy
fgBMABdbZW2K7eQ2P7C1zoPmCx1WkiAKp93oI/1gsgE0EJRdevl4uCsZheD3
aVkx74oog+tEzHQc2GYhCilmbCGe+xhCvIyRWzOJ5QEkh7dn1/8+FbZI/ABU
LgKsxo9bE89KgUaJElu8pFVZuVrvP0xzMuWy9wDQzrupU7BhZb18ZV/ySY2F
au038PBdnCsnjrOjnDxhM48txho84J9ErqqVOTv3dzS3wH1yHJTLnX6upLjo
0+xRPS+yk26WIbg2vVQPKz7eKzqn49chLzLDEwGZ0QP09mU2dkXCmOZcpB3c
h6hquCr8Zr8PMst9PVzg6JTRN6dLGPwwfy7dHsMsIjue3Y8LzGQXt3qiUTtE
y50N5Rmt6BZu1NjtahYo5WSwqmGwm+km9o1e7D92w45KlJa2rtl+cUgnxp1Y
CBWwntAvavtpXZAmbCjb7p9rBl9rQUI5roRBokZwuoHieMtszL1+xTIaMiVD
944EddEgUg60jkags2KV4MPctnjAQTY37/CtV/eVBWG77vun/UBCYRpUKaku
k//QXi4VxvOKyAa1yvevt3GPBGbKA0N2obfSZ9q8g7bwduQeKCtRjaswfc1y
WS7LPgGmSKR+1cVBrC0zuK3TWsQVIom3hVQFi3zZCEHEeW8fi2HubfjWnc5m
4NDRv+1ybftr3SJvOP8HnPaUgnwlg8u4zPKufT07PMZzI2h4WUzy0LvbkoGb
aWf2GF1wVXwFhHo8ykt5Qt02Tavx7w9QnflrK78o7ODjDC3nXISiwTiUBkRl
iGKCnteBvF1PALnI4xArWfYFLpseb95anUO7lwX7B47BQtJrtuRS018qqwnb
7oK0/dB287i+v156NPC/YZiV8dMe4D52oJvuri8GL0bu8IXcsDSDO4R0dH9g
yBf6DWXhVBS6IkUB8X3MyD3N2xQdHuxdN0lYsyJn8jrdq+qFBMZI8iXmPN5C
/TgqP0tQK+ULRcEnUuWAk6DnKks1m5sjbwJSCJCnf+Nk/uPQxArCSu5CYtkF
6pr0jomTrduMIDVwO00nl04T1L+ZqpNAktLDWufvvMMUG+wjqpORLa0h16dc
COLg54sk111OVCuqchvDh5ruUN0+i0JIxOU/cfnGLgDSXScLd28O2qRfETJf
Q6u+oAUgkHnDoogTMPX8BTHT0B7LJ80p3XPIZM+/9Lq6SCubZ59N6gWLy/UC
Go4+voeti4i1yikeHoTbijViOHixiits0znq7DplabqYVwTH6OgsT/Hxzj1b
Pwz6DTwq8tPiVshz3dGzsseFO8keh9J8FEyO0ZXkjKcXzkjwwgsOlbmHVHe4
joaN0onOi1bXFODfpGCiYMbNo9OXAwmCsc7XRu7OXcAM+GEw7htRBrbnT65Q
k8Ins8BWPXBpRkLlmBaQi8xs/7xB5YqQ635Fuvh5fz0P86umLm6nyKKzgFJj
lFM+jpR9VjiPMz86zB2bKUjRxo2zAVqWHtlYT/cu8G/L6Lbqt6TMcDfYSJri
MffZWo4EqD0fTvrDp1OKSJaAXLPFTsQR4inf/BreECdeGYe1BgRS9fnO8Kr2
lvAjztxQF7wO0jxBZ31ROaJuUv9VKPZXSt/Sbc7rIzQZmPg3yt6YJUC01jaE
6AezSz9kkoH2ZrMNxOce06TpUrn0ElyTK4f9wRjZFh4zVXwUu4NcDAYqkEwa
y/qK98k9NjrR6dWq/mz1rIR6GrDixEVFYhjtsrZi/IwDRG2XGPvTassouhSI
mAL32K0K3/xQNBOE7wrf9SPWKqjap1AiNd/r0VZKS6IoFVLitSvF01jOduep
SKXZ5z6adI90i8itRQTHiQ9WFfJfr4z+KxfUWV46J40UUoz4imFdtcbF/NmB
Uwv0eXtDxRtIyRg1Pwj3RCd3pc1Dvcuhh79UDLOTWsAagzB/hflI3HrIoacV
/Qc4QsmhbirzYF4X6KkIKX75eiHrQw3UC4moBzwVgQQvA0Rt8W8Tfdk5wz/H
meXSQUTeNFYeiOq0Ie0Sm6mhzn9JE9GJC/k3KsniMA4lznKXRpr1HVupNBCd
jquYRvgINXRej1umyl9tcJFnhtiWWqVSnPE0Gs/J9pOZ/HUWxTXfWhp+bJ7d
gWp1J7OGVSaLH2+j1OUWewsrGMRI3ipxxrvOaNdtEe9XbC6SHYSUEKDq6jzk
kwtdCauvM+EYpXMcPg+yDzH2CQqMlamDR82ttlMEUUYWoKGQ1UDGpAtaawuF
MhOZDJjiZkd182vuzM2Xo7W60H4uYoEK1P4eKNI/ZQNydcFtVGBkvLYHk0pe
XXfC0sZyHciTx7TLctjc8siTwh3kZDY3GSQMXeenXwjCNPX2MvjxnJC+5WLL
jNWgMRM3REXnm5elnsaznBbd+Wi3WOn6tyjduPwS9GGc1aJJ5JoJON5u+0kz
EHs055/q9z2GAaq+4GeYXOVpINzxmAQWr111oIMQsHzk7wW4QIEUz9LkZteK
Eav80pXl/JZro2v05liSkv4J/2wm6fZXTis03YJOBs8onxtkam8+GEwZevbH
Nb9DZ2iHECqGWK3nztwNfwvPIooxZJd0A4cJuSmrShBa4mIJcVGNOj0TMrfN
OTYbia/gGFhFw+tPdKHFiegPtPsv4OcfPFfmz1kOY0sTDnDN1D8BuXteZaT7
WtyNs60ytHLy/mjbwBAZsjfm/AD/+MlZVKlfpT4C2PV0ACPP+41aTA3HMJZ/
prOu9Zymb5vv5HbLE96to6CUmQaDkMx6PWqWvOf+MTf2zr0D5fGUirSS0b4X
Cf8AOE1pcLlstwwNFjR5TLTuISeEESin8+eHbwLnL21F5g82ZqEsH/sVTKqB
FUFlnmiJE6+UfCbzidYDyBiwHG7kXmGo8LTMmntXkXlN7gRjKhqSKg3EhtSh
2lPXc0xkop+AnxKgoLn1neyITpAz4N6Q5DNUL1a9s+ASSpgeMERZF75a4MpY
j8zYUFbdJQZH6iaEnrHOxzYQ63hb9MN22IoRxtrm8JWILdk9+a0HB6l/XQT5
OAhiAY7K7CL8auRCV8kldR+0+j9pDnsJ4zAdJeaWW1GzZkDRweI7p9a4zhre
otq1xePGHe9BOcm5c2h+omFWUIckDRy/x2ofFRZ8CXbv1FINZ/1B2ZHw/sge
nmjTHeFXhkRi6j+WdMyDURAHqHvBvNx/+KXMk47b9OISiIo5k0cvjcTUVhqN
RQC3+AOOl2Z2tzXVyvhebLWzanUWMhRYtdNrEtWZhmmhTitavEXWFQlcNNua
K38GPu6VaLxQMemUClzV5G5RiSUON6bLR1262nm2KGJvbzWXCQo5M7GHqSaz
aJvwMujMrcdrcJX+eVIj25Mts5aRsHj9EfSsRlpxb0RotaK4H3ypIILZh+sX
QK9JZ6sYSRqnnqsjEPEcatOSLH1MvSXPDumVFxksT6e03mb7WWxEtRuHAm09
1uMZ1XOUZNwT0oxJJy40AYQJCp1WmJFC5vp5X1eE/CsIJKStjAKpnbwJItX2
T2mFW4NlECabYvpgIWk74Edokm8aXp+HHHVO9UtI33kieSJbZnoHa3z1LABD
Kj9CPmxJYC2JqAzGSFCKweEdj3IWFf5MswHWGcN1eoGj+Qnmm0g8sm+Pa2A1
LfVSulx7o8m9n3Ki6a+ZcpOl2pIQjsuOE2gNmWI0VhXlzXvNwmWgSEC57xYr
nnZkhS2HTJ7UD4NcpdpgN73b+5+JM6AikgmHcdkIckCi7huEcPsvUTH8C4A6
KulYScc04e7L+estKK99D4ONMNi9h4TrVgws/ZNJK4xmRFL2sdBiC8lQVkHU
usNoTPsbt3bLf78deVWPOur2Kp4NEcCcAy+ZFg4/8uKWojwREodTZzrbXnGD
kXO7k+r/W80oLN75qtLZTQUhdFWWA19Q3aY4OVNMXC5NylKAfOc1jpQrbrhx
XEjWObZcthW4S8mS//4FMaO7KOCDUKTlVK+DOrmyuz0KP4V5Zq7CeXqGT6az
HVKWM7nUMLbHUH3zojo7pLVMt5NQ06prKaMnQQFUxb3QKa3n53nw4oopnPSL
qHjiK+ukCsrosMJwvtiE632w8aDymcpODM4UQWK9gWQ2EisPuRQAs1qQyNC6
a+Jhvv/iP+bUPRYhsyN4c/iLLPUkxZc2I8jX6pPferf0Wgl5aQKbpHc1/RSf
vDb9XHt8SbG9Ps+psXma8WKlV4v5uKvT+vno4DEJRe94K1ijXlbGoTm4eB2s
pOsfpxPwM5W/XRReY6kKIbJhdCPFR9S2NGTun40nY/gVJE7hOtGU6P1FAF0r
DE6VAOS13TUJklJ7109CxRaqvQufsOn0dKsuZYAtxjWbeDfveRS92uuWYNqu
AbacHFQrHe7jRYEkhA06DI3HuoJ33QWp31ZHxZTDoxg4UaGKt74B4ycPR6Pf
9nBmcVnqa9/CpL5V27ojaK6doA39x10yDZ+g39qDwQDZ6ZByzvz+s1F924SO
dy4nsRVhR7K9A95xQPXfADdNLS/hu2tsqDrg9ENIp5dkk/wicwn21ma9MAGh
QY9EBZhodpe3O15KSp5FzRM7G9/2jpiUksZ3vwxCi05M9sh7yLL6AjzRQn6b
Y/djxOpVZdzmQHMHd5ibsNPMUdsLtYMW0cDRQt9ufr6JKCfARW+v0n9LWZdD
Oj5H/wuiOkNTGfv5+cR6lMXg0kq4T6wWWupxzNbMt4VGKc35M5xh01pOtrft
H1QZSY1ijYnbI57+tC5rJ41C2be77AvCxHx9Wsz2sBI4rGjx0nTm7HgwYvEL
yd7iKBAZBG3bIZX6EcuopvnmMBBTJx8/z7C0P1ANww7QOvWxcRaVPdrTHXnH
gIcJJjx5Ava53w2KGzynBKLYm7gjilTehBh6pQSNxClYALXAdtwWEDdEZgmR
A4qyYbBQdlypXa/OKU55VtMsfYNPwAmgrTY6xeSgcW3WC40hlh4t6vv2t3de
PO3eX2p3BF7CiCExebty6A0jSuAfmxvDjYRa3axYKs/+NCFOucXyjpmjsla0
bJFvbMYWZhxRuosycu/U2QrwIvvpCqdUWBpP4LBF5ULeRkByvaXsDNmCiIjN
huOEd7pEzxeE79+H2xsBhoItgzwTDc/Z7Rf57lIHtw+DJj9VfWCYi6/gt1nz
1GUd8rueJQCKuiOwn0Q6uskzXDly3FRx2VEVD4UHyWV+yZtSzvWQ3t0laAa/
kKs94k2ytulEOe6kMAKIA5UbgQDK5o7MDS7b0awvWjOgN2FTOu2BvVAsJdO9
CITVThCw2IIk8M74wtP41EeByETfxLZV1f9s297SHLpT2efaKjPHX8gG17GQ
XkOBettTbaoPHIJGdUsQFvYox7klC7mqJ160ujnDZUQas8Tk09ayAe7gZN78
o214l7rvKdm8UGkaJxqfkqhN0azwUEf/uJO/pHp7Krt/wg+hfoaj50hPaFjw
Cb6Dha8bKRirgluU95at3ou/lArNd96VOAJzdm4xQIAzDxPfeKgQUd9vwvEO
J4cPPbwTgXMq2OgcPB037WQ7d+QtIWVGWMBTlobQM10jSVMlmbnrkM9tz8MT
LrqKAh33oyMqRgGBmRiozpsZrDX+xojfW5rTO81C1fLycd0MUXFQlBfLyYUd
U7mlZNGigIQhhRDPjzAbUoUL4HFKnuNm6/9dJIBWmAeZnT2kRHmsMy7IhrOF
yQIx8puWjEAUy1UJVsOLZV7gedluDhqB0Hlc/HW7tFmYWtLUZIlUzByQa9JH
LnOeRqjFYxfwe6MJFfddmiuv+xS8yIG1wrJxqVQU/ErXPLtZw7/Yzyy037UF
GdSX3YPyvFoF/rVshdcORWdWKXm19W3eaJmAlnpmrGMYWnI1enjzuF1t8EY5
eSm/R4VJkKuCNwGEEfhzc4RKO+sQ96zrJiENRAExYvy6Xnsfe9F56zj4iNuE
9n+8Ei4Qn6n91/QcoYnixjrEh3oN4I80h1H4DZJymkERrcrWUVSUBkUbiWP9
Er0lbc6SlpIJT9onsHxnfo5f0mnvHT96IdHijs4+xpvN9jaFzhC3JB93GeYc
93i4X9hoOtpyku14Gfe+3dup+qEekxN8JRrFRqpr8q8L2uECnDby95PLXmCg
dHv6Qba/9gyObemZfgS9kEi3vFRJ3sKSfqM0Z82MjTGWhu4+GLppTAzQlDIy
fZhXL3R6RurCieitTOjUyiA+4BAtz38O9AWKNppB89ymX0w1gehXY5fXa226
6454+t7hH441P6RwkUBaVyAXVVZ8vJVLbtIjoLO44it7UVPutxN3QVGTcRDf
6cVnG0ocu7D5njceWwits3JT/QAIlHsyNf7/thwKPhbcbBTLFZQ2mxdPVzbW
Qcoygqsq9ucC0WObK0nLgO1oGpVALBlqXl29KeDxOseCqlfdtmamtJCAABLD
TLIqvh0WETnGvl+soHmq4WLwcWKmuC3Hluo7h+qJEBA5xhAl9jZlZ0plZY1k
PACHU0v70a5huJnBzDGw6pYAF7NwPbU1zf+r7twcXO3Fn8NW5C9j1vKwgu0Z
WOzIRlybnfuxbNIv1q82WugkI51NVgvawEntkK+8juiNo8lkNIiO/uW/9Tjj
uNf7sZMARkHAIOUMcpUgSD8F3UWnNAHFnUmtvX4zkblYY0ZhdQ9wsQdJelUe
YwH8ByL+MlkCHKFz5bzwjFXJSWUEVWyfKFe1P3DUGU+7+loRn95cVodEU1Bj
LrAEjZ7nmJUQdPcK8lNNgScWh9SePIClkchhgQ1hBMNV2QMyfLoXDjPnzkmR
5NE4MjoPwGtDph4Ft8tEdtL9OMiqS/NF6v4EgyZtgXx8C3oOIcVw3751sCaZ
Y+/JTNca1aNKrq8kxtc6h97QeXbZkit5bVSubhE5Q/dGmY0Y+wMpjCesXnBQ
AeEi5u1O/13fcLtWjATvyvukN6QcYOENUnWD+SkCAyWXif7qlKU7Vd6XyS7R
pjm657903GqjCsFMnkTMbCVm1cCLX+95+wNt89GUu9GJgpq8rJyjPLOmjmN9
BSD/S2741oI+i1xhDSBx7PEX+FLl03cf5Aa+seF+sjVoR+OuoIGNtrbOv4YQ
CGb4cPF/HqkVCcEwStpyLDihQi42bPaN0Ek94RVrJLq1fREfytHGgyiAsJk6
7qsN+G9+T2nuQIlkeiiI7sKF9ilSqOOtul8DQVfTNVn8oasSPXb95Gev5H9M
YmSe/UfnPxpX8K2PDjXmo2K9ge5Whu6utH3Z9hAqF9A7V5aqz2baJSPK4re4
7clFxQylRv6bBnckB/jboJG/oIvmB19b4dUEyu3Xhxlyo+M0+WqAEZ5cvIdA
T7HWJWB+NbgjecPj+a8AtYi9Qb32PerC86InSHzGjjr90N0WUBa708RSAJQu
deMo1URnT/ksU5aX+c8ihLMKFOPCarrJu5m0r8sr56Uiqde76s2CTt9enYJk
VCgI6dkN4Pucv9EJnjFhFHTj9PKix3nm06Rb0V14F0RPVxwoLK/iojEQgcY5
jqtk+XfDCXYGkVQHfRAq8VTCTuTn4qsNrjhYsuuTWqnu5Nu3biqRpeD5ORF0
yFEnNzTAHTMfWrv1VIVId9mM1f+IYdQ284ZRtIgrJfy1AvATm4gegvR+sBCN
OT/MDxCotaBxXTCuDadQGXXyBrUmKdDliHSDAv8v9+i7TZoVPGYMV0ioHvBX
miEhSeUL7vK4vULrzZtOfLAXE3UISpRBZJbKtXTeNXVCN6ydo3bCErM3H44t
uidXmttaA5J9AmbuHSsvShzDHW5BtKBKgNkgdywwlsK2behfMc2I4imR9mwS
OETqtY6gN+KMTQg5Xmig8V34aLf8LpLEf3DEKk0H6OXMV68Ajz5wqoqMC1gU
GUa1iUcU+oaaZOBY4MlbE1iOQYDsLAaOFhFSIys5CJhj938xBxreeFvRTVsj
wOxLY8nP9nd7eHjoHxC79zlW99hwYQ/QPgWkQbnstGfM2Rjg8jMi2WBNDpfe
LtHnRu3/7ytzG2GQbRgUCsX+D31nqfrMx8EalbMe8ZX8UZs6UOgMORG1vpv5
ZYdfYud0dK9AGUzY39HkYmDaGmipKIs+9PUdam9VTuGVxu9BkD51iqKl+/ej
IuahThow8agzZOQhvBPAsFT1zc4/jhxmpVaEhIBTyER5EKLqQPxmEPz4lMKT
kw9siQMXFEbf4aJZRaxsmlMPhCn1RpbNSa+tEzQ1V6ybf41OWQOEiL4El/Ci
2tDJvdRN/4Zgt0DfwiZMN3Q8aTlXetHJKz64Tb9S2hvrF3PBuoph4YtOwQF8
Smp/tlcZRC8E5VFfE3EOKo9jC54+CDrVdK2X6LQMIJ/AsoSZipSNRFf3/y3X
x9OyMDB9bvZ43lh4pu9B2fbr0mED/cvyq5TARpBmE5eHIxmz6BmBujlcsDQg
HX3rCi4Fmk7ZOOcgEnjljYZFml+WKfdXqt2WKPbJmox7QxRoErpQB+tQIomP
cYW6Ydz1Vu/LhBmsyeXrvFdta+dYDBFNetdU9zy1CxL+7dQJHLDqIPeSOz/5
Tt8GpExHuG75tg7PtUWgrfj6na2hyAt6gd/m95WsXv9do3sMLym1uyak2LfF
pfyt3Hjab9/kaVpDA/9Kz/C7DGWIz8IW0L5YlRt05MhsyikRNlVKnQYP+Zho
KzLzG88i+ih8uXXdhOBg/9rNFNf4M4xt+YBSNhVb7WJ8Y47VJcVcSBYTufQs
tXMWAHqjRu5C5DEQbRPfhp7UKov4fRyTaXQdIzl7GihY+r2+7Idn+aNcekjC
oh89uW5RCqWzc90OAQuOnimy0nNvI6rbDUVENdFlZYkKQv5YloGIAQ9Ks2y/
V96cl0K097J/qFYf01HDo9EZhcYcIRH8c+hOueBbjgSv04wF52xvU9QgX3TD
q0nJlbIcpYX8LBrvaaVSdHbYMV1i+QbeP1rIcf2i6FFZ4TsFS+tIPTRTYT1e
aYFpKJi4u6LGEeZKNXcaUrs/tVNshJVAw9JiGcSKTzTSr+WhAHEnaNnMbMvU
XlXyL5dhdD70JjXvvKCYfHaBpp7g6rda93jSl4e5/6c5jef8FAwk2Ew1sGj3
Aq5if9QzZO5l5RktaXHZ4mqFU2y49QKGeNcMxeSKi1hFSDxmHX4k+U+dyCD7
gWbFLTLeZKhP3d8E6vceNTNBtf5n0Kk4Kq7uyVEGxeR7YfENdQ17FRTv+AZ0
ovH5JnSUbRx8CUYQxyLcYhk//+W3Ir43pIB+OYkNepPZWmDX3Wuc8V8rqMuT
DVoKFuqmCyYHVqPFX8GqzYHXW4V+OTuR2S8MnEmqDkh/72E7b0DINcZdTcgd
Nwb44l2An2RX3psKZdDDmtQQjmwyFttHJY6x8f1D8yFmpPWBJWWiJ6k7VS+R
etjuaAnoLyPoghdtMqV7aGt7Jt+ZfodaP92tVlZJggcobgp/kC49q+ZaG/Xy
gAxvfe/SQoFFPs88X6OprlANS8oQr/nsOdbKBIPQfZEeRW85M/dSWNU9bZ/w
J5P9Mpj9PALYpj6AL67ZjJ5ccWK+qZoOQjENhY+MywhL0GYiEglReSdy3JGi
DT0dNs0wMKlXs1wP2hKeyiSAMd+bHTQbbBsTvrvyFjQrJfSqGaqKjG3b5hTe
SH8EBRigUFxtXomzOWom21KraZ2sSfp1me1y4eU9f316Q62fZ7/FKlMmCwOg
W+X4VN1JDuPlS77t11GuzVWyBUMm8AE1GVGNUNLf1GCej/Wny3gnCXFqvPn2
jI2Selx+F4BdP3wry69S/uGlYdkKPHj2ulQfYt7LkH6caYwltv/S3a64cErr
Z71Rh6t4m3DwalzTmV9dnkqKFGb+KF4xjOeioEVHr5AuAn3i5rVcbLshPAjz
aM2QV4nB/nBNd6AKxZ1ucrBWHihPQjZaLP/lf772Vd+iq99jFJYX/e+vEYyb
6u87OV/hv1PqgCpkekx1Tv8mSV1aVPzM4i92opwjgBo7n/7iiRBKVnvwGuZa
h02BntjqBoRTJZilsy6QBKrF1uhI2n0mxjyDCb+BZB03ZVl+kh7geHi4hp3l
sJ0AvqjF2blUs+QXH1/HJN2X1DNpcW4CMH9pwX8Mo1OeyIRRqYqFDBCbnykR
ZwqfBOE65x6+BKsE88g6fOMuhGyin0mwWTRpD8gJ7ah2KEJFugfhHCMKxeGb
EcOQ+M2EKZji1C2uXDryfTY+X+B4znuo5oYYQMFAS+NE1R6uz2WrOwhHEQ+E
9LHNMf/V6vWo3UQWaJYQr5SqfiiNFQM2MeoeEoP/7nRZd9s2UH5xLSz4yMaL
8OIcEvC7FroJclN6u0g+eW8iucPWZrJds4nHyPKJ4HePA+sH4+dFPmXXjMT4
Q1Sx+2Ck+I10eP6fY5aFTFyoNAgrxmSJ2tz46BE7NKkQsUonDFdapm/xnoEi
LZjYBJohRrqolckB+WOtjCQBdoggTE4zzZm/27seMP9xUuw9af7JI7qPGaTm
2QlmWK+ipsC+DYu0yW5XMY7yeoQXvzljPczzeY49yNm9nQMzjknn/jygXj7B
/VrAFEU4r287phi0/AmQztG9mtqlRX+jsDZ6WAYPbCi0D8zhgzTXf9pgheeC
mZlqM0v0BdlQ2+6ecdfQCibtUx3Dc6MYCLmKVkPWcovilnJ6Sba1cJdRqc5O
pucWC6X/KDkbilLU54Flimy8ysXlboCJtJhbfDYdJl6vfmAb0BbJ3hm+5di+
EjkVRJOPHdixHOIQDX+MT5cjn01Kovxm3Dsst/NByFJGT06sHUtjmxhk+EE/
/xgAHTNV+8MNEAie1mw53+oDN1ECeFagzXS5+WGOdEdi2tQ/mUX79nwF51RY
25d+pgQU8K/tbUnhCiwDmGJFuKthiqjy95bqjfG8rAuRVCdlELT2/knLy93b
iF24YH9s0ojaoP03iPkEb3l+yZraa2ZwmBID4AFbBV/CYMYjpRuPIwmJuE9h
nDjh4Wf+FTCNIh8Wyk+SUCzaNPhSSgEESwaqIoiWDmbjg/z/OBmdxaWv//4O
rMkZTQfzTCQ/ZeAtVIvRJy6xRODYsu3W+na1ka4DRHeTUbH8r3EPNv2PLw1v
7pp3+D+aob7FtwngRWvVZbRYCMVwheFRdQbIoAbhrC0Vq34c9NwZRkOKPTUH
VosDkKlgw6Z3fX314eMn2H2b6KA/PX6iptMT793h+kqcgDv6enUXw+fcjIfW
2Mhix+NWM+fVVoF4hxtnpOwaW7teNHFDr3ALefLDZKpgpqhQ+N8l4Gfdf53F
6RecPFY8tIDUAqgQxHduxd6bXu4MS6IuDutXJZwx/zN+V8QYFRqyNmC/yse3
GrYvrqj0BkbTjyE3SfR0owoms41ktVfJsc/uJ6blf54kPTyZaY13arPtzZ7t
wlCszDGlczSfBV4UQGIh0QGNrY6elpSFaVgPT0TevgaTE1xnd0VUrZaWjW2O
KhFfMGUhQ3PLbi9IUeFkIzsBwzBuGkcGWSTe/eOGeKKFDg7QJVqYhB5vKgff
bL5Xj79IQCpDQ7bHNm1JSTD+EfiQEtXOcpENNauEDg37Zlrh0embgG4UDfXr
lYCXv4V0pdLg5UFM86TzdYoBn2PvasyRIhLhJxmf7kRoYCaoPFF6Du06Hdgs
Ma2mooXaX/a7F54ZS4D5yeNK2lHffa9N5lgAUqwcmOzMSXViSWyN1iKfD/Wr
kVxGFSjzR6wfygKIlEsj+TtUKSdXjOFRZ57r1NsH3h1i0Z5+txHOzS+IQtMj
0Ug6JLM1wYCcU9HmpdCqkDmE1aAMq0N6QstobSx87pwF1PR8ojeIUxmajr0Q
Js9mXBapPwpJm+JPckUg2+LZ+BkcvYrAHzMZ+CAI6C20XfBl4ewjY/ypiuaL
un48bSwX2wOCI5pNYUfFoWZAlm/o7eAppg+GnuVjh3ibqV/tNUDlAeLsrz7n
lwKxnYPPNQEu/FqCHeDcMMeomqOOpvMUWigihmNk9tPIr23cj9IQPUWOL+/E
g6x4i9P3r5ZYGsmyYjO+UrFoH1tPNpfw/16t74sLsMt9dqLzm1J0NG1aivSN
0lr6+hJ2JP6I9yC4RXsx2b+tJDilieBsbQRXbKfiPv33Yl27zJbuzYSN1xaT
VZr1YD4St+J+SZhzV77nOVcKcGzguE7AYrb64Nuujn//P0k59H06X3dAsRuN
NJUTGGpTjWhN0uhkHnOeh0UH6foL3UaA3I92+mXDUADOtjmrGIuZ/SOtU9ul
KUAj1mqiyqEa0mwsQF+HVpw8yAVEoV0Ly0A0yOWn3n+2+VfOLSz1W3EGxSjk
XU/jRwAe+kUmsWAosQYq8fPrkVZ46uoLIt3UqYvd7ZuVC/A2fTdtAIx9HV+E
8kefrt56fjYO2hpn/Ld1EwJEGCo1gEK8ZBqAUfwQl4KTOfzOdx5dP69TmUSm
qeskrbtnj1g5HdYYAtgHP7xkEG2R7EAnLt4xrYuCbohpA4m2imI3v+EuUl+4
GxfX3Zjp5jjGLAl31VC5NMlsVJcLMahZpvcUp2G20R5F9uevCp7RrSNxfmPO
AX3RDinHIbcWGDxNubZkz/PEMkip8hkletJUFe35oVi5JVZGPBK2kzFdVSLh
M/f+ON14LZ209NAQ9pYsLKQJXVOz850f0cptp2JPdHtlfa0CFQAY3okfb6a+
Lb2tkaJ/EdthljkXdH/cueTUeW+ohCLANQfZdGma2gWEkUjcWVTDkMMbETpK
7vE7Xjzsg3TumjR9GFe65Hx92WmCtFjW9Qfg/A46U4vVnp6po0dca8CDqxmr
NcPz9WfNWmg7BTMjv62A7CQ2Tc43LjS2ABCWD4C0Y1lJXCaDUbDXOiz9FA0O
ZB9RcF7a7uHp7zRDX96SZzcTchNeYbOvxk4VbuWXlx3Hc3TqMn4rX2HYmvhW
xP2PczDvTjHhqZTDAzxBWXvqIrMkCaGHAZ6ZHw2uzPkePEcU2a4ukNI3aMF6
PulhAtyvahS4FPI8W+dALzlajrTixjfuWZEltoh8f76SyNbd2a9PyveuCy2Z
Fvye9tUh0sl2khXbHzFV9mqWIEsU67v71OHbwjy1IfaiQJHiK/CLPOEkYM2w
F97l+KBf4Z28AvsRpRwBDgP5P+MZJ1abbL7S8qXB4qM0iglrVjwNcVXTRFGR
XytoRAmJQSf5uxjkB9PCUw4NlOZEkS6Em7D2C+ajpDs5xRkWtukvCLbmL7bc
J8v5ELT8mfMihbN+RP8MoQ17PjPsaa0d438zk/RV/4fRCxlxmyl+hIBmhXuH
dHQDQ0Ea+rTqIHtaLg7hcJZ7tEeShFI/EVKfJbDnuE1CEqnalFqWKTnjRg5F
YAxXlcG1ud8efC718+GZ+hz1tWqB4cfQ8AzWym5dzmfaU6O38AsHZNppdZqM
EoAHkI3hlmFrLgkYmMm4rH0kFYXnhoDx/GSU7i0MWhCcqljJg0aDtlQpAKa5
zNELXcRP/Ij+QoVtlGBvSqW2XgAoDRipIcdfWY7I0pIpyqS9Qbh77YtSUPey
HVnf/jdwrKfEnJKPICqzde2sNf4BGee1rZz6KdgqHD42fKYCr52ZEVcV8qeV
RGnrs7/mo6ARJR7CtawV5Ee9sx/G+qhIzmqGgzRI0TmLU5a5C3nuankAi6dI
w4nn66wzGu2CgCc0zmAWZkEBy8n2xgaWqYNLofobKHiVctDQJ8hMRg0RGHuK
qi1BioJKTJQMoUiSIN/EbUBIKmJdoc6qX1fd1TGLmXpPwHE9TaJEFrHcrLPl
eRAoaBolUyxGskq5MCTE8mMVuBukJ0T5w2/RWoVX4UQqQtOXCvpEdR47xVln
w2jTmsFQj1aA6u74pb7bppyulmxjCZdqRVLyGpsUL7Ad26F8Oo6Ns268F4AQ
ndNWF1P0gotCJ9vuYE/LeeJL1XmRkMqvjN7Mo6IsvHFl0JxHaZdhqMMhKJKX
4cncRhTAOzrCuc1dpGSnmkZddTMOsff5wkjdmKxOhc5fY66v9GV3Ogrp4OC4
odN0U0pFpo7xte30H0cDqrln50ftg0U+1aU63fzN+pV0DXjAr1zLAzkeFUN7
FFJqNljiTuZnpFliLHXItkaA9vyiyB21thJBgvaai4FzoIu9BZ9ohKGhcVMc
KSG/OZOkTXBpbhgEXZA4EMHCHZbGhHI9ccxdVSK4FWRllT/HozHliymm+ZCz
rjddDIPsmgya43SwqZYoW0Vzf3LgvshspPYu0gHWLidT5nUTnJz1599k+SNM
G5mpOy4NmIxsP0Eggk+ryF7GSsjBZvuk2rBo8alDpybAeFpMHsomz3gYkM+j
ocsCwywyfKzTgHRQxc4l9yUf9nH/RWDF16rVXi8eAHJThnvoNwHzj0TFoDtB
qtWec6M5Ii3uXkg2Eawff9wU5elGYKaotLwP2wvYALjfBJSoVsWj3n0lQ2vX
KgAMrEEalwX6PLlesjL9u4Lt4zO1uB/I4YdAMXFRLG5a6du6lBKyZuhwVfvy
smLdZPVDi7DnneT0tGQhoRxlK3RHZvISTE6YIYmi7IV1YeXflv9V/+sNBkKs
TipckoH1qVKjFn2nmBuaoE0VmN7SLVtVnC9MyWfR6RllhdubcZ9XbabGn23v
68xuWqdBmNkPWtbQEiNM076UxdxeM4jZKANypPgm9ivGqcI55wPeDuP/MnNb
EvKq4q1wvYI7yvvVY7+BqgrLdZLzjxxUtvgz2QedY4iLP82g5/6cpen2+WLp
KI//u5xAvDNGMJGyXniJIFcpfq2fASz4WqLiBJGXjUIQIp2+gWJeGoFMLASm
nmw9CzrHGRwb7UTHEqvyQ8G33RvD4LrwVa3CGi2v3paShbqZGmL3n7Hv31NQ
ZcBXXRm84ekbVOwgxqlCh0yKFLcZUyF93qF6nqA2JNsxgpafTci76yN8GXDh
t6ctatZ2W4AfIX3hZ/nHHsGhFt2dWniWssrSsqpa2cEwdI9G/GbbCee/gwU6
Klpk6YT91b9XI15fo7zY22t2rGZUHDBkdI88cVciwwE72wnZdon+zvXbXMSh
s4xtz/MPrPwkaPD9I9H17LI7pZKHMyEzIkosxJ2xhn+3HFWyCD7is/ERGSyw
GlK7PeoOR6LiJA3DOeR6j8Ebzmfoz0GUxQT2gYaAYRdfxw5LmdXwyy9m9HH0
+8BBvzr9HVk1FBAisEjCmpfm+XKU8pWpViLJM7mWc60z/haq2amdVFZYLp7h
jX389rvCY6TAQVY7zr/d9n+M6k2Tukm2EycHCzIfHMoCrV1Lxt0sseUjXQ2s
0uMBYvKDy6BQPgCU5BPIbSPMqt+O+11XPVY6bFlYbgs59IcJsT5/SKQ8M6ZY
TBhi3Y//laSbueg7HakGfC+B67k1TByk7Ohe96OzlQY2xlFvRAO6+VsgvgPQ
CHPqCcWjp+MwbIf3F3o1/VSyoC8ashMvRm4Tnha+0vvuOOJKuuhHJsaoqOTh
ZKK4+s51sajPjCCZi9JYqoHkmKnej+Fi8ldGXox4aHY1NlCwBXEtS3XJHD1f
4txj9e0tFxkuggF4jMWe7SgpsPUDq2axTPrxIpVoaEoB3FgfuQ/ItxMp0SOn
mVvL8W2LzscKq0V5p3nA5/77kRVV5p1Jbr6eboBodVpI+JHPrg+JVxxmNeyU
BiaJf/9cPGlq45sJm4b/JAZwOnqbqcYMlaeDllEZB5MRuKH73A6vTQjmOuMK
OMK/wwNYH//2V33v22AfPntbo8hk7vMP8IMlANE/eXG92tNxqhmDZepigVV9
hH08Z26+OLBIRNNUQ+SQxTyccz5ZUx8U3N63mdWHdoqx9AaZun8TTdDwIWqo
C0bNPlFCL9DaqeTQZaTgq+oGI5Tu+IRt4rbMHJPUxBMgKjO89FhPl6RCdNFE
TeIjouF2OUa2NrWPbiYE8FGxLInUm7XPvsKFHwc2ZWED8iPxETM/vw27Szmn
rd5VGpzaofpewFKXAA1x1dAuIm+0+OZe2Gci8AN0VR++TXmUKwrxw9yNw8hp
2yydBRMg+tIg/kVQocJ4Pu6cGbH7ohZoxzSFq6cZEoJItIUB9i5Zbx0x0+6W
hzX9dYzIWoSiRDIrUeGiGlsTsZOmYBBRKsmU2rdfE6krC5GFwbOusYsasZ7B
iOpfMo4+2GdXF003MMar51exm49B3zxidlXPAo/kcuJ8E7TM/DX2LmcpiY1z
cbP4tzslLgF93+jqmB169XeUfqT0F7hu2hVAQJVeW6lVoOrV0Ae39sIzi+Fx
xd1Jo5DncSfxwBaMB9Cj97UHzps9Fc1r9gYkzD6KMRYekC3Y9WulSTowZDZ8
U1pauI+DsHTpg9Bh7gbPceuSf368E9Q43az1K6UPYe1JI6YjENFMnnww+qk1
RlUZLxJDp82bVS0UXIMNuJQfnybno8HblmhLTti65i5ef6JriAx+9aUtmJO6
Z+oijilbTuB41HVVOd4gKCPaAlDSLAcdHaL0HFBpMPZi11xvkkYflIFXUsKI
0Vt8wvV/jZ7KlqG05uN991jGaHbaVbjI4g30gx9JL9ebsqWRYiyQOTYHrqo4
YGQFdlhMa6rJzVCtiKLF34WsSs1RDdVo4AYbbuyw8icBF5k2wYcdsNwxeL4w
+8Sp/rNfoAsEz31rDOWAMR4c7VkLTEsl1h0PXXqa1tyh0AbWv6GGj1iVEeUB
RgiL0lv8rXtzzuULIBtxjpUb7ZLATdq7uyGepoUNWqbWmwp8ZbV6sGaslkss
PN9Bg6PHqiSKvoua072nGriE9DL525ZRqjEhilCKpnBggr4ytt8oRC/WvkI0
eOYImPNWJPcBAvCGrStk4LSDk4aDxY8YRrsZiUu3KNZt0clYvrMgAK2ZbWg8
MgQsa9858ILj+Y6DpOqcOJBvxRm3kOrzfwn1qqOGzTBmhvlj9Eme1JmRW/Hu
fjDtUJK7sdfK+3QOyWSU99o7nmmEp3WofG9RCixuABRJY/v2fEly+W6DLDbR
TajVnFOfKXm5UWqCKC6H6FvoKUrtBKImNl/gFgFtUUBL1EhkmnAcIYEmjuJG
vqs/gppfQQBmUClH5zCMZEeCsqM01Z2q0GAkr4gV2hU6fFFm/AHVtrvY+oq9
fLv7lI2K2GKPXCg5fz0GPzyR/l1Xx5IHpWOIZegCUz9Fq40Yosg+I8Vgeeme
rvjcS0eQ751tv3nnmFuwXkPDvsnL8pl/YDEr+Hcx/nEuhBIWzeW4JEffx74I
0Z4Z5WLjTAN1svlhDPPWjAqKhnh43bsL0opM2XPL5eNx7uF2fYdGQh/OcTqH
ZAiwzmoJmekZHe3BvEtBrT4X7ksHSjkbLi6mRxEpXhFHGoYJimq42zMum/ro
HqOORMX0KgRSJtzfKHPg3hP+geixU9AyjFlvFvGR/nsm70yCscf8drhZ9AvM
iY08pmk9gURoitPj52ayactKq3tAg+JfhMq+rX8l3yzNQ0I0nT3Ibo+IItos
+h8GXuguExwk+ZG0uZr1PwNoxJBub7Z2ldjd/tVPfEeo8+ZYPj5dyH7jLT3X
+FB0qZa9owzdZcZAEclUW6wnirGPch0Pgna7ZxB4CQO/VGPhUr+azZhcEDDi
+1+h8pF9REYP9xSrfCrjDJPXGr1IZaxKwbkpGzXk5B3eT2wCMj7DTJ7bsyhL
cpDA5d96KXDrCFVjFgrsNI/FC+ciC6InMfMyLg5hdXflj0ews+odF1MR1NMN
ST8JJ1bGz8HsTWD5ytK+RjrhQKOG/4uHoV7/hgSdt0ifS+cmt9BOWhhhJgyh
aTT3ZI6Etw1aQUT/WGNh0Zikn0xHNpLafJdI2rx/LeIActfE/ILVF6dRYlr6
f6PWFBNaM5QI3Ffiii/W6B1mCffAthW9fA5wpH+E7uaLN4iavBx0cW/cL27z
FX+2w651of99/xZObeB0E5uXsixFpV+oQn+UD+wzEE2dMtYR1XhT14p2RXZH
MlfwAFEJJOld7/cdUM6sidcNgT9O/9yh6x4/j5EG7vSUg7VZEaiGN+HQIjU9
tujt1zQ/4eCJbsirtG2ZDcpieQpfKC+jCe6GYJejXoA4eNNZQ4aHv+lX/2Dw
tsDjEdFGcVW2jiDhiWKSEy9Tw2ANOr6TwawKAfAb+iTFz6ZPPGqbOULSS0mT
YTNhWGLGvFsV1b7WnJoyY5gm56DfwhKcGRaLrG/aeRF9FqXEHyARWOMycJ1A
8ut0jbcCYdnVvb/EbRQRS7DJmjFsELL9Hq5t6/7vaTpiyN0Nx8hBiOIB7NVR
P6Fn9hX4yE8U3hZtnFnd5EdCyEulZK1/UcUUGpkm1kmM5I2Z5nyoH0ZSU4vZ
BY7dJGkHpUrAzLMqOcgtTgWQXOj2N+NbOuBhbQzP97Z/Sub9IFjb3cTqkvY9
cgPpYfNNhaHydq0YnuqldIALE6IJv6hn9sxeuil4SgGElQdpapfifwn3bVZN
rWc5+dF9RYMudrjBIlurGOCbTrANSI1SlRzJ3lgXY50SaG/i2X3sJpf30syz
yTXIwzQ5nrSqWwPApWRRUTvo0Q27Q3ihtfgI6X+Bk4QCyp8TdqgYWWjMjH/G
Z5CRdagz1DkJ4Oh6W+tIT0njRlarV3FeipR7JA1sKZZIzhyp2hD8O8PaACIl
LwZ5nSDbdFMRNFJ7wAJvKIKDPgiQYyWI2aSKBB6je8CCNqDuUYfY9qvaVg1P
JK06VankWseGdRosNQWMeJyA3zNZOP7wTML6FZKQZuqaNEu+LL0EcvJOs054
BzSQXiXu1ry1YCqnKRCS5UWrkccOjlp/nVgG5bPFd2PSq2d4OvlYjpfzjqSt
bSMhOEECDwO/vED09cL1Q5EDdsNxF7ddmpKhb2dpYOGj+APYr7VEulBN8sgg
2jier+220TM0AnCTauQWTEjNECBchtQEXnrDznrMtm0Gb2bTKmSqzgxv8ocZ
Zm7DmSyiMNjlbwMWleqi7JBCiw5RQiFvg45BFjTn6h6QlhjnWGFE/6rYx4PE
rpY96KuKV1bGlcrCyHzjEpTNznnm0JqJk6YyzHrGBPF3GdQ0IRtw88/yyq8y
gQK78lei5R4N1WXIqzU6QiKwfTtFr/216ozJpTrDwbmzsIH21wZOD/XWRzCv
JN9qGdhfHrYMtt7nywLZQPNA+Zdk1JRapEYeYHWiWDW/mCHgAFuHiCcW7gP4
U4IXLJF41Qkt3lOYDkq89cDzxSU7Jv4ThTapNrWmxXEI9zEHCircwhyjJlW2
D5XNocfxTnjVjUs6LZ8Vm7NSSXLyhHLWL2TO+RkSl6++4w1JrviItUs0+dua
Q26gQW9Ga44CdYyokXIBfAt0rcqw7KOb9YemhJCkiDX5RRYFYbbN1CPguO8s
rQj5fY7BNnBFykV7EQ+VY//Dn7r+NlugiEOC43Rgfybwiw0BbS+arscu/Vhk
v0ZOFbbu25JMNFbDvQqKMpbEz1FgDJ2qeZjpmUDAoaHJwrWkeuhikeVAinB5
L0Q4zAYtB4ari/nhBaLwhtUGSU5skaSYYTTt6K31/LQMExChNkT9abuQulMQ
z8FizU/rpRWXee84iNyUwvjz+LylC4r4o1ePKX6EeHgrM6zbO4U9+LRo68aP
n158BG8dlovJNPK5N0C/U3m6cjgVkGKELhw0AhcXB509q4/FKuKGfWYjSSsp
z+8+KNHRtve/hLkyAP/4fzmGpMBv7KAIFBFNvFzQ/kfirVXIWla2DYqZgG3C
YM7/64ISEs8CJW1vSJk6gd9v9WsxDGYgxD8lJ4FQ4YmvuVbFrH6D+66RnDt5
lioFASs3yBr8ropeG2DciIUWywDJ0SP7E7Ar/08xK40+UJT5C6A4geIY46rH
6bL+FDlZlmdQ9tEJTwf28VNBFJwNpwRSFwawYq0f8Wz6BAw5xzoVISKeVvgj
cJvuknooTtegRTM/QUWehWyccnjbtPSnAq9qMUOA4JCA717XPYOoKvcAHhdt
Wie1jp1zLEh5lQDB87G2AD8vg+TDcnkmvmsHHsS5xZf4cHpQzn5B4qyQXuKX
dTiDgh6K439AdWLL7ZSiEwj6RRgs3BPWazTwZwres13ZCpputfzGvBVxfM+A
+troLoCiBoawlOCWZTaQpm+SmzIDaDjJrZHwNkL+ef2nTFy81k88i2PnAgzN
ojWOW7WuJcuIna9Fdda+d6x04BXlqb2XKhEr88au0/ihUcmcGF91k3ZcrI4J
m1LuXAm0P9AOibCz8IYAn8bXVfyPVuVCzuSlCTsNxfNDsbv48xhJeOdbzSDp
by0uXrIjumh8KGvKODaHUWrT9iQ/Ymw0yg7PIyHSTYwWddrp+3Z3J6WMo/44
l6+h7XVY4krIOLfMMOPbnhAv4yXvNdOItw2lRMrXiT7PdG9adsFTBn1LS91b
97wwAWGdiBsD6r7GcOl5q+EFyZvZ6WBTegpC+9tmlc/Fg+3tGLcs9fVDH/I2
B6uJYoH7355fLW3zJCRgCKguWY5J85PQU0W56Fl+NH/6f7WLDdyaDmtWDVub
8yeNbjP8eY8IDSCFgMwcyiAgfss5iyCsxi5JgaPH0xg4EofF7wwV5KgkmZ+E
cQUk4KGFpe0Do5+ETDW5N9wSNpU1p510zfNbkQP/E3EMsGoSRHgUFPmIVEBP
HLUNMouKA4iE2/4QoDt4x7PCOagRaWLbuhI3+xBb6Y6l/FN/v3JdYS0j+VH+
0sKxMSZxXJJYPj70/ZjY7up/zqaAr+HFfORGQyZU+aAnM5Bq2h00cO7d6AiJ
gmaJPLfnItTIzgJj004Gp+FuGP2Q9BAE0dxln8hJb9/Crk8bU1MPZzdatAY+
jaNKa4aIp/s/YvAE4PAx1Rf1zWJprDoICIJ3+Ng6Q6h3AG5VZBXueYnfEwGh
XSgEBU3OehMpgAtAaneLad41qF2j04NVAXel/0YPNudc1BGQwMu1f3MnAIvO
rPJ3rsROQaKZfG/qz1dUHz6KgprXNloPyo48fkG/ePGYDd31chMlqQUYi9ZS
16MjUGX/pyswKEQMbaPnQzqUNH9YkBpVLqZ5cUriv//GJrHEHH2/1VoxiXMu
jFIMc87VLuK9ws+bfZwwrc9gd6ptZI2VEqXw4cowWbgxpKPNEQpHJYs/kS3t
AcOkOj+btRDZLFxZDc6Otz4m1cNTu0DsqRbhECh5UiZhcfv4MICAd+RPuAVt
2o4UBwOsXPqdfVb9RTQ4fjQvrjVqCIckKmdjMDSAol2ul0EZHLXXhRt2UNhL
8DAAvW7TO4QJ8vZUSiCUS0TeoDauDKoQKzpQGrfrjfDGZrGcbTGIu1RRIBq8
JNUYdKhhgWZWdV6rwuQSfHqS1XXb7RGxs8Jp0736MrsT83lEDY2YvPO912Mn
7VRu/5cZ+nWmrF7JRSbiY4c/R00gcjISoNQoRqAPnxF8iLbfXIyYUjwabCc3
277tDvVSJmXpqW8aVnEifeslv3fPUJBHoghGbV1BVOSYyz0TwtzwuojHBLY2
2pSzVubCuLoFu0YMOCAY9Hk1fyGos3uEicRrU1ktI2vidaS4BzV3A4BW3Ljo
AnF/B2DwG3VClyCExuGzGS9EV0Rct05LZAd+RyYvbrF/SdTndBU/4bVMxoBO
oB88iv2LWbYAOUmTvJficVe4gG0lgODGVUtN2cLxWnyEpH9sg3VwZ4ZNwyx/
Q2ParZqjXtCHct1KwzDylqxyrWPr8sd3np4S5Z9A7XM2k8PWQ2ggbrLbB4DM
/S1qU+1ZDq6WlhAMurZDQa/c2JMquzK9Hh5Ntrz6Hbrqj/zzJU73RVL7mWv3
jy1wblLPfF8RwEJhVRXUUrppEOkcxRBA8MlLl6pz4mwSnNIbwgmI8jYY7dUy
fswJYSVejZzxJOq0cxsJpcmWmcIZh18AhvLFF+ycX6mUYbo6wtjLtoufkFA/
5K4JRHxXJiAM6bYU1U4LEUK/BZvV72hiNksZS+qnPOaP6I4KveiP4qjB90zD
t52uy6O3pJ+88JGq+1zV9uZsDr59FRuifgyc/EEfHAhK8YFR+rMhuFLjFibw
vVgDEOnfgp6qmNqL8uLtl3lERjdwS38ofYv0VadwdToTPWa3iTumjhVk0dKU
StEMhzN1I/pYMOaKnMZXwTPAy78DJkL9jtu5x9DoXFalDb3tkyMcH9/DxiBy
pV5Kqw0wUx2CPqXen2jPN2FIJhfpCgMtZn2uaFnwXJdVdmP1q2/IPvXic9dJ
9gYoBGvezkVkggmtRjjKMeln3S3nhubNGNnKVtEfSIM8hF9g+Mcrlu6t3Gko
pZOw9z+KgR8QnMSY3w+s2p/n+sb++/oOxdb4/1ofrCmdcP1cRw0gAgiIDWBZ
8VWh4Xi4Ei+U4n9K0EFjzbXfR3csuCIW4dxyhYYKKWXiC6AFaaEBkXMG2Hsj
OZhXk9eOXEeg4+WuCCSGwA1cxfRX6n4zozOGFleUrEEHY9hOuGS2czjGzRUM
D8tSbJ7WW+cQHCSwyLdsIC1Zkn1NkdGFJ3lBYXu6enfq1p6ks6MzauuZe1jS
Nnybv5YHtIK2VotrA02SYEkxSHa7LEwQTdXOuplWCbJ4U1ZI5eqxJbD9KFnh
+pM0Q4RUgYopQWCLrK5hDIrVkgIm99FzlpsRSvStFrt1gC0R15YGq4OYWmJu
RtULI/YvG/J8RWjXjsL/wKCktKQGyRzfVoyM0O/5X29jE18im3M6h9LvQBPZ
pw4znwc8KiQ27OMUvyzgzl38TlZsI7DPFGf8/zpcbiP9Jo3j0iBUhMT9zmVB
5VzYN7fjwfSVvZxwo2pTa7nuuVpUCWtDs/NETh7aqyQ0jy+JWkAQqKlfCObj
NAQL0Nk09qW1WLmBKb0WO1sh9Pp/QNmRbBF4Azczavx6BdDUiK2YEHvp2/2Q
96WdJyz6OUhxqaMNxO/7M33CfR1hYJTXl54BcytooXwx5R81UN4lDUWsNcBy
5921LKE5Uy9FPJQ1BetaS0crBrcPNd3WlHe8qeDrNcR6KtS+uNwJjIrVHHRo
10QD2C7yKXQh40M/OGhGSV7zA0N6HSXZPGAKowyFzSYvzgjBKHqW3mTOuxvr
BnaZ5Ksi2g8vDluthGaq/kaX2E4RU5nZOAb7tTrxjiQntgq+7O+oJt/3wPEC
lE+z4bMgyF1aTdwFw7KvnzrwRonQySjoDHx5ELKuqs6vEZqVMwN/uEA6dV1y
VXfF5DbIMwGwzFqeE7pMDzKlac4uRNsWXE82vXI3uOd0ruE9p8IR2hHZMqmD
jy6D0d8DfGKovBTAkpRlgfUMNssZM0lqpZ8YxFeKod3FKcuNzMmLozD+PvH8
4gU9zuOHQjfhj3iyedT1KJco2ILNiVstYl1MYDSC4RshZRvVe2B+UgmHLSLb
Uz72vCdf4TCTlQ1GH9nXq6icMAy03FtpY6FdAM7PpWSacnkuyMEDrRM3R86Z
DaHpNbk7iJoGrNcsa0IMKY7yadlRZ9NKxlLfB7Ox7IRX9j8bVlhgDky/bE09
JK+2mYBGZ9s2jOrtIqABqXDcKiplLU5Ke5s73TLIU5dxwEQZ8TZUs5OSYmM8
oSSERUaAsduZC/42zmxPkqgFGudxI0Jz96KxBhziMWDwoglCnrzAYs1DxFPw
tGz0FaWzv/ApT2ZvNUrEOwCePVydow6/zFTB+qkNZ3vBUomJFRrIXOb11ctL
kAwzVVrdee97GSyfyvgem2+AdwsT5wJBr1qrkDy1uoLH+EwokvG1KXxAdWyw
djbGiUOMwI1bBzjpRVINpbIJSgQTQlVZl+LS32YZY1cN5qj0XbVUSNlB8dGc
Auk1o63i8+qQZXtsl1/7txlWY+p7HMzulGjIh2qkBaBKYXu50+YmE9Ltw8kk
yPX7B/YJGStiBjhURuYPNDouv7DEeBH0dPSvs93yfnR31snggc8zKzEV27i9
l8g7a8UpPhcYmf9fNOyMlM1Vc1epLRh1T2GVB6ROtjV2/1/Vg26m3bNeDb+A
mQRmE8fEq3MJgHztUOB2PVoEtfg1X5bXbkZP3oqjMAdWTWzW6+cbJxr9EtW6
FVnhmc4qY7Xq1Ok/O0bA7VaAVz+uq9NKUshWUuZZ7UkIE7ACCFm5BTKAmg1H
rpMUqJkfeyyg2bF3t11w1xEsigdNUmRmWgWN5+YRQFiE4QDHCIASyTDLMxkj
YcnlRWVqTtGH5e60RH9gSvfzBmSq95lwBaQkWnAsg63hhy6sZEjv2O8lK5lA
grWCtBJ00Xq7yqUhy2ViiBUWaRZfp+s9BITI2wrEdZhAT+uUKQARSrK03Fun
i8MzimDZ3x/xBnqXOLAjU67RtFtuiVLd3gHQTLwlPVpFSzFnfjC/eH9uzlZw
WgpB5oyGC8lDUQXFAeC1fmylf4i0cJ5jtOyTIBKGmTvPbl4UBSgEciD1JJqw
pwljcWUQGw4iVlozF55v8j4UFqAzNALI/+YD5V7e/bmf5bXUkhMBMiEqOLP5
HNxdTDDYG8JzxuoXzVLmo+Jvet442QBJF4zGHcTJrOFNU91zavZ61oqn5AaV
u56mdHOvSh6pYDOm15tQty3FO8rx7oBnhRdpZuWrhCgQRoROuntCSU0l1okV
CUuyYzJAdDkxaJYcakbWaR8T8+fG1P6mGYN/ErFZeNgVYoqgKSenenc7+hQS
j/1amYPNRy4eYVZQw7+6q9ZbciTK2UBOhDcLzzeptani8bw4p8oi9U9I1rS9
gxJ2pefVa1iVGBtEn+JEHM86FsnVuDTd1mIwtjyAWWYqKzNyNalET7fYo16V
M61kDQW3PcXiSc3fe2h2e54y9nisF9GozOGjl2gFRjydf+8uJVGZM+A/ENyc
ET8y0/pjF1n1lQhbb9XnHUiBVdvQJh4romddbxfj+SuglNM7xdcUqnA7s1eT
jPM96HBH27c3NbeS66xs3vpmQUV8qk2Yh2P6nKalMLbiAhb+F1Se1KkF9/67
4CQGkppjdIivsXX+d5/JM8EWrjR/yV9JZcO6ENJLmu+WsvZczsOqXBk2ALmj
4VhRLQENm9KLvHKb86r6wyOwibJ5fTJ/NV+vdw1ZnHffHL3IfLdzvt9bnUQ5
qUErP6/knN5lLLxqpFexfQ01FdCvTfe57hrTBrP5+uk/kh4z+hYeuN5Ro3m9
qTuz29zAdk+JMKZHm+k3wuBGNcamMV62xHstpbyX5ax/9EzwMeYB7ee1EBCL
dgOaor7+Refx9EW+fNF+KERs90YiWUHzCK4wqU5Llh8SJgY9GdqOte0GJHVh
+Lrb/E/mLPp7gsMwNRoqfGODY0MUP/tjAnIs89nWd4xuYyUSwFrHX0hA9kJu
RG/9yVMvQp16dCDKVSpABOdxaodL5fLkQQq1VJwE3sv+RzoGlpAdFxHpsXKb
xzpXam/vlp3uFhEz2qIulUNucr2YXhNhdHTRLeEjB5xcqxz7i/JCoME4pbmE
OCM4YL57q2jw63WEnMETOJDM4mpBxi8KOw27MCgOVVFwlReM6daVSH9gN/Dg
FRrVg/dYB65tReJa7LfGRXi92L5+e3j/HqDy0Pecm8u2ErK5nnhYNfdrF4XJ
HGyzHG/+2lbq/a8PTEXR1+mpZ6QD+ZtyDkArGvkhPFCbsBV4soDUzBqAvOJL
ZfDK01eegRzF1qW6d++XbLoKCb2+aebNTQj/crMNQDSU51Y7cGnAcrUpKMUJ
qjjgYvJp3CZUcJVjnZf69lDaAjxfn8pD1awbPqNgxXdlj+3etTlfXU7d26RQ
SBvbk4abDDVCEmnV2wKpUrprBmW3G2pSSA63ffc2FpmmGSkttDfdcRF/0wAg
lZLHEc6nTpjzJnQDK4HAR3NL7IaP0X+flq9IPRrQd8xaQsQm1eXXd/rNOLgm
61x1+9fq/m7HxURYLmLSP3431ckjDPd/YENgaE70DQ9VhQaQa7WRXVWiHp6Z
E+cUNZNh6gS2g0WX9iNromCow4dPsdYgqxGUOYQ8yfz81OYvUTx0/zbAEwcX
zf8zHBDBrv9TfPMqa4HmNPRRfL70NMcb13PufzeQM/m1a/5sGTKCwrhUPq7z
y9ctLfiMb6FaDT4kJkpTf1uCOKpYhVvzM+yGo/ZorCukzEFIBuv+o45gbKok
u/QfQO22ZReblI1eabd3wFYXRFo1TQK9PP+fJQDZW2cj10kNFMVjSDEZkvjP
qEfGDN9gJt5cw+1kAB00cgrDp+EDTgK+SqZ5c3jpsJRXmzeTUiidTZfNwrL9
hRnYzbQEJvykYvQ6wbhqWZYj/w+SSidJwvwHyOePEfDpR23rVPMEmDhUdJY1
dlnc9imjgfIxnkx4x7Gn1NZGfOOiMnP6b3zyHit8o9cTkAg5fBW2eweifXH7
cobZ6AAlDRYrUqrO2x8is5/qcWQvjRMxouQfEPfCDEEc0V2bUk5uzZSbyJC0
1rWTnazvQZq1B+e/N/tQpCYddQVmCWy31GbIYhVZARW2kzVOlJ7V+5EoLo0I
KpqbFiJ/NXdeoLXHcNy6Zj7Mo1bpYH2Jw0mPd1lSUVKWHfWMwuUeqQWZabpa
yETwvD4r7uemKz2vNwDWJ8ciprxW5LwXlGto69f1aSGi+UevQBTcyRKMaw1/
aFxy9r63L76ByIaMEMrox5Wqv5p6gAu3Bl6lB//1Iee09lwHRVP4128fKVyD
zpS5opsscUEyIg+VKnOhY7iDWDqUHeKnuoLSebtSkzJ77U0UdfmIouel19wQ
JsMdVlNp6MklAntUyo1nE4vwlAHgvzruJicZIwh1b8i7OmXHFU1xpom5EQUO
egfu0joy68C7ZAvKBH19KpK4+UnDOvoKy94yArQ/AS0HRlv/y9hLjMFg6v65
M73fxiN0TFUTng+KsP/ofEJJGrVzquKe+udic3NzPjXt3UCOJYkfTAulJriz
aVNN63sHt+Pg4+832i1Iu3YSV3zs23kIuZ3bF4GKtuSB3fnji09ERN8CfXbx
Ty4hWwZNpnP6pWiJLhzD2j2snCNGNTpFpeQJ9cp0zyqsX/+J2+Ps6AF/hkbI
z7SV4KWRVPApzfz49TTGBo4ocfiraouPZJdlI3sMjPuX/AbfvN9FFaArdDmD
m+ZB+74zJWfYdV+2b6iK0+bg0MzutofwLRMY8izAm4TvrivRUMd9MgNGXl0W
XxXU8VuvDSA3McOaOjOXz6FH9O/j6LPjVWyUXw/piP1ux8W3pXqAmdS/sHpg
JvyTCDPwwKFSjcco9GThkKOygVFBSFS0a81+ePOJETZDcAsjJfbMm1up9Qsh
403W+a9c92iemvSdp6grJKumsKuUDmfkTlY0uqKIjkuZz+aeq37aa0d7PEnT
kPASD4EOF/JM8+4UJEmEKrlSV+jCMvCbNHRBeyUzWZO+n9LqKcWi1h3WQCia
FqhcDXjjSiV82JuU7f8izo3UTFqrBJhn1vnwfUT5vcCIH6q+CzkY88SFp6lE
OyZiHOmFHmslCXAr4WZibgggOuhjga3rtGYHbFnuWSZgjgKVJZMmfZ6rVLnh
ZylyvxVXygX8MQ26o300/9Kt3U6mOK9kr9W5G42FByZdFLyPVS7zmhWpnTbB
QPou9WgXTUf2Ce5qLStMsj8fRzRHwC1JUJUe13cV9/9Op1n+b/VAfHKLefuu
pWbcQUm3eaxZmQRuiunpbnwOW0dzDkqqTYeS3Q8P1S/3dtkEB1C8atJ//HXa
DRoifrbNVo5m3yGtriSJ50Ok96YuwZKCx+RW76/LceFG8rMJeuo1sH3UgtPq
C3XxKiEi5CEQdXD031oKBkufH8nOxYVOaAZr37VVTeC46IBQ89D8L7dVqQBt
z1B7SCGH751In7ZFXvB+z+gTV0Dbbxcw2X3lab+VFKaYDbvNSXRYvfwrM/Fx
ocHS5NyZzlyMBcCaRwed/z/9VRvufY0k9kVWYuETPVAsFVtxEOuFuLgZNTe5
FhNFabCXAfqndiYT/vZbTy5h+mR0+NaFbKat5f6ZIZZ8ef4BJ0Ql+GPTNt6L
NIJbYJWofewl+y6bFx/zZqEesAZTfi5eAeiQ2FvczdSSxiFPUhWvZwRP/flV
MRUbCHcanm18s3IQe+UnT5CsJ3mQQehuCN7dxQXASuuNpK/f7ZynQVQrlLk4
xIClQ/NqzWQb4m4S6XUZXK6u2wUt3ZMjYXN19DyNrNucuigIhj+u+Ui4CwV2
ZX+/ubuWyrOgCE1GCbGWDmpIjLrQtqysEEdCnpMM4Gva5ntzpOCPUt0s00CB
WqaGTBjG5ihBGQIwZFf/c4ZUJKziR2OfIEhtRyZ+SOnLW9ghg/iGz+3TPPRv
sMWNk1P7inZF0ae6xn/pDIqmDR+49B+y31NU1QgLW3qoUNjLmnDhcxPm0zCt
/NnP++/z1UdskI5fWRzTaNrlVq0EwXLGDC1YZXlJgua6sKNaCFPSPJV2TX0j
+Jmr9sXr0kp2HG29c5RGM0U5r5L7mElDVxqacqBJ/V/ogryqUrbywrY1gX03
naQHR8che5m+fzS4nu6OIFAh6cHlZtoF929OiE0F1Pk35fIEEEFAYatBBV6F
X0J5AXgYnY9/Anz/HZb0LE3fK3F51qvvoYIqY7j0gUMOQgNem1f5+q/qF7Q7
INmX3T5FUYHlQIoVTt1MCgE+sZeVxU8cqRyOdfTAjsfFOCJRwpppzACrrSYF
aMiXo/L02yghD2xq6ZlwDriZ1v7IM9RRtdjAKz3f5Qij+mA01lCA6kqXIFoc
rANc86qyQlhELddGHCuojSiBWEX4hjKSbxP3nqUAkS4+U6U9HEF8AypUFbX7
N84801YQdkidZ582F95DU2qM/9CUov7yqkZW/k9rF72wlHa+8CLr+iZ1W53E
PfNnjjEdadk0u4sF0f5nGUPMMO7r5PKCdYdesydxAaj3YmDUOcUKyRKYHdKU
/zojsLSAEHQpPtEZG87lPaNlJ+MVN5ZQoWv+MEt4dVkEUNZZhX/oa6855lvK
Pn0NyepnbfxUEdHyCy0b3aPyGuVww0yV+S/Z76jexuEYR+nAmjaYZEZbo00G
4t0ntjkWf9YiZmmGHIxMNNGZ2rZmfy9+XnUcN99u4ODJ5aIZQByNaXZHHi53
Z98Kcqj0W+SHRmO1PiFc28FkKBZtqQrPZ7dSjHFSt1AnLF7T2PxcoBT+6M3D
0VqIrx6ATk61cHhecex/FYyQZ9lPtyR1jGiY2c4Tz6b4pi5smn2VCAmhw9p4
b4ALNqIn6aZuaAXOM7DvStNozJr2NFCMhIxYG35JklgmReGb6GhhaTeaJZ55
Lg23FgblVuI6A6MIMvsWy8TqIKyYOVzzwAw1eLbGEJ7hFyxl3GhBLeNJOPmw
KTNgW/dNgOeqHnfRnDOryVmC+JVNbUzlo8MS/e/lJ7gWeUSepR40lINzfaHy
4iVPXFgc4dGDUb7903A2hHKs7jFloBHR4WS702Hkjhf/v7FFWU6/4AxU0Wsv
nvot3cJx/zZdpxC+n3K+vCyKkYSyujgIFpTIaPI+zd4Z03JPpM8a8GIsp4V3
SGfDlyeXmJSK+YI6eymO33xSsrxp02tDznEMGtVujeYedzzNqer/gKPU8PRk
vKbAfVlanYMvaK9dB/Njt4uV5TdoE6NoNhQxum5ETnuQP4L39KGcd66TKkid
DQcCZ44RSR3axx0q0Sx3Z+dwTRg6p6+eC7O9QE3nxLSImknnxU2CIf+t8eB3
mtWD0z8XZJYMhcSEqclE1W0kfFKg2i/17G/bZy9ZbW6HJ63ptE/uI/gWJI/V
CNqTfJdGXmxIeeGTktUpIluA5CD41FlMOpVjdc833D4aAe3buXiG2Qs+uZK1
0V+kq741VqVUtCw3udsuzbAl5F5YUeMPpg5IDth3GclcaXKGl11I24oPXzQE
hAooabULFQuD3J0AQP2Gt/xh5aKpXiyr2mjtHUJ54DpWWc4Xhe/z/hFKamVj
mfZ2iywvHs5H+wK8Xo8cEH817EZ6Y0ZQj59bfXxi964m22ceYl1DyQLhMUOk
ZgpqCH2V+yD1y+EBiXYHUWNHtZW1ma4MVBnCJjxjbZzMRXmjn0Q1B3iZlE1d
eDK6u29EYtUUZXCwYSwzVfgvY87aXGjGigydDxjgkKFMas0umCOE9Ymp8NUu
ZMN3/5a1aqkuBePUijyHn88kLyaW0jnCdpF9oonZYCtmk26Bsexuk8ojgdD2
KDF+Zw1W87z1Eodl4GuuzZDWWjXqR5PEmM8noFiQEhtj9xlRGKhqXFXVjcWC
+LxVWw3dGPXrBnvD4l9IviDIsifePwPaETOA1NscUGT0Ap28bhaWtqD+mEp0
I8aEmjYtOBDSHUWIvn5PnvaZtUAtmVW/SOXQXIA0C9l9uiEnYxhxOax0W9Z+
Q65ZbV8QtqybwUAYTCXr51qxil+8cTR9oQDuBhzBQSdlk64HRPsHM09U6Rw+
MxqbIEE0kRda58c0mCrh0C3Wvkbo3xem2GvdMF5wENm0USbqAyQ1nqYIOBTM
6Z5Ex1xHdc9xWG8wZafRmCOn7H4w9wWLzuHw2g2MC8lIOe7lzhpAHQMakIFO
50cEqVdA0S7AlGm0/0Ea1XQaznlsR9j9vJ9DLPbzwPcfWyrFIWQavvrSFzS7
+mHw/GT24VNjkY/ad9XgAxy+X/LIjaHC+as/uBaGfNZbx78qlRqIWN2+bCe7
71f1eqeuLK/r7s+qOPYq1kMH8FRO4FhMLNswhHwP6Xpw0759+FP/OqO+yWaf
kGT1+hIIKM3BiL9AxadCjdza8VZ37+BEVuMvSjgTkYHMU59O49el10cMjFga
boB50YJFaQ/1bLNrh5Or+GOMmafYFs4EEyfZDJGfk2+R5BThD3NAMo0ZSt+R
wL3yXIeWJIRXbgR2o4WgOanJlsMlh5NKcgR8D2YTzrkJRn2VSesthZCn70Uo
cO7z81mBj1dnEFTdt2PEtEjARe+nLzA5gKBa5x2TrbN2ZMhrkAWP0LZFdW5V
gwvoo1MeoIXrngGcE9eFOHsbk2FyaSlWN8FMBBTIP+r9a7KsHjSl03HtLdPp
8doXG6g88qBifzHJ8s8sApPurlwd41P06vM9d7zF/ALuHjVVqiZCOcVP+0Ez
+L4iM9XgjBxzY8Vugjn8sMBrIPdjgRa2DwPHlEJnR/ng/Kd14cZa8aZEBweB
3SRDPGl3itP43/F024MVzu1Q1YgoqMhaZvaGV9EqMyV29/vt7MVUkbZm3E0K
hIpZj2SMBskI6TEV9/n0JawDUajpmPzdx247E/eYDW1G2lqvWjLP4BzOGUuS
aSt5R/7wf5pDX5LaRTEQo0AenOEsWCwGtY2+6tO3GbMvTRgcmmyzK5GTeP19
6bk5WThvhi1GlspmEi/QHvb8AXmlSsBDKBS4FxyRU+PbRDPaLEVOq+cAcXBV
ZYJK+xg4MldrrR5/u5UENa+nX0Ry2VNoZ7p5gvxwzY1EczcPWNXo6oS2woRF
uA7psc3602IX6Xctw0IUFtdpE+kOSe1TKelOBBydaoTeLqcfIzoifY8h/LPU
8DOXrGo6kVVGtM64EOCGNjE8qJ5Fd7ZEs0+kW/EaJmnFUDcsDpsIant9fElE
Pb0gMebU6ShrBU8Cn5amnCkPnqUKuLODyatob/q0Vq1bppt3+90/pbhSZggy
Cow4EESbJsfQk7p2wPu+SwrSsJm8FOnlZtdjoa15yyz7EaKC2wzz51XbtkCo
4Qu9rvE8XmSTSfvYfyZyItAYPpFnzFoe39RW1RyJVTKB9MVykZNIn+n6FHS5
DXwMdqzfn7nLdVIEuTuvgEaEzVkP9ze321KzTv3yY0Qo351UY3B+PhCDIVTR
+OR5xxxqFl/HrX6GVlY350KVnQNile1xg2F/qJ8+OG2ePzUUG9yKUNymtQJI
YDgRTh6msqlyGmYBmvv8FDxmOM8TtxWrG3ySinK90K0X6p+4rz1EK0rpEOrN
HsHQekCHlm+Wq9g1JaP4oHlhxMKmIj6qtfOeG3L++4W2VFMJVtjLjdGQPv1h
UtA0bEffvISGLBYldwzqQv3HnlYBTOW7BxAsYHmxSaM3YPf+9oqp/2w324Xd
8UonwrEZW3ITWAjLePhyWYTXnMpjZk4L8YYVd8ovQc6XlyS6HWw65033JRO6
DCHVg9uUzOPnZ/PMWhJ072rBPuYNpVF/BQZCuZTm/VVl6CUT57xbRPjtS5S3
mVDpKUlv6id5YLeJiDoO1jggP6xxpgcRxocEsWKA0klzAZiKbWYaApfjZYpE
a27JH9yfpHL8toRkbj5OiC+72eG6TBCcqPO0LPP44c1Fe4xbrbMLEhywtkOq
9sakvKM9IYxSBDMkowBHo5r7kdB6jvGwrrb0BbH0W6EATzqrDR3z8OXxFAyW
hkcrYldoSvgy2/flJFMokcDA0B3/FzpmKD6iGcYIeloC6tTwaUhzqXKhYIN0
PFp/FMBzJbdbETGuq62JLvFgEW4HN0pF932BA5hP18BlQiikwpbsk3MYCNsB
lqATSFSyrV9X1qsXL+9tqh+kAIkBh3QkvukhEdCf+Gm1vtPnHJwDt53hmMQ7
1OtQZYq7Al0QxglHjp0KHU4GTz/iiCYTQ2T9cILDRA9bQ158Sfd0QpNa2DGE
c3KHw56dpCff5eMON9rSRULUsFWvKH8KRAV1MI87SK7eFTxm46w+5cQ2GMrv
ZXY6Pv/8vZJ2WGWxXohRVQ+68HXP7tiwW6Tx/ZMqaOiEtSA3MqqCJbZs+0+h
tG1Nbr929pIyeCpQ0TkDUNflXE0B7swN3rdkfAyQ26XkQR/rpTRNsrigrWpM
U+ztEo4IqV4wcXP5hfDIWTZUTwc1QaAd5ax+kVwjDsUjezepWTDGWgUc7yoj
ed7B61OLPcjA+BHx3fLOciufSkmbUJZMxXlfRbJ/7xIOIQk7piNudwGnLKCl
iknGtxPNQnBVKKv3Y2quXS0J3xJWtWvtyWHUbbO5cuBNpPNbW9z+cMY6SRc1
z+JSyRaHlRVmO2BhcRfrm3pqPJk8HYEsaOzqCn7kb5SVEOczuIiY75G6fTPX
he0R6LuGePPf+sjzRp16r47C0xaSWHPh8DODaH7FHPrteHdJlTsVLJh8JNrW
q02IZC+1TeNYhBUj9XWYBjcJIFXgqiIm5RfhiK9H4yOiU7+SzNxLvY7wiUAU
ycyban3QuzAurfWMJl5n/4lSxofmS5nFocDwGM0IWDz0kszUWGCJ237o33d5
uGfFO6JHY11mOiVeUhqwgOo98pK13Cs8TFEHUO2Kqou3paL4BFjHDQDqnZhY
ATgMhRGXkDQEDdsmlGgvz+kNVO6NXSmGDYx4QWj5y9YT1fjgUAw1YvgE+CvR
I1QlkhAoRmvjGtMguOOIpidBiSSbaCwyryItUAM/mrPG0+oDK/UKXwdYuSeu
zdnYJj6RgGE1arGFPvMm3FXu5I239fXMRX80prbRkSLlZNgdkW/MVuVYo5cq
PNhNJ+YcBE80B7F1onRcim9gOHkIflmWgGNvCC9355FzYtvKN9WeylDVzB6p
2pPtjIi43Qe4cqB8BOsq0ZBjmbPSNfQdHAROtDPdKyqLVhCsMhyPI8wTolp9
5ZBRXtDwHoM6Z5lz7zuodhKYh9C6tErTXjh2QXhyWXiJuKN28GdU0L2YuqF4
f7moxU/Mu0WDPkEIiRfOBP2kq0B+pcdImekT8eTsSFGyQA241NR2KOTQlJ+/
O5LgN7LWVLY3WeVnpNvvYjg1jW/r9Jlt8PdpkErxl3oKMWl9evu3/m9XChOT
1aE3S05qypZWBHuZs4sa6cWcALgOtsOqUqCw5PSMUqGjbCEYfpqfIDxkV52T
IgTmN3R0f1Lj4Ev6JFxoz61P/cRdhZdDFySbOBgSZqdwMIngOT3ASHTfCXvl
xF/Hdyuezgf+r/ym2vyfg61f3aaRqnRxHir7N/XjyGk9cHIdlT4dfOOo7SJE
vVc+WQIxt5GP6b77ufuIV6OJfcRDI/dvynynC2UDatALPy297bzLT7YnePz0
bh7B/+N1r1CECm21RlaRcD8jUiw0qWE246LuTz2Z3V7XBiNQpIiGbnCKeWhV
DTi1RPiW3Q158x6wr7RPpzB2HLCObcnXvKvswyHHeIRNng05bpRAkm/EWKE4
rl08D+NIlbE7rgizBGcEId58aLJqsMjsyPVc6xnRQBZWcPEhDnfpxJQkYqcr
heZUO5rUp1p1aa6a6llBsDps+gEL13ttXQBMfJzmDNj8WB5r2SfgNPk31NPX
8uUIeWIjB9OmkVLBFRg6TEQAo/+Jacc0WR5FYfWEGl1Vqrqvh0RJhC6XroV2
U+JJj1ujUxZnXVB/gPlIUuv4df5q0Krfb3Tz6wd5T1QST+8jD2Jz839nh5LZ
X+RjDelAcSLhZvp1bQggAL3VYp6kpmYFP+L8OA4vcAghUI9wx0k0XLTNa7gL
AOjhObWG2I7VA5kLoYa+v0lLqE3C2dLVBz9ipQj6/VQyDpcbrmZSMxJTcbsU
qNfskJVYxdMASSWosqnZWy/jFvHqD6PbI15MYxzKQpVmZ2L6zcxTZ2+yIVij
xnUlFqgPndiCPHnPR8hy3nyUIFdfdcfqz4Eqm21+7A5fdO7L1pjKcMxuueGq
439VhUx84JdapegUA5dJBsn7rg+ltMTimmcVHtDrgUXjQYbZT4DJDdFfpatt
0pC5b6XJHJkQvFO40VtTuRgwp5BvIbtbsMcNUjom19P3Eer2SvQdstuIirN6
8e1WSOc98k4ya2DCVVNtNk4XRhomtvXihRep8n07HhBgExrn7QgCKrFac6jS
EclMhUdbnEnoKihT/QY5mlYsdNvyqPkPARJqJ3Ni1A9QGhxS0JBqzxpGmjc+
lgsBI8LWDfwDyU/T5UPAdYeqfjiVV1b/vtaCsQjCpT3TxCY8MiacCT9bTllw
cpHCo1GHNgF3d6JlAQJXhXkyG1Ae5g2LiBAYrty4F6FSjCkr5Cvlpxc6H0uc
gvs+XVvGk/jTFjP+YSxDIKmwLgej4S4il1hc5JXA0yiLxtuS7UO8+R4EPKYO
wurlcvOjkISod3pp73MY3W/ucxXU6uDgtKWOmPRxZ+vtIN/45L+lyFTLSQz0
JcTEI/FQ5NNn3kew84sGShAGzoKlJw+3XyfYkPJBTm2zDlIiaUq08cafID++
AO666kxU6mdJL2exSiNf7ypLGs2g3apxDbs9TSeh/ALpZKHXLC6AezALzx8T
JR7WD2LFnnhw5Xs7ZLC2P3yOOOab0K9iV0IoZwRP+J3pl3fQCE8aJA2y+Dd6
N5hHfIKS6bD4GySd0a9UhVbsa6kyD93XUtUMPwTozCWP0rpgVHuymT1wZV6h
bZVkyXGolE38qL8yAFywd7SEJZNhsOQLCxxX27wISsJ6Eh2vt3/lzgRnAGPH
5ASllFSfbsUZ50XozQVEVFFnP1A6SLfQWJ3NTNpT/QIis4olvftk/gEVF9kq
W8ym40v+ar6DNJK9XZpcDM4sXVG8y6vz8OKDPTo7zI6JhPfUdZY/u4bNPrGC
4QeV3nJhVYdhV4u8wREdqJw/wWKuEk0wP3fDkQ+2vKmT46KMdY1PFg3o1gUS
yNT7cb0nMAZL7yeJ7RyoYZMyebkpErr3aFRHds8BQT3x8lHwhkOu+DuWdWJ4
/4esoAFb20wSo/D0zFzvjZ9bB/pNLomozhmFOOZc0pXDwLzJsgGr1NaXupwZ
+1umIh0YMgGvjdUAbdOhqM3hrr2IyPs9HeOndqm2CLQEdyA5F83VvxRierK7
/CwbWkAnRk7pzrbBzN6sYxOfOnc85/voqUfmPpyXZKmpQyW+xpAHsr/K74qc
s2y+NgSz89cKV0qlU5tFr+YBnN7ELRXMYHSnQ3QTc4EsJEBvYMaZJ2zv4aBv
qiYP6O7P50jI3bAr9ndzB/LdF+8mEhxsVIGkYkLTfwx6WpClVPBxOEW7nWLe
vVffnN38tMvgXtgzaCEHukdZDDyPCph0yGlu3rEME6n7Bsj/NOyWW8KUCxrC
nrJDMEkkOIigJMArYFE50dqJh50RuhXFC32heuO3TpsySPxC4UltcAkKLLRf
4DmogHrebyjuiEZ2mpYzXBRfCKEb3sW6bcLR7jCtyI6d+H7ia1X1S9v0rJdH
x0Dpkfy5zpaLkqvCRvUfX1S4j+rRrvKdw5e3GzHjkIDwOzV+tlLx9ljOkF55
TT8zK6AQOTswKcHSt9ltHKXtRzr5o2FQ89yv1zZeOoxSC/md4M/trXi+sUyK
UJgpVT+cqS2oc9y0RBGu3o/iq03E6frfwc6I+k3E4IFLI8NVP3uN7jHyJ1ir
b9dysjCaB3Ee0zBCfImB+110K/pmsD+NOngEQBOo6u6U3ynO2PfMUOU8W4yE
NyeHqXwG4/QGlOeqeCG6/DurxO1tqiveQ9OMpq7On9Z03rWwOHHhcrd909Vr
pUvXAvRdDAbMYrXGFka12/jBgbBGfMiUvF3HpA66tZKEgywqz23B2/kqhkF8
2qkikAPx/4f0VpMO7hGIMLakhlwOQYq5ibxYtTAJ8wOt+VKyqUriCBCiUlcb
JKqs0M2JIMOS1yFFSCQGMFnQcVItYqZezeo2O2/IMOh1X4f5tSQSukJRXpKQ
mjRBPeTMsCAjGxlS0VuvaFkwZxYsctqqSFiZYsUsQ0Snuzb23JOHgC74fjPR
+NSIHaXCDKwdnFBHzat1CJiS0wtW5rxXGE1t+HHRFaIljEl5hFztaW7Wr1N/
u76uKn/qRXc2qJ/7tshgK/AZZIaBC+ozN9PdxYrPwDe/XNEkyAWeeTr0g5FO
ZR4N+HluB0esZLygjG1RSPwE4JejD6GqcNkKdUTX9ivm773NRMs6p5aF9BSQ
gmVYBkg/FB10gHcDu5OoYuzt2CnOHd9e74i8PRNTICQRZ/9f8HIGEuGlNCWu
7RYDuuAPgkCF2DcKdOkpWqyPeXMUVNSRZi6HQnYBAEei61hoYj7jIwlfWqYu
j3vV7XthINrawRmwndKAO5eYw/Hxc1U8HkhafunFCU7QYr7uAXBIFVNyl/2u
zmU/Z9dgLcHJFQXpwxgYxQEYcPNP8j3ndAs0Xrrhmex/CSXOqCZAGtJLzOyj
+N8mQpoRBKy+t8kprCa+SbNhNQ2GzdoNbg3QKfLwdFBxk7tAB+Z4aui8LDDF
4h6s9q2THmXDyu7v1NQZH6ZmBOt3TqkKQ9v5Gf0GCjHA7uLTut6U3GPr3n5C
H86OMTJqd1H+lgJr/8IojyGVawZEiB5enm1fvCrDs4NNvdp32IGpfN+zQSIt
8RXdhZFU/6U8coju+bZMVd9x5eMfEQulK5H8ds9uklGfnrwLTUA65gBI+6vD
XHai4xHgsY/lcE287Y81Uu8iXeUdcKT4ZsQ63ZgRBNowleNgZfUAiTqutpfJ
eeS+dUvyEBRfT2w+bKLjZaGLdbEoa3Py2UrmaAWgz/XcggbNMMx3tK6q+rps
pZbrWYUTjgz4B/Ut/dbB6SiqpFSvWmq6KApBXOfs/TiyxzqSiT+e3fIWzzA5
z54Jm7cRvg65UcVNon6pPfzbV1wjo+5+C9NXx6Z738Rdo29q6Q5bV965e7oq
IuNvYe4gf2tN2BHDAUFwTVtRvCJqtUrbcnxsH9V/6e1GMQ8TCIN++98zRMKq
nR2b+inGoGpY+NGrzmkA3uttmNCYkNnqCy0tqYcYKkuQEw3u1V18k82DmRZt
dm5wLqH3d93TpRqvL5wkTXl6pdCAW7YBlhXTy+sFfNtgRIvTUBU07bJtlRLb
G7puj6xxmn67q7yc+j6XnZbdomdUYa0g7tqNSB3A6gUdDqHRTXsb+hI6G4+C
jntQ/XBGoc+k5Lxar8Q9NzKBeB5jfSAnU4yPyINvsz3Ntu+TNfpv1hrnnkWO
wcKLYSNaAr1cB8fFrHJS1wU/WtmhZgeQwov97vA8PqGneVJ93vvhTKJ9V50b
BKH7TEeOSzq2e6vHnCktA8mkF8TycBqawu7w1k/3j8dZVwgvxt32Te1XHdvt
KdKplHMAv6Go0YGat9184zCr8VdiSzeXj+BMjwEihhks4I6oB+ulbwqR5oy1
xTdM/aBx7tsBN8rAyKfcLn1UYSGGqtcl3xpBRttNNPigv6qxldKWBiZLijLy
p3zdamOoz400xAh6BuuP5NTvBg0otIRnwVhpt+xHgtkdGYk54nTP7Hm0IuG6
sU3AnY6opw5Rkh6uZzBxlpMtCrT0728mMtGtWllMhbzDLG304vSXZYEuyCMw
Fk3vBcT2Wz7s6D7XQvguyw6g1VtW4JrN/4LIuA9YvkmdGBelmQ6zZRymSQVj
QE7h98mTDjc6phHrpfKBio6jd5krcB7GvQXpJPJTDKRUyvKynWoCvXZujUyb
U0/4iukmz+RP0kLr8xz+X/0KaBL5j5R+F4IuXo+hgkGMkOYhCWV9gsew/qKv
O11Ylpl3sada+dlcJjb3SSPRkaUZCDIt66RQIUbrB78+pfHwveN7GK4wxIi7
m3TrDd8is4qT7YI3NNPov7oxi4YWA2GTyRg3M0YazNTJ+DKD4Ug54OhBHAoj
+afzbhvWf0VoIAzS7LrrQ93vd0PcYZvFE55CyxBFqQ1oeSiSHfyZxd/51z0r
vFPYkGi1RmPtbKmcSRE6yFjXo8949HfXhwp4oglQul66iKxZsUk6eHSibGLD
ll+//Z2dIFXdY1/xDc+UPUhjQPeZKwZVOxVz+uQFyX68JW6aLc1Cr6LmN41y
iG4+TacERegKvNEbb12IyssCamawlnzUgj15Ldd3Owi0hLTKXs09hL46aYWM
OIuUVHBrFX2pSYKqDT3MVisntULkMF8JiyJHLkPGaDboPVPFb+jSmFs3diVm
XOaYHBWG2ydcUsMmFsUY9roNx/bGzgEHSODo70Qz8bDf5wHWkTHfogtwJyfw
jCyEc51XyNYjgdx416Hcu/UaHfRoiPuZ48zrZ29zluQBfIbr33UGUWPV/RMs
Yj9Dpomg5yNr4MoC+HTWg62M3aNGBkBcJyqUrP2+wpWvOqDCpadCA9NkatyD
E0EQjTrytpJhL0xbWoLKCRYl9ostyIeiZEimcfsxtF3pu7sh8+JxGZXecLjr
m1BUjT4lKP4w8v1z0oehRLE/4hTa3tFOwWm+TeQpwHfUwLV0hg8VuMfKuf/U
pIB/TE+E6/M8EcwvbkfaxRrt7XKU9J4w61WP/y3co0d4aA7wnl+JUbh2ZROp
PhIosAFPRw0tM0JvHNoP5ohL88JV2tzsVjYkpo142oDmPGf8SEsYJiNXb13a
jk+dobbFwL51H7/5zeuFpg5wrHHZn4x6hUi2rHxUxImM/UKt+9zxqUotmSlD
nws5FBGQgtT9u8ODOEuTxW42HF2p8DBBd8gWUTt+0sjYDcPU8Z5XOUSJcHP+
WneVnH8A0kLDmv3iRixVTJST1jG95xQzFlY4OKbF/anmTYVjvtUwHCtisNRI
vuMD7Fohw2VEA/lbn0obwuTdWup3p6qjOp1oot4n0VAe128+lkos1hqBWiUe
VPYfeSbyhDDHYrTQryLTE/KnLUrcZ0mGGZ0XYhflH1mfYyih1l/xCEA7G5Fg
NJG2KzVQJ9mzE1n/nyUNVWgCmQETopLE95KGh0vZ2jxGTNZ8s/8g1smVZqQ2
S8X2UL6HeuQcUd/LknKQVHMjGzl0eNHzxtnp9IqUUuYwlVhEQ8s6SD4Hw1rR
IFRZgmECxqEA9mcBQHA3ObN5gfz/uglmgD1mR6e7+yMoFzwKhbbXkaj2kP2K
IqfAl2WWczH9GLrbC3XI7+6GbmXGyXxJqWl5CbHr/lAb+D5zrswMcjHj6WiL
5n0ISSK0dCi3H+T2L2gdvHrbc7bmLFac7KC7ueY4rvN1zsjdXpDBMJaqFOWj
wp7KeuixSGJPOu5KGCkggu6MlsYcDX8CfRxWF9whpbOjDToDnJwKVpH8O5Rg
aH8WnrTcvLQXJxQBKbftITLkudqPz9gNKbhDpS4SKw+aD8z/iwEBi+CiJBt7
WELg4nmwzbdpE0yOx98gIveBJ8pZqIzmofaD7r+Z9ChBUnO3zw0s9Exu14sN
2OoOt35nnDVm80r5vmrB/jQH+f6wdjsVcgBToZq6DNvysfDiKkyoumggJ5pz
PH+/10kJHC1zl9FDoNbG6BwFCLzg2+5tNKQdAsDbAYx4llpPLhRAk7r01x7D
jw8ceDtxr+AA8gghnA8+fCM7yiI6abBUIcDMlzFJgFnkxQpZBYko4qzsvrC7
FI3wxygbsFIdksZIJZBITIo53ptKwsagMO/NuwRw9O/aKTXkzPp0vhQZS1Nm
zg2lRuI73OgK9xMk3kL8L01omdSmYsfUHK85VMJatg9g7RacWhYTzoGvVkKJ
B2COaiFmbzqrD6Kvee0jO5/hInRDclYEBa3at3iSZamTFoi0PVb6sPVEeBLW
XSIhOZMjI4OSs3aVa7aPhD5d6/yHnN57A0+/B//H7Kuzmxf/X5wxNUcMe8h8
S8FVMzgbbkvCs6opuZBkDoi5b2TYzc4/6GTX7nocwXCYhd0Jr/bQFB30Z9aX
3xcw3WZyNvTdT/t8g+A3PbkVuwL1SZdGtPVMU9kX4mAOPKwB9EX6Jw3p/qJS
TAWy+VOkIPc4RJHyW4e3l8h30Q6TK5tB5rbEdrtjwtYrgCYDvD+bb8MNQPF7
gRC+VZUyFOX9PY55D7QsGHDWnvx1nrOZwlrYAwtODUu2jGycoPxql/E7zZuX
bro5ZkiTek+IgWbEjTUok9ga7QTY3BT27nW1wlh1OVfTQC5eTMEzamtvuPv3
3YJ4MTjkMvEqGa488/3iCuXzdvgD49JNBUZAdwyOG+QGy7PTvBsiuprOORVI
LRncxbB841r/T1Ok7NmhoxjyFxiCQcx3YhpaFFZA5vvqvDiRyj0w44b4WEC9
kyH+ZyUIFKUkjUPvV8THNpdLREVXvXP4bKCc4Y/UZ0Ilbg+PLpPRMqgL+dA3
vVAzh3Ci9nLbREOlbW4tlzvIBUyCuckwfy9+8NDh9CcQ2FupaP6c1rWQcUDf
SSrI0pEd38jSJF00cGaIA9cxtC21yCZmLJybi74cNIw3U6pbMz+jywg4lxym
ez5Kiiyq+g0qZ7g2E2ulS2zKhxaP8jGLsTMGCfBjmF8VmOyCFEmjY63rNtiS
SQcgeOeLMzxGyWUzZcN8CWwUfdguAtyXnQzcKhM/OMOnSXnZwAEaY8sHhF2i
opBpWWPzy2pPd4KPVunuREAZ8WAfUloqRhWRWQK7buyAWLGuVdCHj2i9Phll
WsfswA+78Z9wQ2bPw8LPDPA5aowInFfiQNYCTSeKPQuq9lM9iT75qJ/ciWUd
erAkvNXZz86mD4vfv/+I8DlsPVZfidsRynpmOQZ9zUCX5fDOE5kf09AH5FyM
KDQMDgSkmQi+B2xi/VpKCyicOaDknLIASyzrKSjZ5JJwuzMZzP9xqWBVOKBK
F/e0Y2k5Gn66FzXxwzSwlN0iUkK7m3HcSS1kfxbGfCSVLnnobVuvaODIBE7O
oOWy0/3cxjAznAA61uQ6UdsYdp7/eXZIpnMzdbRNNZ4rC0345QHEVWiUZHUs
39T80DJlpt1EueqMRyUMYWf3LyDEepi4ADTjnQfH9+3rXncTUkCPnIz7em3Y
gb0Czr8sBhULA+M+WN3R+/ZABtspeME/IlP070B4yXR7zbQkY2iVeplP9QMJ
WVqH7TagkHbPWXwbDhMbPljtV8D25STdI1aeV2d+dR+XpEsVCyqbpF1HNHvR
vC3OyUKl2FYVShzE79ik2ZHVy3Jggud64aay+WSSIKHSwqmfIK/GMMI90tnM
lgu0KnQ7hcnpt25kcO5KJuo40HXUCzkoqdeCUmqyjuhrAOeaZkRcRPlcU3H3
MPgyHR9v6eW7zoXmf1u01ahYLtKF4cxRzF4FQBWTEsOKFeG89HxLDAQeROHh
qx0YFcscwSl5u53RVcEvqEpcUpnEoroJ2ZiIQKZ0WJzIetE881lUIZieZc2O
B46xdN2oOaWf9wpARg0FlyZQdvCqrPiWzh6QxIBWUoVPG+TjgxtZZLUg6MWl
HSmd0lynmxsaVUDrrCa29f7ONXFY8rhyTLad1pTxfo+ULcexJS3afVSePwSp
j/LlQC+ZFnkwzzkzaiyytQZXi+90/4g7fim1y+iW/nfHDiU2gDoWrmLggXYJ
C/j2bWudj28KCwGiKg8N8wW6V/z5hKS44bwHY2DFOYcUiHhlkud6WhNxmBCf
3I59nJ5snhZFMoZODySK8yDO3rHz75H1xQ3ksZRcLDd9Ebx3+Q7aLKY8a74U
FgdXNzLd2dYEeeP0O3IuWw49UlQ2gQaUUh8bUjaTZtzSakjRQRUMnCn4tTal
NZvOIy/4k0RkSGBERHnp0R4ajNjCC0gCkT08t7+GWqzUUX/x3zQ45/AQDgLJ
2DRiDpmc4oA5b/Ze7iKS02DWo7MiHJjIiM5gy/p/2Hy1uruqfgdh1/iswqC3
a1EK40pk5E8D34hwVevTByd25uiI5thdnZew/LKveXEJ2DzIqyceXXjOeQu5
axMjNT519EsayCgD2xt76bVdN79J/ZitgEA5AS2me7OIuXMm+tuFVWiNLkWY
Idq8/LWHfH4oTnvawtn4MIQakYwrBCiZf2B3RqQ/FYaddolmf43qh3hlMoV2
GH2Eq+F5FIcQRQIaErHRARVN7TXdFsu/Nq3HW/rv0yABFxa66y0nf5s8xzSa
FF6mVopwNpySNlUOD2nsOkiQE0vcpSH85e2GAWOf7Ceywbo4FZHB61zCPRlG
YQqUR1a1sX9chrpRQXdiUakEPyHWum0/IEWnyZR0Zylf7+OzVZqMoteX+28N
NRCUS0J6VbAx+UYDoQOyOdfX57ua0fNYN4Ro0jiGqIoMPhlc+hJg+MI5Vd69
vUcn4E/F8IKI/20Azc8TZvTMELi0XlkYSwT6h8ww5RSLOBFSMy5AvthWhV/H
b4NXR2a6s5yUBsFP4g2rYltmyZDx+WU+mLVeMDqVKMPuynW5j04CC2RRQI2z
qDZISJqAIF/xS0ceMu4jZBTVI07kN2XD13BVdklHYQvRlDkwqrlaUHWtXHLR
btitlGj9kd8hq1zVCqF4oINQGONeJK+wssZbyEzouJe+dxE9iGrSPPu1iaSe
LygQ/rDcCWAq6TPKM7ENoOHm98SBmoFakY2HgrjW8usYUR3KRzbTz9Nm3PK+
nrjgK9HIfiTs0L3tKzxAKitIezI0d0ngqjN/sywWuFwqnomAnnL2zPIoKUBL
YfuoKuw4rCK59sGeg7rvY3uyeZLCdTdmRw0GCsbaDY33Hm80BOYFOIwCV3/W
xZt+MrBLfh+0f0Go9wv6bL/Ojl1mprPaD7kk3ICyuCSg4kb8WiqyYJrUt06Z
x4LWyQaOobw1FzcMScs8+xzycQSN/Jz1tyj44EHqrSCr1xgqjuGat3xD2/Uq
nwoY3CiiJDTRcU5OR4Jb+1Mu1GjvhINstoDXVHVQOi6yjwIoTFQleeRd1oUB
e8DKpj1S1zwxyqyH+xYlm/2Gq1Yx9XdA8L1ClIugiFea8wxnJfkzH1jVUhCS
feZct0hvA0Ma9af3jx47gw6qOYSkVyfGXTlRSITO7+EIzx1bjrFxrPf6WaXM
b+MiZeNGzCxdo3mpNseH9ohsrGKfNhEwbz3joLZ5MAlQS1hmcM7sTedaSFGD
txaEUNYdrxwhMjs/cijGJcEwdqlO1tZl1TqqptEsISXpO+zXrV5KABQfoCIk
8ZSzOZayqihisCdyIbE5hz65nMr4/n98YpjCqeIATy10NBMxBv5lZ4gs06Dm
SS6w5+s3+R/hz4NIkdkuylEqcyCv1cfqphQF2wDCbl+ttCCHpuaQdECAAVux
WYVcuO1qLbDwGYLBW+IzvEAVAfJZ2W9yKtHmltMFsUujE6cJORhET2AfJTrH
Rdlv4bjUsH8dVyshppNK0srtTms9x3YFq560s92Tll6aUjJ+IdigEBbvmOXB
cv2PvXq5D8Qd3Xb21XS0xr9f29J5mQwhTRn8R/xy5iMXKgz2jg9HSAvfVinV
kxloaWoTaE1rg5nQOZGU0ePwIqQnIR0TzVPH55v1/Qy73ZxIyIVryYj2M4VO
M6Ocs7qay8j6Tl8knrhUlrQdFz6O7CBzRXsnOC869+mS1Jx9zmqtnt7N0Rss
iBwXT3YDGOYpshIZU10lL/VDqgH+3/4n8+PlPC3YxMpLmURPPm7k6yy8O94+
cpWhg2v/d+2Xh0YUqe1quqC+MKvoCNa2SG1WbV7NNTCNLl0r/lRlRU5avHvP
bKn9Pp7rRmbLeLCsp8bzSO+MaAL1wwML5EPUysDCXsWtvDCAgUU6rHB8iwSM
ZhPYNZGAm+vA9wm7WC/wm8gIzToElmkzbfJ1dWS1cO+emKsCF3mDhKOwlpuR
AaoZeRYjnrU8lzN88KPuqgE5IUumd30qpqfhwBBvhzAo8T/FdfuobPj4fXRR
3ucxUaUoGmdSiQzxS8tVgOHrzvtkMdg1auCMs4yT7W2BWpaixox0+MaXp2N8
L9HLPZ0XDzjE5JrRsnEnsGkPODEhTjXN4meVzYOCBtf9aSJ2SChnB6Q8KzeT
DFd22DDUj75f6ebwC+Zv+jd70GUeNNq54gV75LKcKN/Qx4T0uQaHgQ7WN59I
tnUlrNddEruCs8ZAIX+ZwkSMnkWwzJx1cD+mlq1uKNR4m6Y4PMGnbA4l0UUn
OW+HD9XODnI19AqsgHZtkPxBbwViKopmPWTjqzl3CVsVS/8r1q/FcAqN9/ih
457U08MTuFVmD4TRIlpUAEY5VPNnRWb/UXX4bJONLpExkIGaxu6z+aSjCNgO
vykerlwhlmqrn7tjdFYCTSrGm1c0rHRhKbXchczlZR+v3G4pSJ8qsv3mO3Mz
4pUL1EawC8B9oV25cUUKQUoEHYr3G9McyqJ57Fzw+OjMWGjt8M4M06zd6yKw
84aeKYLo5Pg9OGKLqTIWrWJ18uKYveUi0Sx0oKExvap0RHBoKGGL0MRTjoR2
Kzb1pZYfMIOIwHQ+aevcqcnd4CLmuiHzKuUHL8niT1aJXDnSEJvb7C7HF5hN
XTkiHS3Qa+8zkheTKvnz8CDLwAu5oxdKOJmqUdEDwt5qmoLDpz5QS04QS4ee
DGYHJGQnOc6Y2hF5LHQPfqCRmusPedX6Re0cJW836DP9+9A2ZEg70Ji0flXl
VlxV3Vke/jlo4W6cTkj0RBJ6mRifggwfKJNhhv1SA8xNqsmmsm8IqRns7pEi
rf03JYUP+b3nq0etOCnuY8H2qZ+zHlmDicBdInf0CzubXdcIyOEh9u3f6uhe
goTKj2Az3zqILpgjDkA48E4kg4bGz33d8umIplwOcgS9ZJ3xP2MsbEbXW51/
I8aUbejYHoZtzk3M3qfz21q0oG/1RH/xvUugKmgS34jhtBwfU2EBswsmyGlV
F6u8EAlcB693GT8xLfrJBoLlcbpSqVHTow7kR2NaX7LLA5A+TTglKGM1Iftg
fkDK96nOgKBiGdkTAbQPV42ALEvrm6zcsmE+1jZDzv4tc5TbCPD2Rwm9iunT
gqzwpFx9QIL1CafsvjZVn1rjmXmuLbraag5e75bCw85spTvev6CD7V+iyKyB
6WM2qgQnn9AY+JHVEddp2OilacOAbhaLPAOPSm6F+HovQ/C1iwtkhtarQ0I0
UHhqnNkBs2pmFkOiixyTet7glZCNQh+miNuqRa+K5KDu75+wxXGbDYAaXdHQ
tGkBWh5TBgQ3B+rEIMJPDZDB0TtMt0aRiogq09gLPjA+kydTGrLl+a/2ycJs
dfRdSrKzT20SkG2/hwx0AUG898/vfNgzJbt5rY9tXDm0d4e7zfqv/h2Ve2QH
/64g0OfKlCgqztX/KUAhKNYwJZZn1mlI44jHtu0hPG3ppCrm8pqzN0WOL5S7
8KY3Kv/IM5T+DVGkZdAaWkcuxlz8n7m1IApfPyWEBRn1E9BhCVrNIA6Va6F9
vyY7afpaVNElRtLB/7gSrYj4Dgtdczumk+9E1pCjwoIXjVmGLZZ8dNwLuWPf
NafKscCCCUOsim8oF+lIp7IpRcZ3Itn4d7u3Y/sqXFergldmNDT3mvE1m+tY
PzT0mlQW3w109afO1EZ2fxQNfO3kwUgDd2lg1CW742wmXSJD/OBSnH+qOY0j
eT4EduLVLVUy1KCoN1Oa3uQFDIfYuwcsOpxVksNB12fLGqL+kMpNh4N9Jb6R
vEy5joyhTNSs/3jQ4J8Hxc4vRu9KjbCioJophYLM8wwXAlNwe8t2kjEcXecB
9ybePTm7All3ZTx5DvdYI8ZCWUNfqdvz0TmQhWegM3NQJ0Kw2FO1ikkpcnu5
WA2lSDWICCRWl2j9/QyKz81d7nztizZceq+gNf664WnfqQNIEwVCty8mrz1Q
NpeXIM6LKI1YSkHva7JcwdjAxfX2QNs0NupKQvOs5BvwbteEcFwIO5anjrVv
xaQ5JXUfZ1ETZkDwhwprR16JRGcGsgB5+PzqzhZVX8O9/Okent6SvlGep0h7
j5vkjGlzhSCeWjKbyJ7bm8RVOWRWtGg5VVnf7DjnPx97EOcvpiJ5Y7gUW5ir
8FQNijA1aPp4XETcvijHhkfQhxlit6OdcfTFHWvaQK2h03InBJ0e7Yt2a2d7
lLsWYSADVIRavwKzN/nvaVWKnIIcOawTUB8jVqNE8jVc813HxdSigJNQakuN
TVWDh31587gshn96pHHuOnqPOxZrHrSnlUu/0hYjG0ql7eNrl7QWUDu4LN+b
tg5JoamhKtGD8xaBS5x1RyF3C+lR/PY7cMfcTtsAKIXVJQUG8F81+3tLDt6Y
NETH7VX9W+thVXblCGD0zKPuHWLLiYAwnGXDR4IY3uEpI9Yw2KMpdbW8hWtH
5lI8168nMrsXmaJBGpwJnIiAJFDO0hiP5uV32Mw0uEqVkoyeC8C4IZ/u+Yq0
ExjZ0FpAKtNIbkFkVVBvBeQb8HUI7HCg5OWN0tpfDF+7kUKx2c9bso0FARFo
yttQ8l00+yyU6rO/GsBiGV9aGrsslFNIjubjgMKdLdgHZQCd35ixGF93Ixs9
YID+1+u2TnJeJNT+kLus0CI2c3LP5LnLVZxlwDAeAuYyS5XuTS9J43bxVB2V
I6upx+5AK422ob/JdASr8L9bwxYV62YeLatCTBKcZ3C5S7tOphwlyfmXWgX8
3UmfPKYmGYcDJ7jcbmYkUaVl4FmnI4RQELiLdaMUQPg=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyKjGRvIjWHcUKmptrJ+QJi8deR/ckIbOwmo/kzr695yc6Km9dk+03+8g0GwyPfAeixlYdZ/J+9LKuca026e1SuDfRwHHNq2ggfuPcTjpztZyCoNHRZ2+2/tN6U+oX+7d78lP+Z9wsjE4/cLxCIgJGKP6lPPoZXJIBG0ZQZ17NFutNcPvfibzc4chQDiqHl2PnxXtpb4ECzeWk8eTUvaOrw16TGemTLE+0N0+ecVeU744nuWobEdcPeucDJRJk1ERuma1AGIhBdLU7sjZ+lstaFs1oM58YhCM2c0+5szEkeZe6z71aOZy6dgHBE8PzGqRLqvqTtyUJPmLIXUa3J31pr9bajpSHqBykA49flXTD/atjvgxX8CTX39Ss6YUskgI9yJ7qggeKKkYGjeYSLxhQ4U2NQsdnTmTwfsP2NNNZOBCbEg8cuo4HnoLUqPZ5ZqdVJzu0gdZ2UFwy9slwSfhDSLNKG3z+yD4cNCNWOsrp6rRa72H/9MFAB9G4LqEGo88FxMOT2FKkERj+iO2dL+2jyzmunKAI3onK0PFzP6yms9wnOo+7Oqgiz4gYVz7vwrqArjtkD8xgbo3vRAIQocD9f/ZRUw5PqKbCm0J7t0h+RFHcBYUIFDwxYzv5hfehMpG5hV0J/bdNDexkUgMrI6N6d1e0QMXKuWQQGBQ+sG2K0r4oqwHssGeEas/6N4gqFFsLSxT3rYg0dONitX/7iZQZxAkogCXxs5mz+BAX3q9RLrcLdUkkGABwHIsXL0u+bpIZ6W30KtKyKy7p/+vRdQ490E"
`endif