// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bPJsEF2KIHAWVyuvx3vawkkzPxRpg7nQ0Uf931ZXJByLKoTqu5TCK2SLbelA
3TRm0XYm97NG/f88qcgF6PFXDX625g7DZLSPI+qcYV2nJIW6jqyfpApO7Jze
oi/jRW2FoiwStKZu71coCbm34APo8H9mp5QabIklpRsJR5TxU4I7JH6M1EcT
lLhBU43VXtcG5gVS3rGdPqdwLVrcQQXDuMz+37sTAEiRNeIgr3O+sapRTmQO
5y6xSLEDmK2oTrkL9Ctg2oplEW8OyqMybUOlhn1aILHm4zX8hJHnLJYDKTmH
PmaKECCQ3Wx5Z9qM78oaEVTnJfL755LXD5/7Jf462g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SuG2I08WrMeS0+U2+5IEHAO/gVCQbWBxRtAC+MfchK65SiqNCsBau5awtF7M
gwcz3TTJlEQbNuaU7YHX2/SHAUcbp8JhB09B5ep3MjhisppD/2rBn1B8YE2F
Y29pKfhfDB4ID//qiFCv5Yx/UEvP6MSAF7CtjTS0F2J6PzYc6oJnvcCiN0oD
IkaogME47r4F93zHmGoizs8bz5ldAhKUDggsUkPbL4ZyKZVwebbeYDEaoKUR
jZnoEBZ86hXRikg6sswIzJN65PQeVOMozwQUMetKpnFrSX73hSOQR+qV2Hfr
BW+w+6afvKBAtRawAuolPUkXmb1jCN09ZUF0gBFG2w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YAiRkAvhwWeFDMJJVT6SMQjiwfYPqUYJoHmsY9TW1n07rz0bWe4N3U4aSeHZ
FWtybhmRPUKEzcAcVxxvAMTgu69dAViAS+RZ1ogs67v2WeLSMQ9iExQ7bhbV
LfRjLZuQ9Yx1kH4QvqGSqraFJJ5STVKYsqnHbkwvuBGHcnHl8/jLHxN01Rce
4hhX8/sjs3gp8KCH6xpUsjgcA4fr58Dxp6XExaERwuE+79ZwAwZMC2OY6x0g
1Tj0CXlWsBhOtoUDsWe5uOShskuPqwrUDgcCWi4y+5cJD3uzMNdwtWJlsXtz
OKLILU0h0d/OlyRA7vVIh0ZgRgtAjF9CjNspL2Jwow==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WaRa3NPkFXwrOaRLnhzAY49mv2dAG+CWGkVCsehcBea7Bbc9YX+cEGbeB0b7
ira5GnVX+BTV56Ui23bmKKEbgT9gvElaKRfQHrzoNlxkfH7lWgw/9eOfYJ5n
KuPNf2q12Oohlum4p5AWhOi0S7cIwJ7MmETHg3qnHFUZonHJ7EJLI9KEP2tB
/NiHBMOkkUSxBUnZuDCq15CfG1n7FychOl2M1DiMoN2vcs9XwBDSXchZX4Kb
vfgrR49KJKgM3WmjrJynvrY14/shLoWOZUflYDlJeM1hDd7c+VmPvhzG3eiN
CoPHOnlgoXYEfIFfbAbxHUCZ9cKtsq8xWbZgvx/pZA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UPlerm8r4EQVFsOFUgXuot5RSyg1wxNGxwawAKHGze3u10Sf9GerXVBUZ0iG
e3eI8k/coKRjENA+hHcH2l4WI1cWZ+mAaERslXXnOFFo0dEN2d5wSb7wscj6
M5PfGUc+4ruExsFIJGpcGJBcuJrpIUj3JIl20ztdr4woRFWuN0E=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
p1H3OWmTMCsOqGJPazBlRP3W2qs5K01bGTs31NkW0ThLOkPt49YDtfYyjh7Z
94Cfm3t8a2THJ9VMteCJ1WzWkhMY2NwjFR5QdsoeR71u6Fi3WO0KGU8CUn/A
6Tr3gVlsJrBKYvmYnUfOl0TwMVD06LbPvsWHM1leohiBpXKxtkgBermCjA+N
8wJnVGampGZrRL17cuWZk/EHgEOlcSoSPhZWjDmSglMvYNn1fWE/ou8FifBM
ruJQWJtnnOMulCPo48PfkPYm1UgpSNhqJZJ+7ahCDvrSygn/JHm7PRrLRP3a
9P4lzb7L/qyR9+iajnBFsbycg/68KWyi/Rofm5INOajt5KuzVwYtnwML5hxt
GbENCE64jHtvVZcc4gzWHkg5HhTe68sg5kaTbZ5xmHm+pm6Qy3fjd22ONf51
ze1SM9e4Hhy4TWlsEzeZzs/mPtlsfGZ4cQcZSzzPjU2SbOPwhaKwBF+ksQ8t
3O3MSFXLjucFJZ+Ev0C+wDRRhNZVOpKP


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qCqg7ftzLehCQ5KeNPu36DK55cq/wuohIz99BFofXtiYw+/rZqTIsJ3CkT23
lLcMO4uObb0hUznjQ1TY3pHvb0lNu9GqxUOllNhiQocjCnHWgtNN790XDCDN
VbLPOy2F6M912VCXm4exZA5Pw8VZKEwrV5ymasDBOQZDpMMokGM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cYdJAww5CvDCIlqRr3CrXyOI1TMcowGGZkeJkPIZR4qfAzOh5ihLtrkWO5gi
5cKtNi1mUGfq7BrrJ03ieQku/lIVjaGJEXLG593Fc1pqt+8Y9ySrtthqmsuU
9OolhV5I4tUXZpzS4e2knb+WPbyf/4YDVj4ePl5dCPDFdjwawG0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7376)
`pragma protect data_block
T3ewVCne6tQ2LnEK8t/ICp7nhc5Iug/M+NxuuMlfp1EH32t0pY7GaTyBXDBl
BsUDAy8WjTvFxat/X4zPldeZWDWEjVwohvgAmO3EBwWT5B/OQHoj4wzF4vRX
QIRqTqJz/KbQf1hsma4UGIgiifdiwYeHuUKPgniUIkOxxxltwV0dV0mOnUG2
EIapQdKUWcj8IOmEKVK+so4kKYIsRMPgINp7DBpWiDec3qEahBW9OyE0RknF
vvlZ1LclAGLvOohvK1miDD7ix9JjBHeBaGr/Xhm8+7fPOzQ0cPSCEUSgAzvY
HF72QSCDR+mxa+oLWzsIn1L/Ew1oVEenhJWmknGNfiUy8j2MUpBVqaH7sS/7
iAht2v0Uacz7qC0I4+yBu/1ToW6Alk/qXDdNLRCpQ4L0tcwJNGjerMymuGyI
oF9/W/4z/uVm5zplgApjJlDg3Rsw0rELoQLKI+W34kOECXpBgFzhLdOWYqPR
mM/WCJ4ZROkUkluQ4ZhP01ggQWY0lqsA8uXCcCnx5m3IAQlIn5u4V62tb+Ws
bHWe0yPV8gEdJrwfnpKlHsYe22WAIlRXVA42JGnkeXdFUWdCjgSkVYoyTiXy
ootQsf9V13OGcAOQ3WcjM9OPGgb265QLo56VGiEuKL0iXv2ifcKTdbmphIEM
logcSiH45ZrR8jKlYxw1FcBvcdbbuQZAvQRGvD2vSqSQGKbMFErBcffx+O9d
r16/QzmvK6ibLrspJhGT+Tdg80vWdtauwRTnNDeWym9GrdUoSTL8vkIDqIIR
AG0KEvLFfgQqIHwTvi27K/W20oteHWNskB3AFeK2BUd57AqS4hJJXKbxQVWD
GMT0igfOiI9MoM/1mPHkl8E7XmMJvWNP64mXKjL2IaY99w52hx7ph53T98IT
ZPQsWkpV03fHx8iirEtC+URd40AV0quqDJsbfnoPyBHD0wpr+OWclDzp5ZGC
5koCgonGoho6llVoc88gSWzYGOzCfhmxi12fcKzv2epgHPshM/Jjg/vp1wZh
XGYb6rnQZSo4lTvpp2QIXYs0erAeMDwAx5IYnQbXRZRClpztiUZTUmUrDHq3
/WaJ6B6nppn2oqkQRa1KPrEuFY7Cl7SpGTbd54JwWKK1ZR+xN4xQC3/0bCSr
2ZjH/c0p/vGNyiWJJYhbPTAe2VNeFwRcqGVepZvYwIHMQpx0fWcLO51Q6ExA
G0UvL9hHlbQm2N+LH2bOFtvmM1KzZeTGZezcBY7Zsfj20MggTaGffFdgkol5
PUxyathU7ivQpcEe3o0v3z0nx4ue+oTMv392txpKfu/rAAF2YQ9MdmcJPkMD
7sks8JOffvz72QckP6FQRBcgBIlqNrX9/VnPjA6DCT9VUIcq7wykhBErgNER
0CPjVwOD+0I8rjZ8dcjmJCX5HaCVOid/KC9q0pFQjVvZANdznZ6DDUHM13D7
wq9Ny30s7scBwp6hx6o4K4Ozw4nTpizK8li3RkXxgM948ronaOTEHyLvjO+A
DLwRsD7Mq7LiUbvVG0PnV/Ww/PdvG56WzQdhQRUhUg9lLV9VCwzE9nyIRBbp
VQdh3y0G/K28S+TOon8jBG0IgMk4H84mL+PH02FNX2IxjY8agSyK74Kg8VEI
csS15ShFSHvoLigG+lq5rXMY+4gxg6eFMSIhrutlqK9jiz+S4Y7n0Ccm0Gw0
zCXih4n/hL1TGDDxur3qBaCqKv6J1HgPV7IXNrTXpjFMk1PcbRtoKtOCtpzx
Mw6x5/mrLb5cssO4Avgugl8iKUnIl68L/QL8IsgfOdINCPKRBRXzf+CHdq96
FozBVIXNXSy3MgxVmWRuyNomPobCXTb9YcZecR+mCd4P2ChqDqew6pvR9Xsm
Iw+b4KP4mdQJ5lbRNAk0vlEmNhiZGifNkeaO+e9rwaCJirAzHW3xybB5nd7y
kU3KTF6mJ7JHFmAgUI+OIyNeSp7Tco0jC00iyEfbf327AoU/8CQxDwdvxNtT
9C+300ko3WvHftSBqNHpozY/23laxKAjI94FrmaF0Qgbrn760iKdPA/7Ig9F
3tiiCcf9M/JGCpuFPUhdN4f79T6y36fdS2vep2NbctksU64B3n8GSrSvOFt0
1NIQgmHGBxzYwGZwLSk9HIN8y64Socu5KmllOYulE6GUxdPF4trv3px6S2oF
uRgQXcLDWwyE/pe7jF0aoV25IP4escaWkNagHZBUs+Cw5DlG5Rs+n6KTc46b
fqRaYJwsGXFccQsonDvzGrbwoJNHztQuvoC3jpJWMZO1ChtyvKODBPAGdiBA
eUj9HdhemrsCOQaFDCumyI3X7kKOpdqFwp8QR/yZepDFVVX8b33ltt1v2GHh
mLdhkEbQVJsFcWPciAqnV1ln2FfEKZCcZdaJUv3ZP4jpFaDzcTcFui24DWJB
ZPnoIEa7lUvgPCj65T85P5hbyjXwB+9cV9wgyuC4Xs5nbHR5VKY6Jk6w9+CA
/VrqmFpwLZ81Yn2Mt3Q1i1igMM6XsamkcrPDbJbYBY5a4ktlDS3AafYvHpOP
xVRTImxdv0c1jcHSO8H9JD4+m1RLsPpwwZbLL1jk8Fl62542SturmH0gUKn6
7OiOL3LNFy4DTkgZWUDDC6fuwVtTJwDKwPmpirfYYC2QxjBxCRE5X8+p8AKj
JyFja+2BSQHWIqWUc8kOhfaEU//r+Foa917FFLzC25YGqFvv2WEK08dbxma1
sEMYxZJXk8sSGfKTrv6Y0ecoWFm24NNCSGTDJpNuSqwJ5mbfkepmt6iuxzs1
RawNLvy5yjUiMHwUxY5T2IGd0hhxj3fe4MZoXuIY5XomfPl8kZd2o4hY323p
p0GpbAws73sJxiByEx9tyfabkDh/1WiIOkWW0BqXruoDg6nfni3I6LUtGc3q
bBwwqIsjYK1UvEzClBPwjcdc43hYxXLqnlaZipFY9N5nWg78TXzR/V9sQAxx
x6pOIxIccgJWYhLbGr/ao1f96dOlTXnKEgJ9CDV8BiDhZMdsSXXOl6Ow9oOv
GAWIfPvxf/1570AWL59A1y9BqJREj3ACDKpue/xCwKuBAPbKwicTIQPr4mmx
DqR2xjaeXVOKti9eYsyVcnZYwgUIsFY4Zqeku8qyyeN/3ovTsJe9JrypxN9B
Einii4hVYJWp2pkw4JHiQRERPFTbAy0sUyIEcV+jgz73e2QVLMWqfjkYzPNZ
kfv9IBYiCn9xSTmqvLQQ1vDQDkp0OUdInSvRU7FYfzE/qS9+ksDAmg9y3dU9
fxoUxpC6SwRAYxXyKPrhyhLEky9AISwxan5qM8jKXIlX/wlxucB69OiYAR22
euOgRZCq9kiVwlLeRGu0LSji1i0JWVdeZQeTXQGRlmX4mK+nwtD8p2HaWJtR
xbiiE56R0SLEFbLwI/DWnOy9YKCgMCMWmb0InvxGHQxaStvtqh7sB0TYIgEU
10opKJQnZIWiTXZla8UN7IkZ+2cmE4qZOthAQTdkzf9bKjY9xf9mpkZ3zWzU
sRIgv0UhgV5Vx+Pd8ODdTU0sciMloZOQOT47SK0Jl0jK/FnoApglpJ8kyzP+
gFKJKvdqBujBzYDmy0Qpi3SiDg2rL3400iJzzqiX0/EfSvZSJPOIZ5jriVq/
GA4KfO089Vo37UGUrya2DBHHoSLCn+VMtcBX5vwlqU2yaxlPUuFCvUoryGmT
uxcfasNLlqVD7sg89n1Dfh98oo53n8QEnCkYKhOXZdnv+FfE02M5ltEzidEz
1UI9W4PXwd7Uc1UXde0Sd2K0KgaeLPSst9cohKvbuoW1hduJfTIlc3qx6od7
wl+r8G/uxH7njxmXHzS0QHU3waQ61DulE6Ie9IMdNWuWsshlpOvY4FZcvSg6
0q9rzePlJmrCYNV4VqR5EoZ2QcDZ1qAUrMdI/HN+p69kYVOJVB58+sAB0cop
tmpE4SZuMhR1A4Kbu9i3Hiumw5Kcs9h6qtac1kf/gW27aQTaeXseyUB48iUV
Sk25z5Wq4+MUnMQ16eQTRvOoKJJgEvHtMUves7AKOx3Jjz58QnYnp2BVBjpf
dUjNPuF9cCvyt633WRb0Cck6hbep+g3XXHN8I7ZmezBerXYrsnc+ZTOfTf20
+wVnI72LrD3kGJzOLoWleI2exLIR/tcbk8wzs4OkFCehxfpUYUlUyc0qlva+
khl90PkjHdfcYCfKdAOjCkvfDgjhXwvUrJVSKXMe5o2cYTALOU4MHD4j83BY
CVsqa/xgjzOGUgmWJjvSZfOBgO9AVRGzZ9yhkRlnrqd8TKlUC20d1vmKcb1V
qCiwUsHU7I+DX0E0AcvDq9ArnkryDtDda3PVytINywTxrGvmQGFhUHSV8NZO
3TFG5amV69P93L13YF79uzKQpWpys/UWs6oR/eKmw3vy6TwVTzVkJ/76I3MW
P9HYE6dwD15FtUCMVMCzibc2HRigTZuNFmkFog/7J/U6o8YJR3oLWQNMKYvU
Khwj9rBSeYA85qM+OjrBjO9T0dkJ86AAU/qZetAhvKrhYKyVfiveXIpGSLJf
M7dMSMKncWzB4u2/6suqpj1dxaSs7ssKsXPXRNAHLS91AzBDB6e+2003I3SR
Qm+l1ilvnG4bBlWU9y+1h7qWjKEMSRKqNFD9pDwCozXiVwQkzoh8dPA4SVcb
oXyIkrkagnZ3YjTr1cLoLLtM5foYJxTh24N5TGy1ENnFlRacqLonv6zypkNn
Y61aryrOnUXEQtHrVAdrrxuX6rFpcl7U1MTUK4n9KTxjhng0gmqkzwBeDfgz
XuiTr5HS7RVLXGwOTsXNu4y56Bw6cAnHrsZ8Mm3laTBaLVLYzO99CqIU7hY0
St4GkrglVdw6hGwDbCwb9lIZomt3gkvSq8+YhZe1ZgvBu0oFuOaOjYTq9N69
d0l7d5HoygzhBizUOp6jHeUSrMMJeg1NIytnQQJFhDP0V4GYdtjaxicy4L4Z
mzqiI7bMDZCsDB8Tvk2AGjUWMZTXKlaKVGU+4xllbSNj+ZlRYp58IS1uqtIw
wyGlyNrZq+5Mk9h0jIDKd9eNX+LFBklWsfsUIHlY5iQU5Gn9unj3zj/wvPRc
NIUmf7W2y2skViP9WqZL4qeYRB+EchcBY725+jdJsni+/UjARBA6QjoQems7
ugz4gqJyLXalqA0HkigHbcH5/R02LIpAxKHj6fRaj31X2LEe4lR5gVXQPcuF
ihfGsiWY8STgwHsC88pdLAtCSM0HjutzLKbyaCNzjm2HUU6MeoVXx5hpv2dc
k/7QYW7SvHvaRtZOggrXBq99EnX8wZhwVUpfkATZssfq8I4xHx5006ZqOr49
7q5wMYyJpjttmCrOPg24X45hkwnmHUX8lAJyLdd59PjDVhqeHvKUr+Ze6pH1
+19b6AEHYe+K+bdeoRAyhDv9vXG8idJ5v6uCzA70wEFidLAIk8T/nazv8f9o
zbsbEKeLo+NTAd4I4uSHaTbTL8mjVrBv2QBRMjJ3iGaJE6hjwOledvGxxiQ5
nHdmVMzExxewELf+EgOlF//Wi93c7CyFM+76mjXktJrxHQFzPxTkOhux/L0N
0EqNtVHAoBDDxizD71qNeRKL91KRkWvX2skWDGymj3NhRxenc//b/RxdL/9N
Fg63AHj89tOfgpvoUc/e8C/FGdXNDLE72xLQ9GfKd6AeINovDBIIG8uy8x9z
VqgxBLrkPZMl1+mQZOV2xPBXFh05Bbqk3hop/zmqGYA3i8i1UJnKn1cIwTkK
6p5Ilyvw4eQjnxR5wm/N7Qj2GvOVQonJCtDfHNZBSWA63pxaGfoJ+KTSs0dS
w0vZ3fnJkK1XO0ICKIc4K/rTH0dCF5Wo21Jpq2gCBhyP7Z1YHoTRgrBXUScK
DQoFoy6gXFOpDo3xTBL1PQsZau3QXighSTvhgf21q8j8xtIuGG67dsoJFyM5
sKjFBt8FIdrdj54hJk4gMPmVncv+8FzGGBt7hgouy90bHGPvHvBIdJYLkXkl
J/iA9wWRBFKNwGJbBI2lFW3CXUm9rvvVZ75Y5czHV6Qea4NtnCxV5kDrG0ti
SMvTcLH6aW9u6BYooETKXmyfdXfZfwAzRfui6Z8ztznHqwN8AFAW5fTIxuGj
JI29vBLpFSgHrmvpKx32pl8G+ZH+8DmH+6ZLphq/SxTTcDKwfZsstMRwtVkw
aiQk58eTqA6nkLP1k1Pdm0IXB0KkQKIFILnfBxf60mJfR/pNIXmEPgdE/GH9
YB5AQkqQbfWp2cfRsEaCo/LJxKIfu+k+43bYIj9emHYzhInVTvncgxTIgXBp
MgqRLvUyU2VVYjWQweUHCxxjkFcwrtC5MPScunUNE34uQpTzBeWiPcM2giOC
rmikLvFwzw3KoVJEoIr50khI3h3eQuL6z5oNlMSLq3jYphhZ9dUlbTL6mias
N9aQDyelqnY49/Tg/n6gmt9IxRd3xPeCV3IPFnuwWPSlRBIEt13vLVyNUpMx
ZhO177aXkmLqlOpIdisQOrWa2AN25emE+aOvtbmF9LGi/5EQSsDEq6tt4DaY
YXhizSc8vlOwbOUypY+XekmXW/c7w8jaMgdiyWE1xeImLd5rVW/tJXr9LgEq
N9iZwHRheyrzfra2hEBI/q7Z13560z4Zz/EeAAnP0vxLorSVhzEaw+MLXxv1
6Yht1kLKwzJpVOgYrTZtQ7z0OynUwZ6aXi0t851LJ3+zKJxdS/rt+9D0o7hu
/r6p7P/swTJiWvYo4GNZcswlAWYCok1Vs/qf7mBDPcrIVEj7IwxKxG4Ivii1
uS29Fxm+qEqF+0l+Z3h1HHSpYNZUCPi1dO/3yzLnAgt6IS57UTda73gyVyj7
KDotDHSScnVIUv5ZOXwaaO9940cxGtqKY7XrFHUTUDnaQxUxwmYGORyncyIW
fdr/zterboEEEZgJfRfoLOETiBpInjxhHB9rElTxKQ51Il4U4WP+y+DTZZSL
UFxIjpcj0F2RXKGW49mlhY+2lPQtdmgM4T6LCk0BN7FrkCWkUpL9tZ1+JyU/
4k5Ms1x1+HMc4BDp9uSIQR7soOnRKPj8nKeWWoyrM1yuZbIjYs6tfTc7OjYK
qCxtAf0dn7REDAO/I29YP/+BsWucDO90s6go8kl3NTSTI6vAn1KJsEO/QUez
2RhMHtixZVOVsrFGB2MbxnIhAUMynpjVf644muKV0UQXij0IXtK37YyJErXO
+E9VPTp3/KtpG8+Pkai35wKgB1dleK2CwJvsZAg49Cwx7X9rMg4C0cHi+qGP
b++C8mvi4Elpaq842HMKUVXvJ5L4Y3TBKaaIgqL4XqhksfdbkRc9XxPY7F9u
Pc3otVi5A0Zw0IPCGMzFgfrGJwM8GIvTvoCLPynXT02o6B62IOrKA3QQNCKg
kFPce7qA14Vafioa1aIeua++ZAFC95A98P+VInA0lqeHPG45Y3/GOdmOZAaS
oImFOgjDHwHvkbpxwByzI2RlCFG39Tlg+3ebdFxoi8sIk3qLLAOCE6ywUpRR
/WYzgecV+rBR8l1PAgYC0Eci1LHonkWbKF7AF173zTyckbWnhgzZrcQjlqQs
A/RYKDpZNIJfHGJ1fNuC9J9wUP85HIVNzHuTd00+gdqvz4AK/N46yxby2bsJ
u1LWq2r0HWW7aH9mWC31AMHPMeckq/CfJ+04D/DIv1Z5S4YcaW5BjlOFMOKa
icxz1nKmX251m2Y/1KPOeW3YJNIBWNzGU9D5Sv7z1XH13EbFAAxbesLhtKLE
mu9ZQe7rEeplCdAqaJ9CI4NaZ+1fiDK7XTO30NEuPlMaoZKkn5cINS4oDrAN
XWLjxTMjMEP2pzfgQ9rhjw6ihGWT6+AS4tw/lmpqR6cSp1tgg1cTUbvZ2Hqq
1hprPiP2dELTy6QkYJhUdv3uVP2KhPYW4uUT/kb3jQfrYr8EH5ydx/9Zbtmx
LFdZv7XWfF9cuMp9VxEXmpmYFthG0vqz9NPZTQmteI3yTILdM8kDh60H4pQu
IbSxu8rLHD1DAM15bY1zj3LJtkX3LqLjRBXqgRVY3LkOLADqO8AKNfuhk1C5
url5MxND6tWbDgN9byR+AxBAO3MhAzd5LZFAVaWV5oD0Sfke0sGhJ9pMNryH
WN/4LQRJ3u9+iKTFlqlZ72ARNKn/RCp0wkqRm+tJHM+Zv81YTzcvjNVxf+Ff
q6EPVsiGNwvJOyhd9P0sd7ez7HadMqxeTeqzJElqp1vMDWPG1dfkyLQerN22
xmOGGe8vmlaNrr/FGhYxEPeHjqrJnLpMczwt0nyafJyorMHLK8tfvPwv4Btx
VdID62dq0Y3jFoj6pHbEiEefqLichsa2ZiHj1NKBhaZbWy9CbIYycTHyNkyw
gdpMbINmdi1VnRLCDydigJde7HQuZoJO8dshwQOzocfLh5NCY9DyxrglFdJG
TuY7/e2ZSIoolzZXQ9XEnTLBc/iaB+U/9Bz0wYWss/9uoHi/VN2Kdn92ihao
ZINNSRWyJjNY5Pcp3KvB4fHMDW6Ku7J0sQ4nwphQVFrlbWQlJ0b0XjKPNzHD
BqcNn/juibb5twfhVQ9BuBbOlaroPlN3DBVaDML5UDSitcfNSVGkUriuhN1A
wHu4j9A1nNMEEumbMahqcAnL9towEhVDrYEiZHb55jSMyYTu1vl8TZrI+j9Z
kDmKUCUUXCNbSLUoCyphhO58D0CBEbeHXZHjgjlpQxWy3DQf8fBthpK7OOsv
uqdRcMmW6gPbRDtxVjqfYP4iHLp2gTgnU4JyX/hOQyfxvcfeCRYS7A+TzlIU
TriZnkvOTVSY0l7bRFgMRgTGfHDl/sabygjxHjqPCYHN6/OyFdcEilYBR53A
Qk2rynvQdPFmvVV1ushm9JBnq8RagvadvbJwUae0Ejydw/ia9jxzBmzCY56P
5WumVKKz0ZInfIkwqotp9VG5SGbazZkd+jQYk9RePtkV8n5R+7A1+bQXt1Xf
XRjhtyswL2Ow8z5Sp4OHctK7qurSajtcS2nSvhDhHUsFFJuAKdPgjBIoyiMd
fWMZIIfwtJFKlvGF3sbcDf/Md60jh/KxBGuhztDc/bZa6cjOsXdlCK94aeFT
/Ydy+111lJrR6VTTlE+kkwEMUCPZyCStcquqpZJeZOfA3y3fv8wbXUeUFj7z
MdRFhqMPTzkSdpJ31Pb9qlQ0ufdyfjL392H0gJkhUFbK+h52kV2kRk9xxhOc
DAZMrJXpXQRT0NOxvFGar+1hXzr1uw5fVN9y/38id+nh7zcly9tYZ11GsqQ9
jaF1XL6cgpB/zVF6j15P4TDaX7SyEqmBO5iCuRDgp5RmOXXduE2cx86jrIAw
s3N1e8ZXheBFMu1p8ngeaROgZx5apcRnXaYEa3Gwl+/qTXfy4fBfkU3bDFbm
obj7ospYlgQsxb1piWzRq16RyO6aBzRO1faIv9c3FzZSnU2YtYPgViaoRazZ
rRLbOqoe9TDOJttjcZkhW+isRuM5zxyFVXG0r/7GRILNBwS3nXGnLOlTG+bH
YoYxyHfVQrWHoYlblwi4i1BPtR7cyjILm9OzP4k1ThTkTuS8QZleviCBG0cY
M2ahOhlHjLj73Gu/rYt+tdYAkP8NoK/xWJNeUCtSJAo3KoA6F1KeCVQsnpCk
YovWI4N9sAXuGpsR9nadqlWtxAapV3U0U3h3BecYPIP949PxE5Zh/CI46kpH
XF8R/qCO221aewc6cI1PMmLXR4vCmtNNDOg2jKxGzHL8owJcR1uKcerbtEiY
6lHdCaFp0z4b3tLdY1BSlK8Im2xm/f0JJ8hqZkl+CD80wmMIkuxNp+ferIMH
X74aksiE+6CiyRBg6WkCDGwcZrr18VacXD4saqBvKCSgG3+J1w/v/KBMLAXI
GBwmwch9iWNs914IfAYScDmcBwznQxZ+GunR9dmNfbzWLwgje6Z3FgE=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzdY/VvSHi0/EobwaSwUc19Xt0ph696gLRwzncpfjM4awO+PGkCMGxcc7NYE7KURq+eKPO2k8Bb4P0YpEokMAXPCg3PEKjy7c0KPXrpjCYLFHLosG6g+CNc9if0oCeabJT9n5A5Z3Jd9F+K7CKO7UYfAJ1/Em/WfJ9rZIU07qcDZUZ+GTAJT3lmJ2OvzAZ5FJ7ThbfZ7IR3KduSXdF8FhdpfGV+3LTkmH2baX+r/QSw7DuCyo2r+jGoGUYRRnnROfpVu/dZ7TGIdnM9pld4yE8plVj6bNyWab2moB96CzmzDLwHEw/UodG3pjsJa1k2RjxiDiibY6PLRKkuJyrsujg/x6My2BYF/M+lXuLIsZTBB1+iyKH9Om+8N00mfAZC7I2KtWMMiNjpL8W3UJEuAvvZPYroO6Q8lYFD0Bm9exn9B/gUt1SV1ioiBa/PGrO/mfNTynL0fPd73wwJCPYwRIy73EnoaQFTJG0pmZ6fknNB/hcZ9brDp4I2MW1LcD0mCNuTK6lg+eXrAIG2MrdMkga+SqN80MDqK+oIqjWaBNW8BF72Io53WKsdSHplNFP27uoiQxo4z1hUfiX+STiRVZ4yYx+FQt480Ccagbf/vtsqk4tRtS2FqUpsPT6PzT1MrdjyC45IR8r8Yk7vfSV6hazbzrmd2h7Gk+T5OD6+33tWx2PTv8VY2wn2sOmyVeoSHTJjRgu9vGMt+q6PJWsikNhSk5Zt92mRtNwcfJ/ieyiKuYlR6sr0Hb1ti5e1pkATkPyH1TVNOhJyulNQGbZ5rwsZ3"
`endif