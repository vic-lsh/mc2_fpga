// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dE6+oaVZPhvJmEBe9OLObh0e5DW7yOHdnxJtyEjnwtrOjwcNUZF+OHTGL1so
CY6dp9FuG/iyB3/zuTxfYD5Pp4AyQP/G33os9XeqaBPKiXYNDGiXV1pO2Stg
wXgYHJOEsIV3/oJjRjL7Duk9hvz3PR5AYTRL+N8BrO79VYLXvkynF8GxPF4r
Jpi6hiPTt89F4NgYUOUC3Kr/C6EEctcESMA3/yO3BqsAeZfRZtVVizDadLSu
gNb7hwk8uTSdoNgSBnHhDifKfmTWT5RNtm3nBszfWuMq8AYM1gZLiAUJdrAp
rHse702wqSnQ9oeHnUjZtZEq2HHBVHPn/Uxi+nGp1Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KVFzGy7ug4Ke+Q07ecP1KloK5sONd1fj3qB8Ea3JsOfFaDfWwAQwqDiqJrsv
OmbdOIoJnvKa1CopPzjDbl4uvam9KeqBIP3MJIUS3yDh9YM0uPeZILTUMEUZ
PbnIuQ4YPdGpek2xmX4E/fNkSsljez9gv2v/6iVs8wOMghy8HPxBIjdHNztm
OLjKOrWxka14Jld2nxde6u+6G1MGLEVWt4fcGV42KTzWM+Aq+UzJaK4+f4Fo
KfCZQXceB2kaXeIVwI9PWGP/mHDpiQmp8XCQXb3EQni5tNa4s3qK37LWJuKR
ACQKsQRs6YR+JJxOheH92FFsecowUtRK4Xpdk7Ws3g==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
L+SUQKbVgaoMLAIr8TBXRQvYfp1lAoa+98Hji5YGlodxJZa7QgD7ODt9bohM
HD52dlJ/w4eySdEpSbMcz+mQXiYLboPZYuneaqoZ/xaTCSX7nq+wXckAAA2b
7XXWhtYYYusyuKQ6EFy3I8UX40rJb9/TWG2SdZr+0N8ltJDySHx6ioPRNGD2
UXdXCHij5O2juRytyQRlh4OO+qj8BAlz6bwAuv9KMqYRkKAjdNClfHYawcV1
Z/crbjG6YaT3iVI3x6IFL2G1HcK5uQWhLAV/Ii+c+xNRs7AiQKn8pq7ll6nY
RloUQy0Bm3wtsL1VVGnNYgRDu/p9dr92D1BniNwOTQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FEwEQOxlEhb7Ty8DKwHEiIQI9x9RqQ77frauepschy+FmTSJTz4e9lUFFBIw
oi4Wogl8dWekDKQzprKG/BgLdEGHEnQFn3KXTmbv86xMcFJiD8Mfi2f+WQ4N
7EiUlHZ/e8VCPxAGkgwfZiArrSL4DhlLgLyy9yCuRpPufmnbVfPCyCoOgAZ6
fUZ7sKI7xMrSF1kvY7f7Ys4L0Q67qsZY7/n2xn6FrPFC+caFwad1uM/dEZuJ
yZ8Bdtot9fGRtDp5+ViXnMZSgmaVALcN1rqNCtqFhkVR/+p2LLcUm8NDjx+Y
pGSllVtOz8DCk5rW5MZnM6WxMzn/bYhpVQekY9fKEQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gQdROarx/LIWMRBAOcmsausX6yfbvN2ojd/TQV0lhanxPoNzCBzoSNvC/tzS
LAn90h39f16Eg/Yah7urNZ1RPQog1M5F/+KV9d8WVMFikrZH6/kaFvdwJtvS
fR0K38EscSKhB8CH3kpTM4fUoKMCr47Tr+TJQ83JO1iWdHLL4wc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mFLGcwOKI1NTIN7aQbkWBiWWw/fphSi9of/AFulCEuq5LNRp2OMeSRol8/mc
ucKFR62ZruXYGmH/3BOI1D6pMKdf31Val5lmtkpJ2ZUYI0V+duFjs0BY1fVO
rExjU2IlU/FJJ6ifm0ZuX1fOZyLikMTy2zfU8HaRD6K//teI7ur+1OQPt+T3
YLhCx08ycP4yKlAkdy5cJbI38t+3urGFrUlsCJT2CCIvUGoWgz7f1xBA6Ov+
+VjZ21OwwKK1z5LEGpVJaiKnvJ1qj2F6pHrjo6bM9Pesu+63u4T9uS4janrs
DYekRFpeqAySLLX1jFl0E9ckmXSfZRSJqJP6qEInlfbnOv6T7gW1hjPYNUXb
SD3BR328Cpq942Jc2xn1iHi4lJkTLzRg7LhNcxLALIirdaAFtNDCdugtHM0p
BuGxE8DZuTKPHYadLjL2kBlshPUAJZ5v1f4XsJsvfT7dbisNP9uOIHRLRGhE
2BCJ+SwX/lr5/w3SoyhVZF773A67kjDR


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DekKaxzWgNyQ/UnlCgQfWBmd1QHzHGPA3g8Z7CXGpBKL4Jcmq9dr6CSsscdj
USAfDV3sMiM4wGqGd84wE78pMjOZp1jfDHTBqAi8S7sL1Jn6qMFf8xts8XFK
9VZUrIt/+uRHQ8qSWd3TM3KB9CtAkSTcT/uGzLM6HthhJCEe6Wo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LcwZ8789F6v3aZjE2lswZz6kZcha2E4Rt2c9yaB/ohao5d6OBIsTXxW74eKC
vdZmPqSK8fzAc3lrPM3TSdsfsKpLAB9RGNNJ/aMA0u7i+zbIr+PbfsiKtJVQ
Lxt6KFi0hRwIUUuEJ+MKsqU7QYizy1kGEmFaE3haunGCSkJXrBo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8496)
`pragma protect data_block
N1nCRTkpj120xgQ5rMDw5Jc35m//rhcIVMuWCS3BdUTnFBjZJGOLz83zG01o
WJxAbRqBm3e6zogeO1d4zlWSy2A2u4zqjL2c2FM/3+eXMFbeBNedIXlyR/US
BMTf0a8EWLUfVHRbGCoBDRqXp9u1Fg0mc/trW0jrPUvG7VIDQCSG4Pc97CbA
6w6FjbPDMRsjGAS5Ib1eTBHHzG4wzTNlwaTEDEcJx1gDEwfH5yBqKN8oqltj
Qr33KwG823McY96rrl1rv3LdYsGoGjtYiGCCJPTr1icrLUo9u2kNosv1u9Ve
7YwZWOHpV5SXK/L/qAGksaFZTKo+a+DgivOVCk3Px5mwOgkQfIjX2HkL72vO
DBqXW0os3LHHNHLNolj51ZlFmHdMum5Ayiroe6DhvyM3TjZYzbZVMzQ/PniF
5KwHnEG0jShL7oXnqlFm2DiUrZGkhZ5TKEIAh3tasGG8ouCfL4AKo36kKxui
fg1I71zjLSkyMe7A5zRXjigxtorwuiQj8nyNEB5Au39u1FB+i/JS+Wghssbg
aVJM1tQV40PRMUUKPhgUrtOvZncrf9lo9t7a67kxN8Wtn6gvSQdh/uhxzDbh
opzCHqVRtQxsU2H7QgEVLxpQKlMtHHpUkJsqBh98FPTAeePK9E35ts6yTSPf
iTUWQZfLsXFj6HpXDXt2uYkYq/hQaXiOfqNdK7S1xmTPVGNq6fBFOsmL6SfW
rsXYeEs/8U6LBPe/KCv5A8yMB3al94sVOmykAJPTMzSMYTyzpPoMsqccZo88
KBM9yaTk/QPvFWcWoFJF1bG2XhyFEmVvEnPTyE3uN5lg3hNlHKqIORF6Ttto
I9+P0C6fKCPPCzXP9ZMBTgLtwmtpwi8q3i/txRICv2RMHJwErjjudT3RKbRI
tlmrNHszpifXmqPF1kPSsMNL6Nn0GFsOIxp9caaPf8bhGvqR/CSMogyrOqvU
O6Bpsyp7HeV8/3XwXZKQ/fO98QnBMm2rw/Ppk1tFj6Xm/Z/9r085cL71f713
iZDXIeuu2IXXceiJE+BFiu6PVmpn0hBKslAFz8ZihCxfljR8ke0g12v40Wkf
Hp/HyMieU88u/boOSAP1zyByKbFhnDdFfXmoAv+75TWc1h2z2/BTkC0djCLD
XffC/dCuUKQjhuA0tdRw61O6dWD6E5qHVlMK+orF39A7ssNaDPPjkjmXVJMy
ouBeRWKvnqUUeihKf7wqr3hOkzZ3xOe4l5XwN5+n78JE7XtenMKfYkwmKd6Z
jsO4IceSTasLq7EucXopOl7D3vIJ/dhpONjv3An/j+xdMn9FWyoJ+8x8UY/A
q8vFzufGl7L64XpHhBP6E0kAoW79jWBRppGTdixwA5Ai1S252fbxRGPQIO68
hWKuy4vP3enzLTgO2uIg4OPdkGy1vi3eVbEXgC8qLFIQBFgq4BiepuARcD7z
PZ3CYeFoReN1zjqAhb+gTonejPTqwluCKtEJit7MYoxURztJYneFLbF060OE
NMcDflA2KNTc7awtwGHmWWCRUMN28ora/RsnjmtOz8bfFwaFCpI1wEbMpmWc
dSaByIUaI1dOOMS7q7bhG5XMa5MUwuGhEbugAHw4o6uKUrzLVOYJthR7G/MQ
37tfWl7HaUOee0v2FxFe2rhwfr+VSw9o2Q+utGhvtsyJFsIiWulYf/44SjD0
b6vE6B7qgHhxQONh/R0Vem47520BN4swjGIf2jd6WxBsWrTI6bmZxZGKJXal
BHDuV5tWMYuAe6zCs6WHaLKNND5rPzRxxjF16bvAWf4u+vOqCnfj08yIXc7N
EPK+FEH23eDmsipiD6+j1eZ6Fiufn1t/gvILL9cukXXBcS0anB/bI9Gm2TyN
TkjpEkcmBaFChhV8DLQpjPGFRNpiydUDAfCVZC26AOrHwGsHzQlkzQYwBRuD
xb74twaR6RMsXkhSFq7/R5gAhNZbvOW0+MXN/MdRDjDD/DjFFtwYOvwtKhTf
HpnP2AlnY0A6R3klAc4T0UlmhXmbl4IZxsWSWtq3I0dDdfL2/JdH9DkzAKPV
1QsaqhFkCAhZoacic8EDusDNDEiSBdhPbLCkDFe53+Gcgm+QzrZlvXIexDsA
C4sT3d4ejVtmwvGSwJUnHakSEa9byJ1vtkpyL0ed8d9tK4LAFtbgCii4u7Wt
rIWmaJjjLaEcigDO/NjbBNmFsdvPDmQsrdafC3Z3XWHi6qTWvMKvcvszXIqw
aAeetkO2f2CIG4Gg40raqvWQL993RvbOzru+ZZMcKcSl4bp8mb/sUNqu8cER
Z8pYtpk4/TGY5gZ3yBIZfX+58dLMEmlKVK+BL/AU2Av2xHEQ//vQe8Ff5ms7
ETbtjx6plnDIaqMqt6p9GaCRUcW51D2Byd/Sknky7jWAbhUzpbWtRhKxsrHr
Vyhn4LkaldZpUQczGBSoN8gVK61eQSDVxlnOvfDeOBoLvby/ad97joeYDLrv
kIeLsM2DR4yTmtY2DJFt4pSFhDD9ZN8RrSFW0MHk09GpR3eKU5ZcbR55QLZG
G4cUtpNK7O2ZkBpoxrFO6XHW+Am0ws8zfJ2fB7ysJNco2e+I0IKj3xbbfebr
zMO2mZwPr6bikGNiGhtpDT0OT0rll83jhsmrhdjRoqfgVN6RnMv35ZQXc9Ub
kg2mtQmiRLVpBwI9CE4h0xlT73aacfEEoU7Q0E1YytOU3tHm3jeIdHy9yw43
LoYhMw+ZNOvUKRGRUInWm4QID93+ZMCzfl2ljjjGRUM+xf6F0Ep1bvFH1jUs
26gi7rxdjaxsBLkNYrf5VoAxIArbLPc74XZf3nFY/faLW5bEaF6Do+WHhQZe
covQqWN9FFfDZFqJOT1tUyywNJvPRh3v+//S9NPyJKs+6AcbFfgsDU314uu8
+hrMrX5mq2Eht/kNjTX7uQibaNmG9KkatT29HZt3u21fnh0cFfaP7eh+UtNp
3KSZ5f9C14Ra7Nev51sYcI946NCxfyZMXnRpMa/mBiN/JSK9AWRG+Tr7n1mM
zS6KaQqbeKoFYrJyGfUfY0uN06rEeLXCo6n4JXzPv3Ho7uzgRfAOMtNrxSTm
OTgpTKkovEDn+Fv7Bv+DtLh3pNsoz0XsuDBehEznbYEy28E/wfTk3runzvsm
zbl19M0uirM3PYdvxbkL+6T4YeApBwoRsiYcqg6UEnTQ75XFvHTr452Gsa+C
UENcutt0Kz8V0S0FkpiEaiZIXXdAhe1UCvWd4PhoMLWHMylvqtw7SSfjk04t
NiNV+7PsiCLh8M5zBeLtImrby06+qLfXoMr9bLQCgzeqEmt4X9hU/7OHcVP8
0fAzUMVz1mdjJTOjEIbBmTb05U3WrTRV85+SPk6QBC1Wtidr8GgAVZR+6KKl
erYO7yG56ulF/q8hvPEiQMimbdcH4U2hU44RqwW3oL85LM8RgrltQzGL3Pyb
gts/QNrp3qyKaqCRrltI3uXA6flO6WjNLAQev6EiSKzNtiPx13b84yxWDrs2
fpaJDqpjTZejTXIGfu+/nmvJI80cWMwumxKDYlVaZys2ODV5prjEa6QQCri9
ZMtaKNA9N/KXg4+UuYJQ0o85eqJSB/B3dqJsJfa/PptKd/VP5UkMjuBdgDv4
ntyGWDEhZJ4/RvGLLZQ3g1p8OE9FAHz+nu8ijJf8iwyDnHhqEeS2R75Xmh8y
bO+U6xixkWlSfUqKV6Rrc+Ec+j1PXXL1jv7WAItMmArIe+hgOS9SODU5ujry
OcaAIma/oUxSZcLWXCYgGsc/9F4eB0geLwFG41ZCIa5qq6QLbNYcTiti5Lti
IjGGTUTAK2PNroyeKw2MAI23P//gM7pHaXVDs4XqDCbdFtZvanTlGyXmQe+0
St+4rbixuAESmHigCctzYUSSm1KXTYQ8Vhqeu89ktvoM88myPD4MsHQg8a7V
9gNBvUPtwhEB9e7DoVqWj3wci89BzJpa+6yp91fhBKifUWpAE3Qt8GuDfaoa
DxpofKfVPzCve6kbk382GwO7Q3jOKQCU+oxjiX+rqLE5Gg0YrQLuIjGn2/aB
60k1PaMK6M4moyqUf/aC/Hg6HjepgLYL0HHv4pAGwqPXZ2jGBcm65mDr4d09
B8EJSDKsTXLWKGIhKX80lnhUT4syE2rrPGuWijZug0YGocd03kstqNYfFgjM
6yCjsXVvEz5Co9SkOk2zC3ghzDinzEBGcrC6sJVYSDrEFoILTekkuH1pMZ5q
SmJXijMOGSr1sG9H0h1aoKp3AVOpUhSkWlKougSth7u7yqHTcHLR1c8jTzqm
mBgjmcQymcbYXTLDaHnH1u1rCqq5va8AA+BWBkDnc9RXvwRp7p2n8EoDoLW4
KQYl14xvEAe/ZizMulHocYdoj1j7721PHVKJ4MmckppEe3xFsN57JdWHwmy7
EymSi+Uu5YRhNt5IN0r8HByrcJBpnk7GyLmyH2AO+Ig7HAPyq8QpB6xsyduL
tQ+W5ImWEIHJyeHGbWmpBItdKqP3S1e4Lkib/sOFgI0SwhSSOPTa+dFpIc/w
VVyBAauQXsempejvG5bL/EsXd8My3NWWD+DJaf7B+Vf/LmNNgpqJrJejHiJr
VUFh3+xnQdj88u+MqZ30WZbAhSZ8yRLuF7Fv8wL+nxhPXm4XKvUzGtdMFAN1
jkutymBS0VEmGYQZckgegiOfJ9ZMAzDUgwt+ybbUqlh5UGD5ZIKt86Ib+fdJ
b3Ck14BNTB7N6EiZqLIeIARinbPzJoYozyKg4lbLab0Su6v5VsuBs+oPv8Yo
VsgVYHwOmWZbLXpQGSmH8wYR+iIl99vOux/0cTZqVkTl+vt3jgO6JPyngixE
TQwrz3gnVY1Co6zqTszw3//i9UYgRAFfIpd1sX90mJ3nUNOcvKBc/j1QV8i/
d0BKl1S5o1zUbWqMdmrG0bs0yp9afuQmKQn2nyskZcSgjzMZUvFO01jlEmK2
kvr7uO9JDzI/Tyqvbun+zEG6nPOgpA1Guc4yUvnjjiMKQXHMnBW8q6w47lr1
bXr4XWzfyYl61fHVIMs+1Kfizrbea1eMziNPG2oKegUvcUfQMe/szJ+SWd8t
yCl5PFcWZWAb97PWAN6dRJkoyeP+2gh9fyui5twjhJBbjP8FLgKP0KmLrSPc
qMGAkb7qsxRSXq2iNFWkjZ3c41JbdeBv10rM+BHUx1oFC3NzRtvLkYZbgeGD
+w4MCXXAWUVzutm7QfkeeCusZIM4gadCapRAJvMZW69TthZcnVjw5vXS/Q6G
gDgZQF6nsw2geYj6Z7i1fevJgn5jmGgkvY+G9TKl3Z9KGBxyrMK+j6INYyy1
JKc53d4C8PgLyPju1Z3SDs+rNVVxEkXviq4KxSVTZt6ZtM/qUyV+b+Mfuon5
dk+WbfFjd6DcbNHeBXmudukTnWlWBwgeSeKxV/OqxmGUC7u/F1dp/naDlTeX
335X92STwWNHT7MUQw1087i07vJ1HmqxufdPn9zdlvpVqenK+qgIuXWh6MFM
jK/GWpbTdfx5YeMqsbDPGVJRgf+2ch/lOQS9wprIaElyw9/4/DiBMZeretz2
Jv+irC5+devOgoaNFgw2irWWnNM9n0PS0OhkG7cmd7X3yHSqIBTV0nm0qA02
grUSj/y/FES+wFIUrxRQiZsrsPRvifHkT4oy1ruHF5aeEzLAC6YvZhPo3a0i
clB98cdvPMdAe19xQ6nXZLp/Qw/CbDkJwvLAaDuMKJj2D3RHLMoTEWYbH0Gx
Hw/Txbt5HbkL5UafNDrw93ImqtG1WBib1JrdeetDWxsx36bNqQL8jWRTBeKZ
P8vdzMCcsdUz16jwVfA5jlwZIIG1kfdByTj0PeIF7ItIvlxBbAWzgW9FY9PL
3wk1XjL5xpKUK02EzlajrzpbSuBGj/SqdtaRBTeDNrbTL++GjthkLFP7FYO2
/QzvxeaAeO8EKmwcuK3Ym0RqRSShppJ/c2xHuRYjjkPv6h6W0OsyNSex39GZ
sCD7Io2mNo+LRl+niYuPqU+SDN5GpmPZIvKGLCedG9y29eD+73oMmBKUqW/u
psPd/f2dTU5s83Nt5YXVFAsqJ4dymuO9nUIqB/jvblB7rula7nM/x8x7fe7Y
4HSYC/sPDg/4WUtxfhV/KirmrXYGrEQEPPlECeIuNQ1qSy6WhfVc2Y0OSZbI
j/By98JAaF9/76SIkK0W0ViRo0uNRVGMAX9GWcGQPoTqLMB+HWTXlGLxSzhr
UhGeeu+nP+O2fmP7nXs2+8FD7VJuG+mO8vYkHhFGjmE0FyIn78JIGlxcx1pZ
WuhI9nuoDuwn75mcez8cjBYJ5Tb33lBBF+UDsdRTjiU9ZQQXABhulDqgvgnl
tml/zbk2CnFm1yseqPTweh4CpoieT8IZAxCbmNh824MU8/IrCsIxE3QvLp/F
W/wSYy3bFiUf2jYU1WQAtRUcWUJbYJnEUtTfkjA5s4W/wnJLgMWFsvrxekVx
4nQFzMNK9yXI2LwaAzxbkv41j+O59zivOiuiKBjVp6hKPyZqu5dGfIZs2ZM/
Zr182x6+HfnHtrJrEuGGFp+G5PGmgaCjpi7y+IFC/teqTQ4zkxRcA3mRXhC7
ixv1PYuRAWbDzDBXbxVDvQXE+fpAbkX5Q9PHlxKJieeBmR7qP4CK0qEtZSJJ
RG7ABYjCrOVRm57mnUePmjyGZ2as3JFHNu1zBPb8MZP6teUhE+Q4vEulX6dT
4zvzBJE1WpfwUsM79aqjUNB67OaEQGIPifSTWvuUwsoJFiLNkXbSatKR3UL6
rGlz3iMaWT6SrjaJtrCiieaSuLhjZngMofX4T0djKwJ7frFbnCsPJXiVQPXe
jwb6PZRYe2BvsSoYtSGj51VtUvWN5+IdyBspwccZ4ptoO9M1Xw8utEVEXWX+
JLygDX1sM88KTKubYaGk2HJ2MjOBCVSPBFJm1MBhiKSfwOUQ/PbTgpiyGbp9
t/tbVAxVkUeo4cOCDRKjtWBI6GUgIuHllPC7D92m/p7kYyHmbW5aHEal7I74
rhohpQHeFNDETpLk/c1+yyvrrjCZ1wvWmzCcj92RiaN8szWW8aAWkc+GYE5u
4mCRzoaIm0DuXC5VmDnhhCUmVJJeUH4Wm3w0co/1DdnD6jseYgXHs2E+KyW+
WWrFrkQc7URKLbQri4Gc74d5pOJrPKZwlIzmIKfl9erxz+YSE56zMScW3m1A
EDd1C2GIDAh1VHJ2ZjI61deSUJl34IkMrGTxQLG50FwOd6kERS59G5L8DV73
t8Om5xglMb+iQCnzdLSwpNYp3AT5n5JnDcWifEXskHiOZf3pjnPEolRELrD7
88H7eu5PeVmoMBoGn2YZ5SZe9RSqMDS9+96dwdpatuuNAibgzYx3zQXyH1hu
bj+BgieqxvVq83HP9/3dvYYTPr/p383nhwlQR//8PIVLX9B5oncxXElOcEjL
3Kb+o63l9GYrvyO3d5yFzO2xD/b2YWBAygU9pApmtPfh4hJqJI/bEkQAJXbc
MSDaYfjCec1kvVhfiYs2gHhkRg+7QO7AbZDV36g8ipfcdxIeLIvd53SRbhQ2
i9cA3+XVaYMYCVsbrjX+ROx5eCayYNEWGmITk3ylXvGD7QPVR1omboqjw2LX
18gO2nkLdhOfpQBX0t+BYCJa9qIoRagpmNTHqOoKNx3RQAthEQj9N1ce2sqC
1b33aWVtkbaiNQK/L0y3YbrkdsW4+HNu0QgowG8gu+l7kqlhmcZWo1scWbc6
9ELPJdCXmdVq3K6xuTSnHQmnuKZks+967wMUGEIYZbfI+IxpJAQ0UhrRjKg9
40Ky2Jvy3YjtxSuwcxIQF2LFUVY188XzfuT/yY6Wc04lSoG+MX5vvd2LfL0k
qUu/zjAWOtLoI3P3j/yRidZxGG5ui4kYk0/eMA/AGYcnX8cM/B1xxibfpt6g
gsAV72M82CHTmMuZFzTDpNgFVX7UnRoVzaKEXrIBg8RhqMOS/WsM+zK8Py5z
1/HCTB7aFBKi/ZfOsvl5oi2pvAloiubTFIVDAgcgtIo74mNLK4U1e99frGtn
KHr4waeAdRlZXYyjk/aqLGlNfv+bvuaDbAFtUWK0GNi2Bf4hmYBeRG/DUMvi
GiUCcVH38UygD05OGcg7DaHK8+p+vvsKN6qsDsTQ848VSAOE0TNPgIlsgQbJ
thghbaiBg6ptGezp97xkHHClD931eWJYiNGTYChHAJuGVFvyh0LG05H4PzI2
uKI81BwQ9kQCsJIUSDY8wWp7yTLKRGYmMJ/Nquj63njG4SsKgxX+VBD5/YsF
uZz6NJxYhAP5/cyH/2oE9MfNYylRkOMn+11KJQK4ANX/wTnGMeqBPrvEGL+K
abMLxd0A26VpgnnsvFagBj4nnLG3mcib0YptooYw0BnoPjSL2lahQ27r3jSm
inr5SH9LSUDnI8dthFYnBN9GJjqCk7GWrvj8zruWXp1+Rho6vddkRvfEdSaQ
/qpAz67YmPM25M6ysFXgHDOXWEom09e+Y8G/VKNC9H4gVkk3ZusFRXrrYiRL
weBvC/ltIQEjLeeOQGwGgCbQh+wiaF285ALUojWRu0IuPnP+ay9X3bYOnXLI
Nzq0HD5tSCkFAEjXahQEASWQUAq4YgIyBcQggXLPSuMxgcO9bV+blnGL/Jru
D3t5o+sXzO5u3v0U/UI7qLZNUApvgmZ8zmgyaVp4Af6Km3Z/yValUkAk6Zos
RNwo9+3Wy1tkEyDEq8WD0X7ciosel5qyRXeP4rjeREHMRWhIOxnzwvUNfqjX
kn4Fnsdy2C/8QN4rZt+YcP2zAX6EOwKzM9pDj/MAoZHM5zQ/C86aht93geGh
6a3teYoMR0Szo2tBIV5LUhk3f8Hf/gM57m8JeDBQl5cnjkIdqsIF/BI4FSYz
QR2GbLXGUUqy6mFukTRRs5qZTimY4l5F8Bx7WglMyxOK4gpodZS2tfWo77ft
SGDajEH8pCZUOIeLZFIxkDjXE2bKMr2p7gZPLu/NJ8wPNtXdxxz4Bm6bGIY9
fh57bEFru1MjGXjQcYpqv41xLA8hbGl+c+BuRLEvxswYK8SStNeCa3AvP9Eb
7A1PJozOwJv4bnAU8GBhEuDSRfy6lJJk/5j6AAgRhUqw53autk9FefWsp/6U
vpru+IOS9DbrFh4i2NEw54s+IwFmBhMqDWVQF6kVHrSDX/Lu/rfYIFE9k0x2
Bl9u3rwamzVXHbNozvC7kZF3VIe9g4qiWKii1wI6v0Yxxp4zZiTRqt5Qs4ea
R/ua0dEIRQjqogZ4eBaIiFamIhmWdg71LkiWUfUIb4gPhRKlRfKXMwXjnCtF
T2Y/KK5/KW0owBLgZz6EQDKheejKJ+a+vc/85ViwOR+1TMECDgmQUgimP08r
QzzZOljucKFnchjsMGpTDrKrtX/OJ4ZYjJGq2zScf5lK9mhbWDNHdJKZkerc
BIDita7S+3d5BBFXCf8mWxo0hW2QYjp9hKf7ry49dzAY/i1wCF6gv6c88tVo
H3gs4yTvnDRJ86SDNDHXMPCdwI1dIkRAHDCcRNCyj1cXtS5Zr7bS5HHBy50q
DDt+WH+nPST0RxIJW0cc6lnRkeNWkFwzv85zQDbWqQMOh3mUkAsG+cTOPCFI
4Za/cUmoNhmcAPgG4oIYErl4l2Y551cIyvr0Z2siJZMlEM2IWLz++1zPYdX0
eSTME2WOVw338asx2hTwk/XaF+az7lIhzFPi8wcVLQB9RvIKopT/foWJBccx
q4vhJaM85pRGVApSZn+w1gKMFf0pJeet3gtAT1RqeSSgItCN1XTX9TbaAmv3
WFma95FCFtgtTdVZ8kxmkoxVRq+wLhmqZR/Ls7EfU/VBOfzrwJu5scIsoaHT
nFyRQqqOqV96QMl6SWFZVc0n8wt2amjD+Damc6AAb5KlpCNRoJMfQuunAYT4
WyDTv34fRRr3pvG3Y8Vt7RjbKnDVK+PVTCOFw/IURvmVW917Il3Qi/LdjVfl
CpV8juthY1GEdyjlahfX/NzsCBc1oB2zGpOIrLb+f8s2JIRYQ6w+kbTl4N7W
evrtpMQ7U9Qhe0WiRBdJE/d7UGYiB9ZFEzF7NebaWIyI0ryyI7gMDNQIE5O+
yLOs7y2zfwqXkCvTfm7cHdtWXeZUrae/mXElSyVD/MEb+CqitSYeqy5q+iET
qwPnMnwMapeYw0clh18JNtPyAhrBkElQ5Jl/O8RLWqj70qQpOdHLHsEwh9pt
/W+Tb7DUVuVsh1NmXNadatfAvHS4cVeyFYa8oHGakn4EE/YPLxPfdIj4fpnS
9FySzMDivOEtujFTPBOuXKlohHt2n8PiaP/kkAhnv1KSVoUGwXThz1fgMgrS
cflqFTcmMPBWx1XmqGlAHwQ1gifvPtAWYO3MJI+fl53NW3fgCi8pLuA9SQjS
Estff+TSC/9YL/aYLLd87Dpu1GzCjlL/f150fNw3WWwDwIk4S5hZMmPWAyST
b8hjzVnIBK9gI9YgHIKV5qDcVUxm5uNJ+lXgna1cMScCSw9kySvmQNmb9KYC
hZu4ncKlx0upqGDLi6wkWFMWn9w+vJLPr9wnFfZ/NKeZH04HYu7/nvjvptcD
AHbYc3VlJz8bE+Z6f+/QXJhudaYknB8bITL/kMTJAtTOOoHZ2wEz9mM+l5mq
thY9whcqli9TanOMszj1qqdhoNjtMA169wdtzglLQbjG77bCS+NrCsjNLguS
zmvTlGni8GrEo/c38gpqpyJAY4GqD9h9ukeK8VK52yADBEg5yQVRvv99oF5R
vJGYgpsmiChHMllcSEy3JgAfCn24IpBCsTNqGcWe8JLnwLvo2130PuVv0MsD
fCGV00fHZLlpf9mnZBJ4kXA8T0T/Kjid5MeOq3N7vV6yiuAUxpPq57MetZ1K
ZLAEjhNsJwWdWCc9zMP0oa0P6OKHkVWtZVucxhsJpIkYRZ6ZhVUTRzqSc1QT
htYAh5PTLvBUsOrh8qN14/QfIOmoZEyJpiIMO8lrXn0GDQz/eULBuJ9jZHtH
/ArhFoENN7dDo3Cd4ZLRtsrxGWJBZynEqC7/gkJDLen8X1odrox/N48J89Md
sR+p9mqJrhyKdrJhBozigVghwT68Zz6IUg7/3zSGKZl5J582muTS7xQ18aKn
+5sCAwDlc3kIAIdeWsBOmL864x5fHvTkb+hPsJVDED24D+A/nNJHj32dZRUC
ehyqIRi/OIFmT5Ho5/VJmhzhGtUZ198oMBEB5uq4R7Km74n6VKnEQpXMQDih
wsz+aQ9OtVPmEjxWPH8zifRmP4zNzR3cmQ1vKsKIoO3k/1l6HCW2EhKU6hAf
wD4Aw3rM7CJRT/52Y7GvXQHvmwdqxWoYzUmphRmEIfqehv5BTtelOCfXpE9Z
DcmZZ8AIdtebMbONb6nSYAR8k92lKRNK4r4nN71n1gdiG/JE

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzedl0faWdP2/Qih3ep4KiY2vZqRsMyQxEc86Xmw1QgPNoSa6ubbjsw1+w106Gx2JUKt9vglfYs2qk3M/tRqxkF/X7oBvbhdFEzr1FOt4Sjkh/lbmOYMmgZotE+/eHdpGZyTEE9VvaaHA13swv89q7PxMAGWXVLNfjuPQK5Q3pXhHqIoFeNw6ursG5yfg9w4S2XTmFSshp3/aMM8Y6PE+S2vE62u0E6IZoYZawY1pz5mozvgej/1D+nVA5xQYlxeYoxhAkvLiK+RvFzP4SgGd9nBaqOCe3kdBJFVWPJdHEMF9jSn4JK8nlgVgiYyYSIFQUa/MU7uHD3rp5YgCarXNXKV6CkbxadlN00wiEENBlABT8wBa1yUXlOr6o6B/ZK72gl2/TpCLjfqsCL2NUKZavWqtW1O/2evZDMe1hrr8FOCH7/DmANkUHDTqVlXM1vFXXlbSiF3Msu2SGNSbGIFMexOyOdAOTrx6WjFVxmqF7gZYdoGkIeQLyNZmarRIiNlLVrNIKyLcJ5hi3glNU8a5ZnzBCVmvVtlUHkLNpm15z8ShNaIIFNcXgnQxPg6tN/Atz63d+It99j9bjCqs/q3Cnfoz+vA6MAE1Ke0SXx9tc6HYy8+V+WuX88jd1EHggPaJ9K59pL2Q/kqW2VrQIC3oWc9qUyETaaJveUeFzj5OSFuxVcB5iWfcIrSalwkVEh1gh7fVXKt1357ONnai8WukKvOGJp5OiU+5BoXQXg6kPXM+3cVzcM/icG4AoI8iE4DIYhzNMBVNDR7l8kSY6CpIEOQ"
`endif