// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tUk2uUgBhlQoIJMCueEz7khkTMfV3LXU6rskKYTbuIjoKmCJ7/nZI5BlzDV5
aY8t4ltvluRYLx3NHxiYTolzD0J5Pt1P0zJ8sQ8MKxqg1cE93GqM+ccU+3T6
PJi9XbC3z57DVTHfvf0EPt8YTyTuSdRCjwYuuQIte2RpmQlFZXEwqYuel5GS
rtlo6wj+uABtuUbE43WQKNyf4dNZzoi1NbeRPBv96nnZHj8jImdcMWkpz17o
FKmVHOahRsxLRdXCih7fenuNPUsjASL3IneUV9fefP+NYb59mnILm7CXcJ+o
3/5g69P6U16y+J65SyjVxFv3+bugR1xsvCr53o0AGQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pzhdMp/xLmPfGNnGrDsZtdLR+Xf2cmdNI7xRmcWNceMHyJjbeHQIOFk+3lJg
+4s2rl1YYJG0aRD++jJCjBKeMjk2tDVF/2YB1KU1FIiqtoJ0BI/tqzETwet+
X6US660AGD+QGdQ9vIyXrcpBeRR3T5o739BzyPhmJHM30+ZRbNTHU6s4Ea4j
TM/SDBN5k7TEGIPYuLQX5yZKqKGVFtOR7rUGmnYGnCLrXjJMSAhf3YyiL8Zc
T2QTTMYQZ6q092bPlMETs4MJTx1sc1y8hZwdrc0G4aaDOxMT4ZFuyhGORcFJ
j6sCwWxNvjzz8nEHof9Zic5QFeE+lD2j4weMRIVvIw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DN9sZ9I4DKXab1zuNOl68MP1fDj8Ye6dA0z9AVJEZEXnlJP/6kRTE58wXu2l
b7SySuBr+Fiwj9JTSifVkJmW4zYRT0dX2jzRoYHgS0nQada7l4FZ7K2qDiiy
vh0Z4unFx1ZhdC2kDRRwYMDVJBSPQ0jhd8sgSzRgDgVa2tOAkEy5N9PNgTbU
Uc3E1zQZ+X97G2GlXWdJP0J6MOMxuuabRWcBYDgrZL7f4mfcmIGwPE8eAZ4Z
Y7tbgrIbE9jGJy0EYoPv2CTAaTkdm5V3IAA9jBOSgRg3xrGY7lzgRH4PzaNA
S8zZ1hSXZrO7p3XDxMvvNBOjZq3uE4OGS2mZ+0H00Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oZbPIW+/awUdwvtfRud2jVYqCs9Mf6x7MW+K1xnxj/JtATC/LGhIiMwd0dJL
le4lxIo+DucmMzBGDfHXM9vmbbr9jg4pQJeBQBUMDGnrcF3nw93RJFbeZPAw
pKvfymgLvN9dOTkwXkIcmId2ZI1+i6PoqA2pn3BVpymFDSjvT1LZh7xyj5KO
QN+9DixZZhuRdhulxioMiZUYROpCCjPXANVHXurToR/xefJECtyQDW+vj9AY
vOEOsSBAcVonzWrR4GsNOQIysGWlc27EpyMz5fo9omtFs0P0AHm0XYRF5hrW
SYNqQGKGBr8G3/MvO3f1A4TdgnH8JSjM/vY75vg1mg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rtwMuYxnEPWkuQcJvQF8NGDM8oFFvBEmEHmamwyJKJeInY8b8xE5VNvPRijU
PLOnI2Cu7q7w1efzlQHdRxS7uJ6elHuKKcuXFJRPG+IkN/3P7YqhxQIz/MLX
pbUd1L1DnRA4X3dXWhgYz0r8GDulu5DBBrceXrExRFrr2dHC71Q=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
rwDL3IM42/PvO7sJZxnj4ZAsnQhrGq/T45oxGeud9qiOw/GZYZRgACS3ltJa
hiLi70FTE/69+/day4WSfon7bHVHGDX005eDWhtq6XWJLv1Edd2/Q6ZjtDj3
AODDLHmiMDMJZ5qKGb5XI4pcPHKeR9lDSSMYrYdkXlCoCgrBcpBITUcQIMxR
D3hQ29ve4DQ+MZgHDzNjjZkPcPUYEoJN3be2BjZ8+sdgKml6giZ2VEROuQ+o
wQhQ3voNwHV1E6r6jLtCoYqjmFxefBSfIk5KXsLbgq6yG5kHJuDt7QJDrOxH
DokM3Iw8QBv6r01viKOc7HwogWMnECxkai0O1UIxZmtoRT793C6xTDyXxa0t
g/5ivYL2i5ZN9BSF3nUpa3iN6jVA+LuJrS/xYcuQ3A+r92hFFFYaSP8+Hlsn
Q9zNWt/gf7T/WGOGWWBChYqL0YPGt/U4Mz+HBAlPseVX6wYRcPWswzYahNj2
S/215rt+hkNsv9mKDcTJyTzZp2MUY6RF


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VMZvX5Sf3pSrIMqDw5LdWmVzdEW59IChvr+zwg8nQgn1NIKyGLgT5dX7vaJD
bYH1UN7VMe09JOUgSdJ9qW3Quaj6TbIJ8+FMNYnY8G1+wXDk2BLeDRl4gwU5
ufumV1WT8ZwthijXKqkeJfTi7GPu71oEJnuJ8Ia011kFGwd9C8g=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GnnjdiFdcz+VH09FyPU5tIxHyAibtA5fnUsJ/QbnVwsScPlrMToMy0IhCYd+
YRxgQdV1pa4KmtUOP63GPL8JTQo5mQRtDczcndvro/7z1RRI2fZE1rxRSlHg
ZGXN36SrfXIXOk1kU+SsZtWP6eOEPHuFSwQQkUaWtl2nYyz2Zgs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 79776)
`pragma protect data_block
rU0gyTOunqkyhwzrrp9T3hUK4Yrik+tuJVRT53zhmIgu30Bqm4IxzDXebZ2q
Gkjdp3juqz3tyI9OGCHya+PNAkGODDLovmmd8tk6MUcfqqvGRu8DdzJpnOfF
BZ0q0Dw15pvSNQerkzLY4ZjT+hlGQ2K5GVHTWtiObPmv13yi5d6GkmLSkhKM
6foCaL16KFNWZOZR4uLWz0mdeCc4/0IldiA1caGUFy+PUDICuQMSAfv3PFgA
LYPjr/eNXz368Q/6rc+NAHGTQ1jR5JSBxmxqmZnc1cNwl3YA8Gh6DwKhQZ/W
dWCp6LxnlR6OMd+KMwubnM7yT5C1d1IpZ8XC1tKTAWCNlYtzoi4zhkYrN9pP
qbldgUfMfKiHxpsoDDHtiX9Mf4aWZ8O50doRrrkDPbt27QN79SheOznrK0R4
4sRsWofHmQK2k3N2APrCi8zCiFHyvgCitWFZzauTkEYwDAy9NnISwy0I8HFT
ugsSlh3qYTtUEvk2A8S9dg9W3nrdI0V+TOuFBHciKN7mJ8uTvv5+72st92zT
xqbrUI9pYuQhgnMtm1lzjGWn9Cr/GcYu56jC6XZu7hlF3mjFzl1IN6hvqT5t
OwL58bW6UU1qJil3vLewDDoBcjWCOP1Q/5kZx3wrht+G94sfMdn+a0coAsLf
+oQb0H7NejPI7MrOdL4IGAhLKafHLJOqF9lNEU6JKsGhYCfQ7yj7senlmp1C
0YVzpmVkOgr8SfpvGK4sEKt26qc7i/OgK8AM2R7VuBDQKTivAFD5Z/MwKWNf
xU97k5SoKaxUAXczopY1dggKG6DV/WqsFdfktuxDmJF6t+Hd5MP2LQ9WC63s
h5Msf/hXOLnpvP9Hj6P7MZlKs0lGVOVUuZj462/0EXMf+sKtSw2KYOf6nynw
h0u0k55bZE/meC2XsBshcWbw5o+Sw98Rda3KFtSBZYGnEMqhXjDbb2J7OLZ6
KpEI/mJgxg1IiDOYFY95lDYEPWOaCW6hvR2eMzSovZk4aL6oPOPAPSDWn1Zh
JNNZUAeP1HYMrh6ci/9BYr9n8UdBAdUAsv+CA5yguZc71BZR8FRaB/ZO21Fg
wVR/75daA1X/w8/f+oVGJmVbFl/3igSP2shDN1J9vFarnD8LrZUo2opy0oVR
cbYRmFqz6RkpkdioWHDt+ZV2+PxrCP4vz4ceaC0077++UiVfnsCZyAhhPPHV
gQ7mtmtmuANapzWG/f0VV8ja800/G9yZv5sIdlYy4uwS1W0sugSsbo4s2U+B
3V/bdJyDtpVhiRocpCMVS/JXWOAZh3DdyOXIVn8MoF9hqHo9fzIqMk4uDDQ1
X0rsMRaVEJ9Xc3++LBH8RK3PQv10yEtQCR72nt8sDsWuFWRQCLSC0cAzSURs
MYYLrk2h0EmpsV2As7fxggf1VRZgEHJuj9MpMQhVM3MZqIh3UsQFTelIGU/Q
HLNfnAtdm/Xss0xu3l0uvnOFXZXYLuhnSFvs0JrOXjD9ll9krGft6m7ur40c
zH1O8Zw0zuWkWrjaLVDrk2thFVFJJzsCRZJkiA3VD/tUO6PUmEUgvLB9fCbb
2WfbVHkMVYGr4mUjVqVKRQHHNuSn46DNccDl2K1kvFTnTdH9Jy8vRxE2Laej
NGPMnRJXtaxo74r9AzoT9v6TXm6WnMPXBNWbFJyLvVY715R/bCPlp8S7nygh
0dUAQu//8gkXXwF/kVm6VWNq/VRvGNraz5RRzBuSkSTpVhyllvT6G9uiR4Tt
N+dTONKQPUeNJu/aM7GUradid8griziOJQZxz2UgV6Ft2CyudVRSewXLbLSC
4VVnY3XnSZiMe3SXLT+7U/xwn2L9b9ct2NlbeTc/cXdgFLfAbfRpQhUk8Tk6
6nYHH5HGNCsy+weN94BXYHN2uX59HbbPbdMP4/m6e/haRkOQaBLhzdHlZMIs
VJ7tYs9cFb5PPP+gt71zD0GLL/IF6Hk4jygvz+t3z1AmHmSAU7iGiYZP8b2h
By+1TcBXr0fiWQk14XUmQ6lBwMvao0nhGrg6o+rLUSAuzmEGRo6MvKgOEN6A
mFURs3OxDZuaBHV+7LQviaO4WiCuC7Ypux78Iu/tc5Fva4iBgiby7HcJ/keA
8ftQNpdnRzfxBdpsrT/Uh9QDcehCwwOcBjHQwFpM60gLxvFdEsP02Fl+SjWG
Wa193pE1EJHbPdeDJUbf5fMQneLpEUoMowbaPVGA/8m96bMgPRfP5r9i+D25
j6Bj2We7betcwah0kRzHt2Pk84HkFKrTaWXXrRnfrd/hLLC9JwzMTjTgyyZN
eRdBu3TcDor+rQuHXeyrKTeW87uCVPxB09hCcZcz55/g/eV3gmyunzrPpggz
46bYJHa7DkaGnfO7HAFdwNF0ZSmx0X/5MhcOjSAnQpxqO97V8bvXDU2QRlUC
bTSIgwwy4yZ+Nxu/7dP7+JxWnZrKwCFywWuD9Yaf0Ww52RpCBbuy9NpuI8EH
5hfCPZAf4+ByZo1J5p+HogoutrbtVqJlQ17TG0NEH9g5Hyn5cGYuXmZVzQhN
s9W8wIJUMBQJHQSX0z77msf/irfohqK9Pu9TmSKvu4Pcb3OzYkwi/+ssWheE
jqfB/Nxd1+LHXnFj57Tpy7hoydl+vYqAuEEARjP81cRNhivi0rTvCo5VAQTX
SesZ7XDJjnVPl/9DtGngyiCUTUDI7UIY4KDcQxewsdBTVo9rVFpMV59eeFK3
tUF4+CxgCUXhxhPOzQgnFteKdh++fuZw6+n3YDHCjcD8DfmMdCds0jKsecA0
P7WIyBwnlfh9KIWT5yHMIyMYU/7ad+bRl8McB6Vv80WxLRVHIOPmNVLrvuGF
7w87nb2oaFB9jakSja41kMs3gCwXbTAWrObJdtAJuN7nz2aK9JoScom+Vctq
hvCqoinxzq0snAswKy900Tnjg85bAGH1zouwZSLbOADYzRpsxeXyw8kVJNH6
OSqjBPNjn2vD7UaidmtJ5v5TNEqrufJ7H8CI7z5Rg36gr94SsxLzJFKoB9S1
LT94EWgvPnBdV6gSBPVAizWE42uQGRORwj3yY2uK65LXvqqBXa6O79cBE+AY
l4oDy3w762wBTT5fndbCs+rk61cvO4AorWHoHDOjc4xhVVt9AZ1XllcBGYp0
ALKN+c9Vn8IPNAhTY+NC4aT+EyKVIc+PRinkrhKaxDkf0LlacJ78Xuyl3Nex
AuId41sTS+RqLTcIa0ENYJB9X1xFKPLT++oE7eoeMMzu+wKCNZS0k4gUbfpl
TwR/uyJYhJzVHyni6lYYmDkYSYQFKte6NM+ZZmAU9aC8sWddnyAKXKQ4SCig
swfROWHgiIvCWlj6h54J63MQtA3Hysf6p3PFvxqvcdYO9r/KQpdzc5ZFzWD2
wvkGjgdYzkCp/DJjgg70K0xQJHMkyVj9X8mPtTcFPr+qSJl+VYM4y8aPCb5f
6Y15aylW1BKwh4GDxOWQ7HypW41DU9aunVtd/VFvjHRrRAV82AI0+MLTsqtb
83HlrY8wkkYQ1upyHvCQSgqhGZWGWhyjmMJfzj5vAkDT2MKXb4cV8WwyBBuQ
XVfQIBFtvOSHtB8Sq1G6JGFhqufIAkwIhd6pi9RUu94bYLB9KT9T4PjoQLJy
IuC8pq9xWIT7QqquZGQsPp38YVZoMecBvO3BH0b9Lr91WjQ+c6esl9kud3vR
wKekotujE4WVxvHmz8SOLnQ3S6jLnbvzMwIbGJBUHOhlVlnbI6hRhpm/Wu3O
MJS4TDjYSER+4lcoEIvfOV2msUXR/y8/Pp9Tuq+rgu/quiJaWBwJ+aFspkho
/lB6jkdAEnH2rGU41GyR3i6KJSTfADWPpF4HWVon80RypuBNZbE8n8udMeJg
3yjSykc5sRrn0548fLkF9h9G1CCLxAWM2Iy2mSfbO2J1g9HREya+uAywZWk0
q365C6owjJdkvF8aF4Z+A1j06e/wCR6Un/VKVjjgu/cLY7xgsl8yatm6GTub
dHtipAIw6c6zKHInoSRy6pFNUiOyi2CZrE3nM25qd4EqlzwhiNiKn2G0V7bS
KX/9ZwUF66akaI+RXNWKuj3IgjjtWDe/DF3ogtnuQpElOGnCmGaDYrfw6Grw
uH7XjBZQerhMAc2kv0cCuRHllciBkK0qNolx8drQQBnxJk6s3rOVObofoNMf
t/W5FP29ELAr3l9HiliQaLEg3iPdLMNFst00OZr7RTgBLyHMIvONj6C1QZUA
QAyoZv9CELxYEUQU1Mr5XdTynG+ouCg/qtROCFUpgyKR81utB8q27klKTHfl
HaXTIJdAYhzhuAlu3rCvlYH1RaNkYfTY0c/DZftqT5XuIKnGgek3RsRrmijb
eW973yqGT9yFj9itz9hZIv3CQ7Z9CGAnWuFDFJZz4RfVCTZX/yCR8v9X3IHT
gayC8wCSbaqMGjMXd36hT2J8YLp4UBghZfLYAyAgWoaaU+bjCozubBV4aqGO
v5EMIg5gcju3gGAOcwi+PEdMreoHzxeyJYHmiXjBdIZt1TAtqnTgx5eXNcdv
fKSSt46ESupUmVBhQ10mTAnhc7nfieIkZNGB1dj5X1G19UWM9qm+qQA5tnUu
LZKkXp8lKFRCjet40oYb3D6H+LJv63FW5xNnCtTaRomhlNFz4dZ+l7wnFnGD
6mwG4+ZAp08BzN/EQ1LDInP0Q35bE8z37h0+lyPK8dgKF9QHwE+xXjau2uFS
JdjXoiTwSleVK6qMuLAeKEk5E9cMkmeK0NlY9++nHus1ayVHcqaSt3P5pcuS
/U+kAGRlR+G71YXZAZCS3bRVO42QAyDtlqZjfK6Lw7shiZHaZHaeQSsb2MDf
VYBNCW4oyiUNdSNZb/isiGSH8iiEJh6wvzPUXt9OVu4nS2UU4fIRwwK4zSDO
rTY3ZDgjGzIViN3eS65UFVF1615YQmxJYASg2JpkztV4KOgVbpvK5N9wFL/H
08q3GLMexXZAZzLZrnGZxNIwyt8HoR4EKuePG3pV0hEI6YsR93ZNuKfpBGHt
7dCNqhJyWBdpuyq+2V6mJR4jYMcXib3kPycKfR2bXDjNBYT5j2THNg2X4SOU
vLugnnC9Z//POofrmZGBuuepMwida/8Rg5CI30jBl1jGkQpqrlIIKpXpHyqP
iwB7alRLUS5tHv76KyYGGMqGqDzJthZ/2hRhTnfWf12pKYtTahNLYfqgMI/C
Dlahj5LrQN3d1oBzwVYLOlto6QNgT8V6Fb9lIPlvdD6VJ9L9SmI8/VaoP4L0
FiDHdM5Lchs4HV0n5V6QEdivTRWpWC4b8u6uBXfYHYWTekZZ1r4PLgB0XElR
sByXUq/TOP3068UFiewjVW9EgZtiZEh7BD4w+dxBMaYCv5xzdTNkcsBaA0RC
xwD+pWpzHduTNTEVyDd8ErtLwq2SdC/CWB6SgFYJBj3O/hUUcfoym8KMM3pt
BaY2rzavSeIRVJcL9ejnGyQ0WF7pO3cSxxzLyJ4JxEHUTQvWoJZigK7sU4pF
zvyNCc3UnQLlpDJJ2F8v9IQeL87ixAtbeg51epHalVGb5X4SC/fchsXiCfKW
UFecrDzNgGnVLtHJcZf0BWO9ivycDb4UJ2ek1wsZ6hj2nw4hhk5ene7w8JIi
Y19+mzMBck8Ifgkp16pqoTCOTYu7kYWkuW2TTNrb5lxusE2j0ouNB3beTnPK
NTkRy0Fs4U+hyaPalH+OMzAU2FoIFQhRTxXO5Hfxhj2um/drd/CB6sCvsfKa
+iCqoVVNzB5wtCorSfleX2H52UuLrMboVEGFKHQlpQvpgu3QmSfjjgKCbbAx
xnsjUE1ck/S+E/tJ4Rvg79n1xkNvyn95IE8Wfl8o/dkkqhwKKYDjwQNXk2cr
cNfGA49qRZK0z4lGWgIJg2KDzq5lpjYn5BkWjO0XS1yIJHvXyJeSRDF6KsU8
OiCV95TIq4RKv8YUTuw35J6DP7hMm/uRZ4a1Czuab8Vzcs6pE7CWoTxXxmD2
ucggClrE0zKQXaZ7sk8qm/T3BB16VX/JwUCIq8r/n9GPUsAK2H806FLx4UMD
72whUDq48n67f9vTN2b1Ic8x8jQFxm7vgtz2dUo3631WjVeKkAZ5BG6ZZG02
epVmq8mTWInqFV4Nn/McfZRGTVncmrOfLy5CFSbNKJ0CvPg8zUxsk67CV8Wv
ei93MKFLWDATPs4KB3bgZ26ndSGAs/qGbJJa47y1tD9d8Mg0fXJUxgbuYhyX
fz18aJxcivyGYKVawKPYYmYzUL7Kfz6zvnhMotr6odDpzUfEcbSW0mYHjf34
EEiP40k0E3jadKfEmAooeY2cNgwtcxMJM+402/Xlb1LC9q8rd07mSiww+9A9
I5t0nM77vURIW5RAvEF/48Lcu0wR3BZwyK6Bez3msqgQ5fh95jviPGUV5pHr
BJO7tg/dhRCINk7TsdIZxz1RC6ENkMAqrLKOkW+L3xn3yliqBuyug/H7o45O
GgbY5vWKKmWq7f3LO5Z1B3oN56WpFukNh3x1vwve3Rwu6Yn7rkDl4J6Rp9vp
6JA+f/3oD51Z5HscsKj3xxeZrx8lA2xTqUHJYWxHU8tvKzF/XgW3oH8WlynD
xvUFpnV7VLuOw4eJd+RTTAf6oSD1HShCxxJyIflA8ttU1sPZcx2D+XL2m2lG
LsSGKB2j/x9vBsY89yU857PoZzIVbjJTB2XGHd9fYslROCfSqHZik6oJBY5P
koRT1/r9WDbSAG4DEAg1F+qbZiqY5wRhyoQ9hBXq+0AdnOji/bZPKwtmNnNq
EuwLabDet9KxdbTtr54/wyhjxyW2o8Bb7lN78kwtRY/eytX/foKULrcGh8Kj
RB80HpwjYDj4Pt1uA4CQ5kUGNp3pJBWcON9kNIWz1OV46Wu19DdgO89YVeM1
GfjKCt6UPZb2b/18mrbQ7bks6mN4LWIIa/majkuEvxg9tG+fJeIVslYhDzS/
5YxVHmR5vcbAQCnnC/F7tyYTRNOqGU3++PTlUQCRdNtPiFDyKDmj8PlFiPvf
zV5H/cjXZYrnDt/K6Z930u5quzpFY02rWuD5MMRIIRCmNn4B7JvmurRnSJ4Q
1kJWzuoPRAdqvsiHDjD19VlAzkCkp2IHr9CLnRL1vxlbR/X4eu1Rtvij8/SD
l4FWCpMEHJ8tehIACHxCkDr32J4Y2wTPE9m1NkDR9bSSLIiwoPQTA7bAOOSi
znLv+Q8rg7CYDgMe1k51EfwJZlmxFJaTDPBoK7b7g0p69011aXAPyESLZGi0
DsgexCYIfDTjvDZBeNf5Vt9UbiJxOPw9QJ+oxpw73Vuqa/LrsnIQRld4P6ju
3X8i4DJItFLnSr9929JYf1n4U5ayXVck11b+2AooyOg2S7f1+bsi0Ra7vQG0
eES9rjlgh8nAR/zylUgVr9jypaOm4dzejcnBG9b1HpgUE1MKX+Oi+hdeTogt
PRogtaYJXW4MW1miUqFVRBQ3tLtwIQIhEbD51gYMMrrBqXu/rAYmT2Z2QQ3R
jWiSUmeVm+waGdRVF0OgX0eyvyOtvyGJgq+skokBKTRuZ4wmH2YMnOyEmLik
cW0o9I9PBtlBve2Hsi0pAAF6DFHbbx6GoJc3/ZedUzZcyhDnVzvBgeuwI/C+
9Nv+QpXk1cRgaIvuiC34qyjuwMWwGKdOCj9Es3rjFG+L90vJvYvfMFNEs3b2
7yjFXtXDtBJBkQEEHjF7apuSopr5mpZW18dL8DihkzRO39JGZsIA+fizo/VG
jeDyNkuMptvwG5onjXkMvmo6v/0u/2Z8Uzq2wziD+KMbOxRgVhWM/WkyO74W
iFiCo4MS3yiDKzCyEJhp/xesZTfOHYrfu1UW2f/qJ+JPPCKap4+kjiR4Nuc9
ZcqiHnpEebCYmOoh+NdFrkOgfoSX1M0e86cMvP7yRLSiWfu7sHFUjF8xyEjG
g+SomFIg08dcf6Rd2xu9iHez9l0WF71r+OYBGac5xggfZLMeZYxFP4WLlwYi
xdsK1ScdjjUnUtar/9yCmzNseHP48e7+zeMBLJy1vU4aEmAqdnpZdMzOfJud
AtFmo2Mjl/wjZGAXMiRd/Caxr2fdj1nHmN4LH6qglESnk7Y7UR8/uukwp9GY
Rov/6gXcFutoe8nxmfiKQa/5LEEmnp7ZKvgX8U4lAb/HJujgGLSJ9rDdpOSd
4L8rQsNS+MCmTOym0l6zlX2uUbaWe9YbQGgizgyc5dW/1jqMbu+165BvBRkr
UVmH3+uoqKinyFEHyXl/ptUNygyPZf/tmRlxB/25T355rN2uyc5sFeVb8Gxu
XG3i9E2p/5NxhZ7CDEf9DGSXZHw9SQkJp64icGrJhgWSCAkPivHtzIHa+crF
8U7DC/ns2Ew4+E7X0t/SCvF9/5P66qruQIgjX57Hdi7uiuwGEkqJM+OZn8Lc
KZqCYj9eH7YajRzjgPRZBcAELHVWY46BWj27hrS24E8JZ/3onXz3uEHk0NkQ
NOrrKqrVX2QgHdmtizfWIoekuQ2U3m+4YJi+rZ+hmNtE8KjYX4qxPND/gG1N
8pBfW+qdawOjZ+iEolWNklV2zZs17HeeHOyZcHg2EUQrfiP2Jes2JPi9+C6Q
31SYgVK09cTbKTvZnwYwHv1yJ8VftOgOGovzPwJkVjgEtWjVX0dXLOp2lf28
JCqiRJIl2lkJ6D6bsXHyUZPTigBVPA09pETib2fv9ctwELdPwnz7CHbxqtpt
BWr97plUkdDMRPvc2E7TBJjZDdnUD/4OvuJlpyf7Z1wGkXs3qNRznLCJ/MpH
fLeTWDfzMcId1tXl8GPexOzppBC3ZEY0PhIucUj+P/D6DBGS5ptPi3KQvWTj
dHl24xkGngLBOXiJ0KtHuDbmc94hRMlbPSaj6ClqG5q15NywnE4JPzYKr/BV
wlKdD+8o+27e+Bux9FL4AqJa54sezrQHxBGz1DPMj+x/SArk+moYcKXHQ7NL
MJmezP/vhO78N4cq/fEhM6nh5VAwggQLbpDCmv3AxZGcot3XoNxyAGROVZZN
f69V8i1yIW1AS0DFeErZ5sZmNFd3AVj6iKvbKSo/nqlX09wpUIfCIPJ941TM
VnUJ92zVv6TQcYalgHgg9Yb7ziCdICFQA48occ8YvFn361rsvKwUkYbAxTOW
Dp++aN0FYL9Zxuk1AHHHhCNZxncfboyB22FMlTIZmP7ekxwjxTagx4eR+uGd
WlC7QH9wm63gVbdamAJ59hEqxBU3Mfl/79TEKavRz/ghbHQJn0kTegcbAw9r
hwOAw/aqVes1y7S2gBi2/POg7WXesB0sk5jXEjzOGnZ/OVps9dEacrmaWvw8
Adoh7RxHtTlFI3D7dsA5tMIQ7sXd7x1aJnWD596eYJjnb1XiGCrcsLjw1RF7
O+ubFdlVav4BSsIQZOTR08+URAuxQ2gAF0wL49rUk2RsPvTTQeSgYBWy/srn
bCpdL7MtAkUAShdxjMeRxos94cDTVeRFG6gsaCgk8Kso0ZrApJ0v/+6KsZjV
a9IpeYCg/ZMfTibucQI/Tc5lxtDayROs3lJfPh18LPF6lFvg5P7NGslnRE3w
zZ9EYg9jbYomrGFvJYPG/uLvTW9RoqFk0Q7sxgs6Ci6Oi/+5V8Z+KHa2bMii
PDECY7TGOL/OA90hXoY73h8zdXq7ZPXYApkCqPNaG7kVc8IGwNVHxd/pSxWI
mYEuoXuViUqzjslnLzhoHDeDIx4mX5EdI/9i5hEfhljTm9uTAPw/WLztJbxl
WbembVIOg3uYItMK8mmhrpK+f7giDEpNQClOCdIO7yoB9Le3jLX8hvT2ul3B
jSlm5WefzvHN6E+U1PzigzXBz/vBy/aHxFjPHhM8ZodnrMFgUJJvNnpnRH1A
ZnpzhxRKRRykASCm0NvbrMdzWh70VmZVu71d07v+KdDGmEH9cX6vDRs8ClQy
tR9oXOBmftWP6bOf5htA0BHFjArYKIJqvzX1N+TLgWImZdHp43nTBhUUAJF5
ABH0WJ8DEfY7YwUeC8u1eBnEA/OvL3KR7ykdzTRMrT+/ApEIq+Wwh31Hq640
ax2w0yV0vnvIxqcxdZaLXRM8ZizhXSHJpUupamw8z2FxBKzY1Fykjq0m7bhF
glKmdzsBvnFwlms4BZkuuN271NmSQJE6Kynzn5R73jpF6PDF5BWxoRPyKdG3
ZvfVan2D6zPqLQOB/CUC6D+Zh8cRnUA/fN4ZFE2FgoCyOjOJcEvSJp70H8nz
h83elptyoDj3buRHUma4XjEhu9AjvIKOU1aAmmuH6w2nSHNrT1FVT/iyHEtN
NLVUB0LdCKBNNz98u0xA2g1nPlVEJFKw4dNYyYxshP4ghxcDASHAwyUvezq/
clSMLumY8TvvU30rPRcl5M4hAT52ZuwbSQtyqtoRnob1iz42WzW+xwre212J
JtIr1vDb5fAHPH1hZnb63ODxUya0XLj1QckI4oDvAzkN5Qkmn6gZok7/aEXy
+XWa6MF181s8om+wjoided1ym1ru/4PEezxkBLdPFRYotaf/jWRBKt3mTTTD
6ouXTg3xODPfsh+gY3daQaGYQUYXA9p5FEHNIvMfo/R2nLhUPHfL37tCZ3hF
rPMFId6WsoLRwPW82Vcg+3Dfz8iCqsN950AZcjGfUFrL7Q6UhSxxii7ORnZB
KQg0gtZNC4wlaDiLo92ReWpH7tFlnHfETdqTDjoS9q3v+9gqB28OVSnAgFJl
Q48v47EhYTWl7VO2+7QXMq+cHVtwn4BKs9BOfqzeFXdZ6Oja+3GTk+72w55/
LRPFKSgp4RtnSh1U+E52BNCeGrP15Nc1l13M8i8WEo5Dxe99WlpPJYBm7+t7
MAuWedg6iy2Hq5wCcQBWA3Vkr1KBXeh9V45OEL03zRuMn+R/JPx7v3nqhmu7
8f0hbYGfD1dvvRiOgixXIdaLDscYDHY28cr5QDHQNmWizqdK4XKQZkOTkxst
eJzRFZ2jSkoOJubQIgfhsM1c4geJ8Uwm3acJUl8dDVPkO7swwEqqffZLG2Gv
cskjLxTU+UWHEB9kH/4L5cxBamhKcSbuVjGmthKdpyCmrPWTtbH9epMw694F
s5emH90aqjvRfe1gz1ZN4H9K9wVmWmocJzfNILLXkWdx6DNpI6QNiwGxaXGl
ZOHyjU7Sgif2njCCR3piEoVtMMjCaJg3rEDDhENw2IVIhR9l+L34nxdY6GX6
XAh2n6jkURtJp8X7K4QcHHahair3ZjY3XUG2OzGI1gEdClsVyvZPvQ/Yn/Hl
gI81OrqSI5sfB7LuzY5SAjIMQywOAKtQgABm8roLLq6TrCtvdtQ4r3W2El1M
v011T8CUh/eHG879KyWrE70ynvDweWzIl3MycGG4fhxibXaE8A9oA3eLXo7U
lCL5NdKwiEtBwgSQYrAvNYm46ZdP9U5muBggVgR78eL6+HT6mM5rbbA5RJhc
oi951TcQmS2qOCE18xglcWEJ+YjOjIWPe/mSVFBE4nHl1LVLR9e3D1lTyqMG
T992QIHRHaYxSxs79GWFiVeF8ux+va6R5PHwvwBIWFOHl4bzVVkR8MFcxCq2
jEsNMcBr8/Yzv7dXS2nfKo63cHGnwrpEmlmNePEk6huPR4+Q84KSU22Swxw9
MlUJjS0F3+uP1X130/Ely9h7TxyMnlwl4TYlCfSzHlA2bPGQlVBsiuDwMI2r
n4AoGg/XaarZEqa9aLzNxdXkuogNI1QdELJUbyp74nZIpdMys9yq3umkuDnJ
zSU5xaH0tFxSITOZYLea+EGtcQlRUxZ31NoiuYmDpru3HYjrTJI2i9X8XmdG
xnl5n+srnEBRAldjsYh+z3aXd80c0dojj+smgG/XUGHG2lE6F2o+AZ+te8I6
dp2wamfOjxS8nwnhN09AGIEVAK5RAhUsOwsC/vULj7LCh7WQ/2dW+2CJ0sZd
ApyUzJEdhO8F6pTdnOqnDKbIaolGq9ucySNtuBgxHnkHQ8Df6bBHysCsbmSC
nROocaDQhN92Q7Ylp8vnRuI0QnZX+V0qVAFpcR8FqaYPxd4uaIF3mOV3iq2N
pxw6vPRXEwwtGkEgo613sUiv6TVPwz57WTh9sEfiuFrS2dYu4xgdPDZZFoYa
CijAfxHHlZrTZlw74XJTmc0v2R2QzO/BIOqzUf02SdCVc/kKgTctmy2zZUUW
Gs0CzNDwqu8Vuhl1MqXXPru50JT7VYnLm3hFOaS0g3lDBGzrnCkDQIhPW6kA
rlXTQQsGEZ7ujEatVVeKhdGRVNtEz4nBQGBST51+pbcDg+RUMApXpxeeycaG
z4Rb5u4xHsqmD6Ty7ZiTr+PHIgDwSTTdJ5hE1JCbCbQ5CnG8yDZb1gULIBOM
cSjdQOBEOWABq8gLJWpkbjalH4nPQ0H1Tw9IKeTH7Nty8eG1ReHYdwHHIGFK
UaWYJfq52R90RLWpaOmfBFD5GePst5mFxn2vtfx9vSNOD8PVnjBh+eNNVVHq
mqWuLEku6ZEVtqZC/+aL7BXwuR/L4IxUZvanFa9Dt03VOk8wpE/Xdb0J7Jns
Je5J617XnXnzjEIuGpeRFvBm+EhRzZzaV7pf8JnZknsAgNrcs5fwpObCcLh8
ys3WfeKyKjGJmzVhjzr6Y/4U8MaHk5VmPYHG6XmKUDaJNGvXbxDL2smcv5fI
IXSutdtGahUuOS0qw0dFkyLXtA1YbsanrqtuT6dKCcgGJH0XSG56HZOSfh0q
QWiNzxq311nD11umWJAXPGcRZ2iOjOhfI8PPJb/j6ToBembbe9y/V7iYzyWm
wPkibujW+0fr6qE0mhs5kYsmcMCXRoHi74O6ejt16FJVAIO+8NaxUw2itlk+
zMedebztxxc+fe3SHznPRluYBE+m+WuI6/pIJFRTBZRjLL6YHzqFn6BIVQlY
REpcbZIx5t4CemJIpHEGtERK8l/ZUbTYUr0FzWcOWDhk78yAA/JE/hi0GrEv
PWyEZiWZ7pF7+5vPvGoTzM6EOl4u4AwoUjGfq1i5NaejmEPKCeWogDSwsL3O
/Xu8SKw7LaQj9Um+ONgdD3nDsa01XN+8uVw1VYpXvRShx8M9Gabm5ReOoMIE
nTqsoVM/+UPUxpX+9OqZBmCxkr5xHWYlSKCoKujLSe6Y3M077XO1YvHq0oqz
W3SR1BDP33AdQ/qVe0Nil6XDfj65r4BYEv3etqhor45XfL35EEL6W38uImHh
z+uGz1M1L49tsCBQxSxdmn6JsRj4IE/RpzddeLJ+hrAXY39pHp+CedtGkRQm
BO4g76ktudCtk58X4qPTsBwuPGdFLAD1Lf20NhBjEfmTmkP4rC/p0JqQnyWc
CZEHbo3E2Fo+ZiYUYmAWN8ccGtzeEG8H6mTmUO4I8bh/RxvNhPxcCpoQLdrw
eV5JBf92kcLtGxpfQrbrFDdcPsnZj2BR3ezYmgYYsSOqXUZ8PGJNPvJ1qMVa
4HN1lxusjSVU7gWKVrIE2YUVi7XHWJf2DntPUqoFKFzhSyLaRjHVt3YcePgK
w5EiWDv3ov+hKERnAgGEA8fdvdPpqW8bwVRlsAKOvw1rP5UlI0z8b2tuQV0s
cNXsRMQMKjg8SIZ8yBpSlGlgkJzCSNkU0zpSQucO9F6GGRdQ7jAurSyJ7lY2
hzdBQe5Dy/yVUbPPkyMfvRthzVDGSwhbJNlh98zu6ZHbb4oe+2GsP58kNiu9
6ATFTpDM+qbJhuYtLc6QeIkFqGaaQH5UTNDQYduGw4S6plv2zldGARhWWYTl
7NRx/x8xRF0W/RIKnZgJjYNRoTDC54N2uQEvsHDmbXiLkjF0hcIn/MoZ1UEz
GBGx5Dp9dJ4IujCKCgBrIj8R0bfOs9CYRsqGtY3ytk7sBqkv43j6QI6PkrPH
XdJPr2uSMvSRrZXlWb65XgBfFRKk8I5Oxd4N4F/PG2aHmZLBStvbJVFYQfXX
Dv2Tj99GnORgH3Oie/HL7MW5h1aDuEjqCsofeTlp1tdAxbTBU03E2fwLmT03
f9FlxiR2801k9FVkaqCjM7oH9mB4aKqDjrCp+ltFgNaldFAYO796/eU0CCFN
sgCC0KZ2xUc+IP6c6i+3lf7aTOWJPs3djpNMRigk7AjeCy6a7SdnDHnoyIA/
AfWdIXH7jNhH7y18C4Albi0SjD9WOVnSULa3n+hwKi4xnOr5EUGayTSY+M7U
7yv5CMQ8TNlnq+KK7bibxDWgRfECSusZWuAhctdaJbDu6zSjIMIKRuquCofI
9eXPEH8KrRPAhvo3CL4jQPsgQrRNAO83fU2ZEKGjpbRsrTAaQMVrQOndj/fh
OzY2fPjxh7uX34VPzhLFuWM+GbMjhsTv1e2dXhchxEMk3a393eDuPvtl13Dr
LZmRb6mr5HsyfaWricqCimilJyz8y0ZIS9vmXTOr6c3nUgb7rzN6l16ZL9a0
vE4bRXfnTXk9i16DK2M7NK+yDDB9ZvAnZTiCW8xKjhGsnZG0aF2RyxX33q0h
XMRyCG73LepyL6cx6KHPcnnwNsFv/4g8DrNiZ4Ht+6XTzkXFxK9noy3ruOWw
MYUZrDs8Rt8kMVW0IGOCkaHTCPQ9lI9gX4CxBYj9JilthoSML2vq7Q84GPtF
cG3qVaqGQzO7wR/q6tG5pKjJv9/MDg92VgzQEG2KBeIzUVwxXnHxk2wizm6j
HPrxuW3TAAXvuhjtEdHqpX3zoe3zxpWaPDEOZmXdI3mgJacJn9UyTW7Oslos
55HQCIiy8dcWCIXc53NZM5VP5e0brC4eMTEVr7QkZx1QmxooEFqc1BO2WB9R
VVmOUCrgyv48y3SFoOhqmQ2vC96lR4bRHNQ/ld51jQlBUKwfyXxLpZWkGh3I
i2M1J4l2geBZiY5VhafSVL8ae/ynFGQR+s26gUlr6qRz2bBbzEnnqRwp6FUA
wQJR/xnvSKSP6x794RNYzVCf2ShWYnA1c8PZrKB3AkyqIfyc+TJL/yBogzQR
Eu5hP1sNoz7sglfXZrnxf1BdgWFe0wK0O02mxypJdpkLqivZIWcDs+2GPm8S
cxn5REik5Im/jcGRno1Iue1EHQ4nEKOjn1264gs+G+sd3qLjtzTVu5/mH0iD
v/Rc9VUld1MEEQL1Efm/Af+cDdlwOkKhIPeD2Wx1zik5h0D7QDfmbt4YxEN+
7V8bmzEh5Kin2n7kUhwmpXoT3urXlZrY8HjzGYPQypoHNrpjF9VT+pHDPUAH
b2NOqZLZ3foTZw4dnDnuNVIdcGURCkTmO/6aeDHFRIGRq5Zj5lGg5tEWXSEq
s6sYg8npLX5zSnqt+w31GqZOqwQ0nJazyyEUC2j8oYM/rrMQ9ixzToopGZFX
Sh+5vEqmkm2ToD+F/HM8HLAyUxsPqaciM+bxakkFeUD+/cktKdinWYi6fSUk
0UUHqiL+YGrlIRdMq2hRRc6QUxJqO4RQCJgxWwrRH1mGIW4uXtOvxoLZ+Fdc
fJpHtrhFJ26lan+brpalS+OKg9AHgO6lsvbeH+DJa5OKs+Pe7cYrBiiBjHTq
tvzWZoSSyvIJe8pIKVxx9u8Q6pDkoB91c6M1HFgUgw81bKmR2EepqxItFzV3
52Hb/8MhmJaTcrdE30GQt3rsralPsZakzwUyap0h1eqBWQEoUxTgymRVkhD3
fq3TfzoAAgbx2MMclIOqfTZQdPbPrIDudxcXIjENw/2E5kGGVSP9i69Y3efA
ATBigOvqmjNC8JYDxYzbXyPuCft67fAH9m3a8ByLVX9pXGH78jrPt2abXvS7
l8P0yxCZNbzXuOT6CKPz47w3vdTviUQaMMLWAJUAf6/gEoDMq1b9jrQW8o+j
WTOHbBmW2+X0T2kvtvv0XyWU8PzMkvHy9Vvmgh0CA9zB3j52E2LOvs0Y5Na7
zWZjQOSxvRrncSDECHOs3SjS7c3KiuaqZXTOo/La+wYiv+//F00TDZuV0ogE
wgNoUhCCsBG1oBMinBGFdswFVJBxz7pbc0Kzsg6vjGsgd5pXdqNWsvXjyQ84
cHY90z/FTbta9QQK2O8aYGS6MNFPsK4Rw4y0eV2vl0657BV0XvKYwp30rAxM
jdz6XIwl3gewpD5VM6egVtg6PPBu/4hXT2K+psJZJC6jKwJ0Ubq/qSvzGS+6
5J1FR5/U+kkqV2ii7rZoreBnqmh1Q4/8ogIoErzSFw5Zi4h2dxFQBP3UOrJR
0mPETCO7dmfrC5HH+R91j6eOzFnfqH6nXoWahFMCq4azr0IB1oC7kJZtD5lA
EJq2n6yP5dk/dbVrO0jhvMxkyp+ZJIHltREqBxUnBS2UZz9lAexOQTKr14nB
4MsTDW4/7Y+c2wbqfj55f9qnLPohrqMUw/hZ+938fanFmbQvU5yNA8NEW61H
jcaAyAVrPmR+WTjRIo2QwXWHMiuumXCdWOFsElaSJBk/y1CbJRaNrWJgcD9j
mD8J/mAfm+p6UskNNRxniTuTRXwtJS0rpZOcSJdQxQ5qkF4KhVBmtZI1HLgO
t5RzbEmmDye4KaiHEYnbuL384alK+zSxzlGifzyejozPNdXTT+1Y0QDEtnzI
uZEGA+o9oPMzg76YDjjN/Olqh9VLRhUhWwfyARuy3GDThFN6ic0EuVsm5F/R
s2k0Xx3lEcLGp2y3bRW4hB2q9abMrUinFfV2d39YTtYG2tlTkYOsfgTC3GX8
veQt6nFtSaXc0dKflhb/gbjSib9O3NTa5cqn6Ugu3wztVpZ+Xym6SPJbQsV+
ZzRu6FKhRWdS3QXiASzeCQU0Rrycd/AXrYQObC6wSTMgkE14UGE9UbH62YND
cCEd+ULwYF6cK9Hxra72eVRxe00U978qOI5ggkhBQWFBJNNHsSg41AL+jm9W
z1KcXg59ig0amPSz83NAvzWSIwVEGKhqo2e1YrWqxwVl2diiyHBQw1M2jhTi
3u+g5pb9miX/XexRf9XHWWJAUQkOFg7dtCfB915evZ/gZGi2wTwaS3h8ozvU
4s7FJE50+OEo8nLXqLFe325KA/uXmrjpMvOQW29oXcUcTjil7LfgNU0S38yl
tE/Z4B9DJ3rf+108Pusit8K17FspMncGcbjASR3gVkmqI8V1boTUZIiLlKNR
XUwTzhQbcU8IwxDBzFxZrp4DyFY9dvO+bRy9clZaLEAxXMhN/y5dGCPT2ldY
uIeciY8BthES8k9HMmWMTo0Nr35T2eha6d9jbHzL0fbQXUT27coAgxh1a4hC
yRtAlwBysUP57/LSCiD1wENoxThyqWw5fUUMWndJhNhpM2B0SR/uZqYHB70j
qs5Mcai94UdQeZOm2jcdeYBucZlin7Y00u02YYyQDSPEyPRoodIDG6OCcqP8
AqV/GDMziMBFJVYR8NlY8CEZX3n6VbXvLv2zjujaxAL+eyKh4I50F2yDkjap
DPS136xU2yRFWLwYw5WjFgDN152OVxpAaqWjbNEKremFgm59tt21QTvfQy+C
xoZz5y0EXbBUgggNdKuag0rh/IwaymKmxXj6/3uL85X5GKj/ByL56pcIiUra
gTWtCua+toGXgccbcZ8ysXoN5WoM3KQjo+kLXwrXUupDM53r6TYrwn1VFBrM
P3TkOctqlJD1P8GyvjXpYn2VZfyFnZ/tEKdjErPPptShZ5Z+IRgc0m00ELVq
ifX5YFLE5TuEqbPJnxwbhLj6Lerd2MHqqRO3euz+TQ0pNHKgPBuWmg1SaScc
r+wq20eccpuvoKJsO/edGmv4gNSMfxoE7wrIZRatKfjlRXQYdIQGFHlvSIR2
cwzFjGb4Kb6RnC5yLOcHCdC5AFWD89DfWkg6meGy12VUPC5t+neomqwXLSKb
eOKzTIhOW2r1aY1xU5gXIOKXLnk+qSFPSVGIxnT3cuVu7bp0fLIz9+1WdIRT
4vgjT+g7kzchrx2IxqlnqJ9vQkD6zoUEDZiducT+MYLmlho9Fgj0N4y5JhTw
JjP652xa8rYMc6m1/o23ozGWigGNAF9dYzWCZW/znm6Fx+YuNtjiAhNlqNx3
xXTjY5kf8eOKYIVAfs5RZguGOukwqE1DcQkS1GpPQjCNYCdNC2xgv+xUL4SA
kF3rwq5k5+k8G6oWIKimjQFk6R5l3Eu5fcbsSpghd96dhj29CSgLlaWOGY3u
XOEnwCA6t+z5bq3eTYmFtZC4pVxRZq4BJP2bABj7gy5cbNYSC+Cj9c2c+D6w
6suJgLJgOQOO9J74BfNY+s8fh5FZ5CXcCF9UT7V8S7Z4/EJbj7B9l7MVatcE
eFTDWm2C1cyVvNbz84CaFHPttoJdR4OyRjIc/ZgT4987wICH5gICUaxzgICI
/2kWF4PvZIRjkD9VbsYM3lJJIY6zMrk4oYMDyGqwdtDgeVZ1Skd0a9UDyXE0
Esb4eNwlUv+ma0Bsx137fQnJhdyWhRbSAiP1gWmVZNkmy6q4RDRquKOf4xjL
ZVgjWBCPktbUBFKg7SN1W/jFZEBlFAcbgqXihmzc3Gw7Z9DjQwDl5HPduVUS
5qbz6RNnWtZI4LeT0aIBDkT61y21MJZ3ZHAFk+ee93c/OF8y3jBFFytgBWLD
CedpB8yEX9nG1+f1bovXZog33/JRWQtfBouV+9JWnsXnqj2VVVPeu4K8YG8s
MFwBTj8G+0fvDJjqrudLBFp5qkbibEuWQEXqPEHKROAHMzHW74zq13YmnG6z
VAVevNE20PWSjjbXj3vdoyX+kpcRn57huIHbiTw3noNFqu8PBfjcB6ABH6OU
EIsfe5mJWFIlQzDsQJhuUT3XL6INshf8wMT5mOa2ZECzNAzHeg+d9IJyHW7K
uAcypnFcFBfF5gV8y1J6fiEJTpfdymJxMr0gYlvMLSJof3XZCBYmed2IwSNl
azO7r1qjQEgH6AAIp5SOtXHNNrOylsti0S9A4Ovkbn6h+/aBc+vCFrqLWh8E
Cw/d4kv4hYJn+1hHJWQq9sA/XggVmODSL9Kv651d/NJ31Vz7Qc8/aAKQAYA2
x3cvLQ/HUkWfM8k4OvJ+1HjhVQwyPvLCYTaHGNxjh02MnQfQXE6DSA6P3Fsl
Gn1hCi5yvRezbImhrs1cVlFVqWlbqq9MBrTjYFPX1Od4rl4OObYZNuEsy3bi
rhLRe4L7ECHC7ALy/ZIAFs2RvGykq1SidlGHk328QLcvocNbiuBOsnLMVVBR
TIALqCn8Tq1RO3J81ZAtTXAvIYNpiSYJ9HRB2Hm46Uwch13Thw//IbNoI64i
0tDtB11Lf5/KaWIZhqw+oHEYHB5dLu4FfAzW6AQizT90vc2pZt8gXK/QXivo
sKl6pRoLwoTohdXsz4lTw3SScdIZBj6G/LvG9RP2i4U5xh/DNfcTPgHbcEkH
8VXbSYtI7lC6HKlICak5t+AG3+UrlnzzlekaqTpEnOoJJsogA8SCr7U+qZea
LaI0wBaLhSyg05N1c8ZxesDTletnHpuzeIYS2r1OGv2NqfQkwawU/Wy2V/7+
Dcwb16XKnRfvB+MyKIfH1sjgwgpwTGVasu3EofG+4ZhKRwyR6QkFepKaBUgP
zFl2I5g0Fgl1RYY9H8LaFjYRifv/vBXBA7oZ5v3e/BQR4lE4vepwH68gdBDy
iaRLHqwUfLEg8QFaHe3VmoN1KgE1+CkXmS5flZrooH7iVqwPFeFIBu1oKHH+
jmioElwOuEUutCDijsHDp3F1UE5kLNPg9ymuMqMH6Kxc/3GEpg6uTH4wgubF
xmgh4xAUH/jLUGeYSCxKvo7yKQNsRo3jCkRnBISDey1VKVdJB2fd3t6R2JyB
b647cDxdubCOIjJkgqftyBIa31rQs5mzQsVXYsczhNaKRgDvYbZVQweb8HjB
uGEf/40TJBUYQZGDDnRabARnzjucz38NbGg8Sj2mXijTc6EnSxR3emEh4rUg
7ihj0vvtzDVn4N9Wl84N943UX3qXaIhtiEle1ZYaFPNawAwuK/fQU083OdCK
nKKQ0PXDm6T8e58UbPDFYP1RTf2q7C4S1hpHVslJjQRzqn4KPlwx61trZ+37
P9Zz1dOT8/o+6UlVL4r2ycBnwBipjkEfFMvTnsAXrzEP/saysbEBLAl/pF82
i/Tp93iYvvnNLTbFXUSUfKKWncJ1mo2NIe6Ext1RNzc5TogO4YWpzvrE5V83
eNSyN8ZKBpDXR+gzQB3A5yu2B9MlCEbGgNYwYEbECqZnuM9ZNSg5Z7xUe9t4
R4CpY4iw/YEeCkzLXyZcSkKB89+7/DPOnE6XSZiDZmUYnn6OQof5NFV+BevJ
U/RJEAcgCNeqBQoS0e+7ki6yU7S6I7JCmswqGyE5QnxzoRqrunNs+/C151nT
ar+1ooZN2E7eHUIwegpx49TKsnhR0BiW4WhUsh26f5aHDeL0msBE5ZksM9yL
9/8ep58i0GTEWohNtEnCYgTsj2ubRg5OalyadrguHP0iCTLuuck70Nql+fn4
/omj3xUp80ji9IPFEMw2O5/bqduFdHl2lZN/riE0OlTyL3DVx+my4uI7EUGq
vUNrsr9EsRZi/6DVaUHpKKkOWJCrT6WMZUioqZRt6SWpLCPM9MPrbQ0h7aes
SmkODLFSd15gXjvIYtW71Tg8CdX8wbFOmfTTJptf7eXmmIPdFyZYbe3S272/
sC8uFy1L4lyKIC47Ugnyj6U5K4TsUWPxUaR/OphXwMAWGPkro7UJAW0oFCFo
SDZEBpXnBxVFQ+UpGUzttbkCHP5yQQqAZXRUxGS03AM5qUVpXrg06Hd2qLRV
uUPNQYOSvb56uCpS85/8VSc81x6mvCz2EUIeZr/Sc5hky03xMoigso1fsFbO
SmWEWl8SI+tNXdEldwh02aEFGYZkMyU8gawDNfGikwqjg8RdvV9JuHw5akOk
+DsRCS+EvToEb2EvDyey1MxhsvoiJbfH9Ojr8bGwMzAMxA51MpbD033ZZjeC
rM6RpTVkORszpEax781egWtvz2iTT7UU9O4ikH5nZTgAfD8D+L6+5ZiBLxSg
Ro7h7YPYmqMAqq/aFARLqeieOT9blEJ38BH85WgCyZ4KJIiwhzNTGV+iEB4N
tlBSY6bNN3g/5osBQrikOp5TUgwzVIi4jRVlUO8pUoetFJJCR4NIATGYP90v
BZc/hzG6YaKsi4NzxA90gnG4f81s6OAAODZzulyHXGQbKh7OOGPX3QdxXxwW
g7wuWdDkaj54SMH90RRcxjJW8frq2oe84VYW3Z6eLniuGkUOIUx0HxSzsfyr
XrEx/dzqFNk97ddQlK2mzKrrah2qos1qjgjEUH2k4EXbjvBMvWN2MFfdWaF9
M7YlU+m9YeVyDKd9cs/wnferY0qHlRe6ETXldMDwvi+B8LATQMkujv2szmZ4
Koeuuf6N6/7SDFoJwmZ5zYESy/ogXCukUXAvn+liAfwIvLBstMLCZdfsu8Na
6/bmdh3glvuwG60I2scnaI3fVFjKqWn7N5nYTMT52QcLFb1Sx58gzpkgcEop
2aR7Xiqc73pOkVGWRf68/0yvC6n2n0i6G7HdlnTkpwWPQ1jSVm6LFhfB95Jl
kZG0adyM5cyVwb6+RS3QBrTSIfqc2frPi3NlSO/kn+8dDcy9JnKnj0P587tT
Rl1SV5BFqX5RqRrCLxvmRB6Hu0cNv18JZfEJNPb2zWN7D428R/tmWFNakY4Q
bH2KvkSuA38LAxEJuNUUOJYzR3xke+oIk+jYVi/V5fqgqegXsNB51QCdKBJK
ZpOf+AUINpnbDoIB8kc9tumZEkltFwKhE2GmZrFu9GtV8UbDgWyZ1soxp0kC
bUNaz4y95J+M/GrvMRnpMhYwmnReY/gFA1KLGguwcAsWLF880oW7pJmTcoPv
EQv2JvrLVMtzPEPjOJgeowCVIJQW1pz6jczX7OwjEVPLba62qS5CjG9v8lE1
FXxciAJntRWoPdktU1xEVtuwFjAwuqhQwgL85GyddXIOc4lE3QvrZDxgBO+O
KrMjSnWgthbLAX3gVj/dR+lcML7OwGNehAT9Je+33X4GGp4glhPzw/jnK6Lw
fuf4xLTApNkt6SkNitW8TjVezz4I5surjoHQ7Ti0dktgooq36R3nqpyFrwVL
4q5GtoVzCtH3u5oGWYpaTMO3YLMY1Ic7OeTEGwExk7nz5RZ1z/IXgJNsCoI8
BvrIUf2K37XaJosqspghIFabVMFYlBnFSTOyXKrIhlyVapAVOFaD0QNjz9ds
oq8TJvE+GAwHFxI78vBvx0QLsWDtz6YPJ99bhDT8DVbpW30ivGRfoXsNUmKa
bTlOLJe+mbA3Wg+fObamMsOH7j5xWmUWew4JEOHEkKqsHCitBV9mCuNoR2Y7
V7jaYpwwy/kZkcUn0CZISHwayIak15cDrGzC0c/dP7wAeXETy2sEF+HXGatw
iB5R0zeeL6M9ruIIP2n6Mwq3ixge289rE2Z+NLhM30hgDfuBZypMz1Q3CUNf
I8m4zM8mMrWZtPTcPkKs3979RgtFORHbuvzX9+k2wmIKmdpXT3SLI6N4A82e
SslBWwRC5B6kLxpWxLT5ikL53CQNaEUV/44HxjOYrGlvV1fy0QMMguIlksve
MHSzHKMgrpvMocbDtHOve+jrVlfWKjuqzDh8B9P4U8WHy61SKQpqVeSLNK88
vSFKlcACNppBdLBcJHMqVXzF6t+ra+oRl/ndCMme1m8ySbqD4c32gzUgdPM1
ulLYIy15eiIPKWfTFqteEcJHliXB3TxzyYEpeVUBOUuNmrAzuyWm20iKajaS
7VsU4s3F32HevtkcsbbLlcjXz/082QuphfIwA1CHiOBKOHY5c95RCbCN+xUZ
MXrf1RUgwN98vq0mA8VCGcNpNRjXNcAk8ij7xE4TCPP5I4wm8/eB6jJHnTHw
Pp3AosLK65nKw5MIlituGe8pA9Cf/3jqRiB7fykeQKW6kB3dfZerGeyDIYM0
6jGG7YiZ/yNrXXKKMLO4a4ecL98jg7efC+8F0iSr6IWvIi/PGjoqrWHw0QYe
YpBSMM/iSc/00LwOrUDXIM3UEwBrImQuZPlRwRd7mwD17/tfN/nbqRwrjw8F
mn04jlOGXVHxL9oExvkw80UmOTdKwTR0n/yAtAQVI8awQ15uI9vN8tHevsJy
TRVf5Z/WzoLQ76zvX+eeB0fvXg+YCN6jPMNDaLF9b9LGxvJT6xp4WX/axn/l
89c5RVtk+INw0gnnzHHB91eigfzAfMppnsRs9Nqn9uSkCF7aNn+nANwiUyjt
6i3+noppOzIAeIPqEw4+9WTY88qIMUlGZ3RbryVcgo/bE5ZWi2QpHopJvL9C
ccE+OnhnDMPMYxak6OrELCIlVueKH2ZVQV52jrTtsEbqAs0wOiqf38PfyKh2
ujAV3p7kU0iFQMpFju66yE5ZqdCX59xO8/TMdzqGzkEYwzf8nxgMIsShwwMz
F2TTsmuXbHBWTeSIzScBMQip7g2clvyMJGqiJFIWVclbayOIQXhBqBwlnX7w
n+tg8qO4WhFPpYpV/BZASuzwu1yTVSXHdfXC8+WKjso+vFsFJSGi7FlDXyuO
eGDWDfA+1/dJZvHNUzDRCnoYRpQpZrFqrQXP6Z0Fx7vdjPMu+3e3ZjPm0uUr
KAb+m46TAnjdqDZqv7pSRFHGGL3zHLJbD0V8quG6rNwAWlE2cHS/VfTowmKV
rs/Y8tmN4+kTS+7aesy26YESjat2rU0CbJEi+59ywAUpKAEGy2HWSGpmUKa2
ZOzn7eNfuimhhxSD5O7TFYqZRTGmd4amRluYBhVc5J7P6ECfjLU7D1LZ93FC
ihLM3oNQIObjIPP1jEe8/W5AI6kYaxrc7UWOqj/WeXNtpS1CguJaImYvkqml
scDw2ysS2JT9W58tIp0Jg9ZjgZ/3/nvuyRFbi0/7O4tUu35HuuL5aaVdHAEQ
q0oZDB2/Q5Zblo8ojntiDtfwdy2T8Qg0VkgKkgOOop3ljR7wTWHJh8Lmfh5C
B1QpCMEE8FRvdL1vohqBYYvpHIINDyRg325kdOD4ojSq228fbYnfaUbUIhB3
NG9UadTPZHYwrSQPd6TG6O0cBzAjyM9db2po2toDcwXooVHXRRDkwpHps09f
UxOeaqdEgX3GEC/i+MKvsiUE2KxtET3Yjqekw2iwvTkBOL1rXHNHem/KK9Oj
WA7r9m160jpfiCyybJD06qIqLvzT6pS8sIBwAz/89eIZr+q4b6UYr8eWn0FI
lPvGgb+ggeMSHu6rkJSfu6ftoLjDcOrI46ts14p2nGNZ1V/oBm2cxLM9r1pW
ZLrV//nyBkMBW0mYcfmaqYzvPTqShZ38YL9C+NvRM3bYPBpOntRIGjnnKEpy
Fg+3K508hJie+La24PLIdukY7rqSkFsZcrgq+iWwX+m1R1Pl5XPiknvpo8w5
+88IGEc2QkOAqcw8BXGxabT1K6oz1fxQQAQkkdjeEwZh+zjLciOYf5rEcRQ1
ayxpZUP9QuaMTvMqRxqylB7D39itA0gl6D6XmNbCH03UYZiDG4SnZHfwzNE+
Insz0OC5qupSrcGthIKuWEq6CSVKZtnlBNOpdbEoZGfkFmJqrUcyfhivApPd
mKx3vRHx6oWcVHpiLtMfT/SQu3pYdNCO6YNtTTReiTYURiXPebbHkGqei5IZ
SB+lHY/wMcLojBZ73rlkhk7+5LEWhyHCoVYSxRnB7TZHTwEkH20JGIwvnPVr
LZPUczyaDhpFyoSPzZxXXTPj45o0ZZEXqjj53Dpp+1/117voZhOCLsSQiJmr
2o4/xOpnLAGgDMK6mfxJYLpvYJo4f4P1YNLVxmI25PetT0mbNotAmeGN9bD1
HkfO/mEa7hXD3iYod60kiGl6/+NwgA+Ng3u5Zui/h8yoqd8tD+pRTTinW1Ha
8loO+pwKdK1KEj2x5efYIz7nQBzl05XZju8RnnOnHfdND/2PJc9xqGCdhplA
/KIJPWIdqLPcg/KW9YSYjUNLxZtQHFD50yAWE79+VgtE/We36NEz1gi7bs5v
OygrGIeoF5Widig7yDPZQ6CoxoWtQLaUR3BWOm33q3rXcEJ2UrlR42MPVJZU
kZVEhvYHGzSVhJuitb2d8+aYN98jmCWQQ4wGgoReXS4YlQwZUFgcDrjW8Nqg
RdHUCJ8wIrbICf1rTIp3u1jDzX7+EXBBubHtW2Ru4M50euCMPQaTUA36pZ7n
icgyMDzOAyCwQmEG7RwKMNLSdEkCREwpKeH2LeqHR5nztiMW3ExMn1CI4PgT
FE6T11R0s7gm+euLh5pU+ohS69RkTi+XTl58g1jlGiEumHQYc8RQbVX3uBb3
WgWeREAs9lkIeJmWtDXbGnpjg5qDX54XJ9m8o/24x6kIzfsEpNqj9cbF5fgp
oHwAPjbZ1ZgtEfP0lqusjW9z4wGkvL3Z1VMDmgJ6vvQjE6hsb3hiBkHuC9VE
MhoMWEiH9jHPkgD3lGY6ucFoZey9NtU5KtYz+IHF33bJYesae03mwF+QWnIq
8bDEVYD+Cm29vY2s1qdHPMlrRPkIHSvQkzsF4NqNHg5vLnJBcYab6UdH3BwT
QhWmNwJskZ451rcco/xO9ZDCsF93/nZrBVKGzL4aojGgYasI6xO4eX9G3BlM
fkQSBnR/MXFdKzSygrQ2vvM36Umx4gXdeJIqw2H1hs4dFzmLydLVxZGNvjod
QFWrulcb51hzV0cWkc1olexwa4HhCkMm2iGHt0W5oy/uh5wit7aD3k9sOmhG
7Xvo+iuec8SB+M7pZFlDE6GRQutt6JuPayU2sIczKFIE8jTGLrzyLRrJUFzY
yZARnoDbi3G9b+WY+Biyeq1IQldP6OdO/E7XeSyZQVSA4PgN8SWuEe1rkYT3
KTWRNRA/+1LxWNBjbeP2HXOSnlHfZBEBREJXOJzVZF660WrjG7UuruJ9B8ok
6DmFK33mII7ecx7vEvWKOc3XpJpMCp2TIb+OvCv+q959CAB+GCXs6dWeUEPr
cl3UkcxhZIW+t4XpWQwhOvh7GZivKj//N56bTDvVSBAa6IpxZkzaR5erDUYG
O6nb4rxjwnQXiwRYMyabUqGWT7fYDXqetoA+RPNjrCyR3xenKgna0fxoNDr0
5v/YD3/23mEOMi6etONcRy4NdiVXT3P3sazSvM3ZtLHV8KrJ4kHWXzFBVus3
akcs2xJRHJuhpA9lMMv030XUQrmC7GSGkttdIQfMMX/QHkOBVyTaZu8O4HkJ
C26iFTvzJnenb1btsUYkR6toQv2qWbV84iXaaH+vTrLWNJp5w8reWTHhUTQr
7aWMzobGfLwwm5rMQxYuqYQIts+uL84mYlfjsKB6GIeHsXdB5leOJpbkpxtV
MC1WjRqmcskPw/H+LaVRXuCm3SwugYmuHabvazQOJrcUfJ1V0lJZ/iN8uqBz
Xt3ZffVUG6HD3sTpfTLew0/9vzi7UtfOWSASndu7Ccsmhu5IXDMHBEXr0tv/
mdsi9H48AY1NtrNswWJ05r6nzBg5FdRgBQW74x+Raq7rJDNgrraVV5EztFCn
lAhizK2VbzDO7z4gIrZEqxkIUvgtFiSXZQY+O9W1vfYU8XsOroG8dHlmE1tk
0kc9Ht3SVNlDppP1Jri6wucCtIzYuNM6SjWLGu1kia9J8xNm7cRrCSAY911f
wQLW1Hr0vYnZYZu4+CGIGel/foyCFDWpLehZGYjwZh9f1lMo7KmJFFR6E7Jg
lwhgZhOwZOp1A5yECrx4GZrtCTdlwRbmQdBLUkFQc/j0jTSZbVZxz/IPX3wX
n+6gZbuzDYoQY9czO/hAGANnt5y3xeARqsKikw1g4Z5FPtvoyAH22HdJHhbG
sLQm79sN2sl8RQamaEQBLvPYCIS1pSuFLs0DIbSze9Faph7CEdM3CuLZQmfh
OuXWDVAJMkWXJYplMHBzrgkBaT3CJr1CMRlvGeRKNfR5CIxWxMr9x2c8qGSK
c5+8tMZpFYEoGAEUcRpzkjsXlWeJ0/DKdOwQsDua4UriL2giixAZxU9FnZLJ
phxvaLIs3FaBy7vBKHqE40uSEy+b8Z6eg7cebPPiT4OfD+vLiODuu0dunnPl
B2x8IHhltEvzmedt+mgzlu9PtNvV5SmDrRvEIFUOklGchwYpFr6b3RF1wQek
UJOCFzoDOAMm7qxJIJHUjunU5NTvIx9JAd1A5zXYQt1tJo8McRynqygTryku
skehlDKMwVmBHKSDQE2OioxyGzGRAVeNjpPjl20sYIn4WhfMoHFIs77GyYLv
6LRJzrvyx8YVTUkAKkq7TTO0OaXPNZZStfDqxI0gKTgIugKfy1/P+QoVTR3Q
mKJ1NOg1G0m6TdbbwEUejcghu0MDj5EC3/Lgg4Vkrw/KsFHjcwSt7EubsPXY
sTQA/DVgfbr7SMAR/O6zwb4qITAu+G7ghmSwBgSGhxChVM1pYs7bkl1BV5Pr
cWe1yTKO7v8esZnTP05we32pBGJ27m6m1sBizbHKgs2ogFQHKwMIriJBj/g9
3QlgfWTh7sHEiCS2el8sNh9yqS9xwIcSYuajET6vsLr8Ik5MWqsxBKJK6QAb
/El/jXxo6zjhu1l6NHDvYCZFTsxraAaIuO/OF2ZBvFzZeAEYI3L24c8WoJ+n
9auQPjXrzfU6sQ/3uVjqktH3BmJQIvz5q8rMp+8ot3UAMICPOE93E/OdiQnf
ogMEJNzYeBRufOkr/bTAN/kheGLJWfeNn2ZKMjtWqr0iYPlh90Yibt5/4Pne
2WBfATTB5m5wNwOTvHfDkogwWlqj4knDYwBk+Fhqqc58poaONRMqsEdKjeFi
2z6LzG0uTowcOdLGj8OGijs7yqDqDoaIl351xFzwJW0t6s0htVZet+Z7j3BB
bQdgpwlzxSDpvLp+TQpnPeqMym9YnA3haBLtP/VRXetI0b/XyfhhUUhiK6y/
jhlT0JeqSyWtTlakdmSGNvVNj1nPVtNXE7KmwEgt7TCoIK7mRF7b41gi6Fwf
wBVbt+J6jGf5RpaCGYKVI+lCh0gYxYU1Kd1V54Y3yN6M/spQ7uENDxkw1RCl
SHHE8NHxfwahRJ99CoQkdJJVZ3zLk5IuTQ14BIEQVshynzxJdcfabl9UR59e
Y54ecO/EsprfdhHpK4/1jz2E+hXp8o2ug7RH0riDZRDgaRRSGOMuZeCeJi6K
rWZ5snxjMPRu2ujvMeFHa2p6Ep0YUin/RaR4dPfp5KD7TJS8vOttvgmQSN4s
4t0Vi1lKXTkTgHK19yAR3dtUrxF8cobmx2WWuY+f02U7ZCuqZeXngH6i+ZO+
2XdJhck92rZY+zTbOkIk2Qd96MGXeezFsJw/cyxztBTHscjJAcHZpkFMYzFf
yzWRBahC9+JddN6xqYm7F4D76H35yuL01NO8u3gXG66s4ET9ciIMDNWF71Qu
HSzcQwctDxbiuiBNMZ5vNkLXWVGNq0hNYv33+9OghP0p+s6qGBY1951kXi4H
IjND44yzI+XJZ8RcAvulQqlrjO0zLniIolRSfW8xssBGKcvZ2vEXg+yEdTD4
ImboWfhQFCfVSN8ZQ3jM6BvPtnMQ4D2a3MEaTA9Didd/fkUJV+HixXy/AyJn
7bzC/U4qz02hDktIVhlOpwz/xcIoHMzdSTOKBPKirclNPd6Jp3vEZItz1/Uz
U5oGw9ZZOUXhiVALcKYPrHTyRJKfUGqFaz3Jbjy4ysoarLFdmY5kkZR650Bx
irN75zoVXBCvdH+PM1r5VgDEii6fNipUHLueTJCtLbfkHy7qZ03S5KIyHgYF
Wy/zezfkEGz2k3rkD3mU+EDWQlydAt8LzljRONqqVP4SelcB/dJ72u0Q95KD
K5ewQ7MOpoancKuyBVRfvynAaJX217mic+t9xDLgy/jV/jnbbKDvozQSNxQE
jI+j0thDw5FDQV0zYI3K3ebTNPHtrcQrLDmC7m5yUkfTK4+GG+v/3YzAf0eM
GHdlD2wuOdF4qMzu2aMonUwkCwa3AKXzitwTfHsehZuG2T27BVDOUV1+RGWR
2m0jab4pFrpHC5w9Bi21YPRDUTZfOovfvgwSvxhSHFZAIShSFHcSwITwiqro
212iNoqOkJq3lPKVWdSDCqd3zWeulKncVOr1d6U3E6m4kSYHbjVJ836SPYPa
84h8skLbGS6PsOLNxT3QNoEkLg4EiPvl3EnxVU/hHheGtx/mlluniZ6UAKJ4
8YsQSblm6yxJB4i7QrQQJGQ0/xu0/gC03V7SJxPFqwXmgPU6zLn5sPBBJbVT
qoYzdVg7h9sBb0snw5UqH7GrFbdK6NM0OwqqpZk/cOtHWfiQOsMyxV34w4yc
hxgIuNvFoQTxAAogWBKhEBKH5TkN+J0efZXRVYkuPskk8bH48GX77T3YV6o9
WguEjSEoX7e1kRGFes4Hg2xKO3rFWxYchRSRASeCciCDNz4q1r7RBcgXtXyE
2mYRu8FIRw+UpKJJGPbcXIpqOVhetNTvS9uHkI/FtDAB4/C88KkXxtDvl905
bb73ImJwLH2lBIheQEZ4HVcoPhDZFlfN7RdyWpoxcsLnURNhnMEWxOYm3rdD
Z/foK4/ZJ8JbINgvo+Saj0PJk+cuBSjbXkAEEEAQGcLGHV63v9rXwIAc5ZXZ
y831ugQ3UMUS1SAAVgoqxfdlNI7ApeDzU4xpzGJzhJNem2MYSKX3L8Vh0ZXG
6jhFilY75XpYkou4UHUmfLpT6U8m7AWUeJUsD+iHn+UiT5i8dKhr/Iy7r8PY
Hb+rhi3uXHG9TMGrlIiM0QP8MMJQnRPBUSLSkOv9nhVI+XZ5cNiIS0a3WG78
aMnOsFapWu0TpGZf5+SaH8neDWY6nsNPA/nfBbCzZLK4h2bBFHFETl1DBsIf
VeIQtIn1agkQnIwMNkEFuJo7c/lW1YYVRspiyj1yAf/O31XF81jG3e5CEv0/
OvwzlGCn0YdnyLAUlJ7zpLZ0TNrNJfspp9ttLf+yZWJIK87AMQdUAzAanXQl
3DkJeUOjQAwTGkBHqMC/iWOVrPxQHnie3szZCFmlLX6OqTwGwTQR+DUuBNIS
tsAurgojo0rb0ecxdOp+/fp8pQFSZclUUk7hmrz85nxnbU81g5IoIXLfrW3P
HSIGIBwdn000OrjgC4GfUp53+OTOVpbvxft5Les3CcopT9hi1TolVqO4h35L
zWCpki8TKcN/UQYMwt04H6hcJw+WdwayFu8voHDv3dUgL9bTFMo/wJS+t8rt
fsuH4UWce8JLa0b1+WHMiSsR8DngEz5o7lUYID6r90pzzIqi1HcbjgwRr/MO
Scdn8LDHtPBo2VJbFZ9q/vPexsw36dhRBJbDsF/HexOpdh1iE9S4Bx+jdvqI
gXoibYoj81IxvEc+eiPHhv6a+s1Hu6Znq9KChi/IlW57AQmLe8m7/eedKy7A
w9pmlJUokkUesR8BbSyj0hAMQARwGLGUIau00pRNzy+Ph78idWhjX+wUixOu
QivmBdCo64TxFwy5t6wNgrQZ71TizMsvOlpN6GonugJ/asgyCBiHzfQ547sW
hjQaTBtdOUj+zg3/v8T4WZZTy3rm++pdSMw5P04Rpp9+x0U9jLnbfuDg1lwg
xKXxgeAbkZ1nDVPd2FtSc8c3L4oX2SOLVW2ZdwSBMb3BBtb8uKNtmyomfeLp
XH/xPB1GERdEc4IM/m6RVeXpPWv+eeUoGoThF34MJemWuILbnyBKbYb/97sw
Y4LZRDE3Y+NrCkd2/Vjv7Bqn7xDaK1GrTrAlVqGPLKbEWrlm8N2WN7p5ez44
9U1QxX9CRDoKMYuTgQ5ZhRKFrVYnR/eaZP5VvTaP+tlXoR46VwMVOGn6DLQn
pgSS8SyCZw5isA3NiknBsRFfCsVaPny59z0K+fZMgWgT3rKyei7Hlws2xpog
KHAunO8sdauoGrSwjkPrvAvl3RqJteR5fTCnZ6iGaG9vZg+6QMa7HOPq4H27
1Poda5uOF46NKDc3yG7dX0rPoPW88/sjPKuHtvgR+/m25eJnsE6Y9IQ08yVJ
lyl775Ojt/A9mcH0W0qUnNSTNoomW77Y7lL+pNt2y1rcKTAbNrNWzVlqB25R
os+hbe/1Wq2M2sz/vCDID8lXKAc29p5lPNcBVgz4qhzsCHEnfXx9H3GpI0VE
swBpl7V9rCjBV4noGlw+LpZ1cOkTCYIAnia23g2fwHvGtu60UJucXqmiBDkJ
xx+ouazsldEWPWNzAGw/TuOhQyOfTJW1xWlIHdxbevJm9rtGPVBfWuC/S0xt
oqekBwOuzv+FIYRb5WBsCeIlZxQdELh3DhrLn0dxgJnnTikoHxj3BC7sbtA/
NAG0whllVh6a0odIiUdZTViHn0XBnhtdMbH1RmUJ0XkMeXqoFcQZBIH6L7cf
FPNKFEBJb06Z3ih47gLmNezzDQLKtwq1+59583ldQFLOILEtO3ZgNMzD3ZlU
8KTiQ9F6XKYsV1VShCu8tg9DYu6Jjbj/Hyov2jbzCVLzYTRc0oz39qIpIisq
Qa0p+Bmyr1CMP0wpoUe3yNPyFsyX7c8YiaGv+7kcdbqQCkEeFPCn87NZOJk4
yyqhml1bGYghHv2n+IggIiSwP4yckoEghi7E6fsCgkAZ7BruTkaFjIWJuZam
w5MzvmGetHxgtflKMnR5zSIAOXqXS8bw0pecepDvIoO7O/oCUCJYWAc0nncn
HatrNy5d/g2uwXl5HmubsjMBY9NF3AFFLKo7K9YeXixs6hRJEJ5aFd/VzR6o
Z6qUbcWB5wOkr5RC0uGH3np82CJUb8oEFZWPbo9O6steQ9ZyYW1TAOOG6uSd
k0xZrzLiPI1ewpd3jACdfwDstesRdJ4mwPHnUS64a4NopxR4V8mItqC/y942
hbs71n0ykZ3UGp+Rvu5G/VcW0Nvi98ggkvSRnB/dxRCI9+oL0/vDUhzL29Nf
gvYmUddzyB74rsLbpH3TiWSmFOTM4cb3IQJQSNkFwhdgd84gWhohw9rK+A+v
bJEJy/KOoOa1mIbs7L7ckrE4ukVFpdL0DfE817l6SrDAyEM7beTauZf1n7vq
RTKuiwi8rsAqJYFfOHYY58Dulam3abgCLJ/BZW1PghLx/aGJLnHPd36Y43Ze
vms/Mj/rzrcXM7jNDvH9mIl7ZZOTR8FnCvV2UEE/zcbXUaSNdLTOKYKNSzOA
l0MHg1lA2JsGM7ijXTXn6ZjGB/nIYWy9gsRsbbICyNyV+cZqH0Jmx14WEUv2
R9LcMtKhgfX4mcWPXa7QbO44pMdB54xN0Yqoo6+sYVMrD0O9meUZ+GU/ThP8
CD7ePfJxDkyiWW0fO3qLAFwKwzaHPcclEKVEhMNs/UOJU1RrAZqe3pcZi1E9
dgRYSd8frXgqIKAvfxY+ZNB4vFlI0G2KdqrFH7XBGdHxb/DZ3BtJ7zXVmtHp
q/KmZAlwif5FinvgD+oUadMYBHaZ+9ibzuwzxq0qlnLL3kTTTnWu7riJIuIO
AUO/P5txMfrWeYOxUC2M9uqZyfoDz8q21Q0oQ8FdaBlfypmG2GConhJqafGF
79LUPsq37G6/cEVreFHW0BK77VHU4l2irnDhJf5RX3lZnXo+ritsnK2Rtj5d
xEqxz0Dgpu3vlVL8H2f9ggtetbjsY6Twrmqy4Rl30qxXzscF2f/QZqLXrXXb
lvvX8P2RLvJ9TPAmUWuio3LwaON3HaI7xPI8IwgZQrwbxLTg0z2iQbeqOltu
qmeUr1mNZOi0B//F2ejqE1tabDJqA+dXIiyUnMvjLaDiGjIZg9UAHb27dIKX
FZoCp8OoSx2jyuDHIQ8/fli42R20BPSpQfz9udI4rYii2uWAnGaXFKzGQmQA
IV32t3Se6C/7J377JiFk/7GJMmKYAtGcX9rlk9qkHhiHV0WA28XY7SjfhtoS
Q9Rk5UGmtQ48Qn0MZC3gYYfP4crS2rcS4s1Ez3gheRri9dpLgW9PbFmUjkwH
EiJ0IjcTIuiyAHLHFnYbaToSC5SpIVAZE8i3MVk3+d4O5uIrB/tGAI05qqmD
0yGM7/ZteX6uNEufLPMEeJVQs3N/n84dKj3XiDMXVER2bqgcWhJimPGYkLcv
HfPTLwaJLAejtT2ygh5NWGHDMHHKqcW7O391KhdlMbnMPJ2on3zBpNvyF9C9
VPKnfMgqD1U3Nk6aT6D3mBiN0XDyhQPlZywkQwJKQA+OqEZ8MgSu1GWCI6k8
d0luqcd3knE5l57YuAn+sKKrhQDPXZzLcze8UxiESn7S9bwELG9KGB9OHbHR
8ucFWplMPd/ecipv6Dx+0/icSWNU8LoOMFGGn/z1DTIXFB3U+gxEjT3g6mgH
h3Zi4YqU0FWEQA5KrEgiCgLJ+krLMfoCl7O8wsS3vXYywS+S3kPGKHrLz1Ty
4ACX/F0Ipf2NL4QpVQd0WH0fyfYFifPesjOT1WZCA4ZSjz+Y6TMx33vlT8Ke
kZ00TiVlIUO2rN8q8HEi16L7VeIisSAPkkhspHdr4UQJxjWVsK+nBnHsUSUQ
jn9FetoHniJGpujB+7sJUNOaKIJkPTNyyDnxfyfQ2mJwAFmribIBLelgi16c
SuCpXMkgzyzh3uTkBz9aIDT4VcI1ixIgUvWzPy9cxm4fGoJLWJ7p/mdTwJr5
s0duHhQUyGkpsSMSyeXn6yzGw4t+i7VU4FIN/3KrvqEhZS7vHIDeaAT6NGka
usqskdVI0s0zwCbiPazL4vEKOfq7L+0fMpdqXT/7S5SOgg5Gg2xT8nU7amEs
LWiJwaPPfb800mN9Xmee3jDYa3L2sRrIY5UzeoCGpfyr4pquVzdG0+08FpNb
oEz0cMiDr3MySF/xfsD6QM1ZwlIX/AnrtAwy6WB1mXuIBiRuWzlH9YbXnvfz
qBkw1R0Ywvy3izYh0Dcy4uck4IpfouGZj5FSNs/ztOlBVl3yT07a+MSYCptZ
AhkjOeZg5MbD5nXYXbmiRWVsTxcE1AvA2Mppdri9KDv6nZqwr3ek4PJ6AxPc
UHRaxMhqC3t3jTGlXUYdizIxgqgiFBv6ASKZUD7sZUlwrPnl6BxjFF2oMDIh
lJ3jxQ1SIu3xPJylCM7k13ftZrVagVBXR8HCz69r2PJ1qh8vjp5IgG278O0d
mVA9vq6ofjfc7CLt0cm1oQfR66rlzYYb+FWDfRl2cP6L9IifHN1FaDXTAfyM
4pA8seKv6pf2blRGQxgALuCG/VzzjPIi7PG5iNAHjp+PpMd7gpcz/qCEMKAs
aIzP9hh3GBfhAl87SiYMJlPznxtsVDHVpxpOeymZwjpmCOmlskI9jyW1gMLk
ZpJqVqLEdZxUr9tjuxaEDvH3fYO6flBla0s1M6oC47YJBr1UJaemWMrKhDc/
QNo8VpoViBmbLe0OAEJ6aadYAJ+xpoc5aqMa/rmxZqN9ULZgooeRg+K56Yo3
jAmzsUytqwN6Jizzyfn1GFeOAqOFGCn1dd+8vtP0gnHW1WCusQB+r25EBq/I
N8g2ei0GtUPwUSFrkHw16sRoNdI6iFYgyW23YEmComX/+mD3NY0OAlacxxbO
aOV9ux3NdSMUE27XtOpaVZzSum0fEmir0xW1pUM/O9/bvJSFzrkTIDBTEgIM
Bck4+7DT4xRH8ZuPHFDe5xGyWOqpHkThp+yNA/Y3RPIP4cSb88KkrKkEBBbA
4F8iliN/qpAy5UL8JeNbXFmYQWQRN8vd6MQBWF/thUcvchB9j4WyTrO4Fj8Z
n6XJ5tIOxAMb5dzAH1JpyrcBBpW20xDEh2tMzbwyp47OpEQdm9XlOJMFrePk
5QKBrSbPzdZ14/T+N5Y79ytSVzapHeuaQCrZ3jpMYxxlWXS2bvGG55Wbwpo7
YFFH7YVPBJPBchnrK15t2dFUoxZfiZO+lpUGy36U246lbfRGxdbrotuG46+A
RAkoKPJFigbkLFt2C6sUNAziDlqhcCDPBF1uQdny1x2uiKirHMON7EUZifB4
TIvircwJMha6P2CGIRofby3d1ItDoDTLS+bRahZaOSQ8cAMlTbW5YgbxcS7O
qCltBHoPDrbiwgqJc5OetYftSPt5UXjPp93BOlgZCEQ855TPa+DHBKCZPCVA
i2gC/27/JwLKq7O5BcFv1yVDRgl0z18jm9jInW1w17LC4LUrCFpFGik9N4li
R4zJ5t5+sFdDCIkmdostq4Kl9Co8Hsna+9YapFuqtQiHYUAVLg+y5OAgRFel
cxP68GO3izMWEL9xjM5HHTpYQEWU7kd4JUb8cINdh0H11xcmY6H1hXMYUNbo
GEfH0BE6yBpd+udjaAQdwc36l87kjDDLowfjoEVlf68YuOxGxggZ8FkTZ2nK
3LhofFzHuHRV1dHXhnbvd0HKErojBedCGXapQs83TJ+Ab/Md2w11dVe4ib58
zG3GH+MZ+oPdWJPK+1DQWapM8WumxNi02vSKmYzIhFbk14ImuqkT1MBI4xmw
cBHMFOJuHi9Z9fmyPjKb79uYzJ7zIHcgsoFtkqLVGlm8Y1O30yCi34+6fq17
HUHX4IDRzSZ4VQhggw2hRnR3bLXmvOsY5XRlCxMdX49uaEbToO+344ABEcj/
bECh7ud4nX1AVi5L0XVXvY0gw9wKprOeojaluEgjBYFyaWXCwrkXdQL/hOli
vGNe8eqre9HUd7Jtvzwvp4ybI00YsKW5iDzspH6TfQZYjIiumk2oRwO6P2m5
w7FvSP6Dr70UmBrBRxXDb1Zh8uMsn63jxQEaboOMaRUG0fLy9D7y6XAOaWNf
OsWycE5HcJcNCAIk621UbHS/OnvVtmRLQ5yMFiVvIsf3JXePy++6c30Q0RuT
S6wiTcn7CMZv4rnCQWz33c5kx5U6/QWMgW4bR2Dys5FHVIJtcoigrMqhh5tZ
b5sWJq60aVjDIuKjQKFKA87ZkxX9tSZSZ9IZYZPC3sunBAzugPEovcBiAyRo
wQC4QUAjBNAhRXGC4oESzffbwXTXPoAPugzedMfdNg6W4EPNuw/7vGpGkHoQ
Cc0UvkRJ8E5Ri3vDPfP8iruD3xJaL0vkFhJF5qe2LyAohhBnVpnZDgHELs1X
j0cfOoaWQ5NZydGq6rT1DNtBHRGAe16V1FOtc9cJ5Ej0NBZHv4BcpulqW3WE
1c5aA77OybyPKveb1Q0cDDPof2K78SSXedLspJ+Zi/NclSX2tMLUAbqiGsri
GUWctwIinYowmKdgZyT11xNsp6U6e7FkrdzXGvApOARWNrvUr0Q/5rEvrInT
pKAw8Hm5vsvruf7a8kwD8ButNtwABSETivm5CB2ShC2Jp1MQ+/K4+xUe+dv3
tqniWRf8nGPJkCo1ktLca0j/5k58+SUNlFLvd1/pd+yBAzkrSbWGWKDYeUC/
BCdjmpdWet6jndqdtpW+47zpiINxEP8yJSQMXvz0D0li2za6IAKbZJC7HbYT
XMwLb/NK4bTLHjuIJwNtxPHsmHqCp3Kgi1+TSMSA6WmJ9XAJF5cROGyWPMi8
sw5Z3nVEWyfN/LHAWiKfHrWulQ1EY72GkUyQ4Vo6wblnrJSvM1JNyNcdCF9J
SFq04urpZkAoJfTia8Luwp7hTObc46M7hNmmtK6qE9a82JMLHJ9dOQf5VzWt
WyFFt6TOa9ELvzKdIcGyF+Gzo/AcXvCDr6/zbo92jRDW8VOQk5kEi5fOgK/l
+5Tta9c7umcQC6O+tBwlMB2m1P2FzWAgXoW8FFuqbWcsjBsVSAHf2bf6zmuC
nriiQJYedTHjK+JRFdgiNkjwIO/FKryUs0KjZ1CQTH1qxGCLjR4zfxDOeIJB
V25XNQZS141fFIIM1fBp409FNF/HtEHaViMg/Rwaptbeq2GAAdTLDERmu/iA
qL1+wDDpgRKFB6WuEeLL8m8LQtV1kX/uVfB5ql1aAcfE+0/0tskDq3M2KGbH
T9j1TAWFuJdda1LGDUuFJyaea1l2JdJwEMM1otdq9UU68tp8rC/h90B1EEGN
C9IVkIkh0IutgxZ4/wPs9Ptp0kJrj5Si9nz1V+HJavg6AKUZfz7yuXPyB57B
ZZOzovXIXnWEnq62F28F8ydUUtsdsYkrUWHsAOgpk7iUhPZORxQNSqadmQEW
pq0oglElLL5z0QHx6XATKgAx9PQSpGAV2bzsreW90Gve01ws++Zc+YQvnwv0
Rl7SmjxxUZCnuKX0cOh5NoUsV6/O7AcVhDiRTDSGxGFWK+a2DqJ6UtOiVzm0
s5zwk58NUMO4Icnw5DROpznZWf2J7Tcyp7iB70/PVP95l4OhJnoyTpZzKtNJ
Lgah0mxpQXMd2MI5IjsmgZSd3tHHwthNCpGQGZ7JsoRqokHxtWzCU1ijPk9X
rEOaGNuKH6SILgWI1A/mHz+4LVvrnT1mlBzBztNCCDjo+C3JChAOkovtPrpi
WwPkWnX+g9yPQZQ9d8URqa3DKd7NTwwV1H/Jx2vUNIil4jQ9M79s2jrMJgcE
JS/anNaLoEUU72JufdACDfGyNpAmTfiQO97eARIF9+vEHX8bSC0QX9AfuiLk
hK9o0GamlcKZ47ptRg8839019HG8GbVEx8EkIIRy8KMV1WlwGTcP5XfOYGcJ
GLGOWU6WbGWp5kf6Q1vgLm31G4dh8QCoC4+P02XGlLxy/YR1z5asQH4ZNowE
WqiUvDoFpAtblTw+dNmdXVPY0uGP3YUb4v4d8X+n3vtdArAQCNH1mmf0mGOu
YR+NdPohPu5mzte9d/HUMRDk8vwSqfLM3iASNGa7Qeaopiskw3sOVjaXn7hG
3JryMwJxGik1fcKoywOrAaHCHJSWjYuSpMfEZJU2T9xTUbIPTkrnbhszdSPf
PtAyOFk5na4VeFangxe27yn98kHI6nRWZfTBK6xA8RTuqEZd354hJH5Fbsn0
6q5mxDb5jAyIwSlz1L50qHp54aSApQdRbCm9zn/+xxCXU6OZne+KvoDz1N4B
n1+mGWmux7A8iHQ+fKkk0huq0n9rfDCig+Oqpu1palhowSz+h1Fwz5vBbef0
b0/rbxLGL5+EYo+Gbh0sTDtPFebj6TlD6F5glt7kuf/chqxuvffoG7Ah/Xf5
bgARymUrJXaMSqOmyMIHg8lNwZp2XnADfioAH1qV02Fmk8wBQWren1Z8gAKd
KH0emlYaHiUP+Wc1VQBn2EzApMJexoohtbrBrNlWqhuPKr18NZ4Qmt7Qinet
IvWrDlJ23T94LcDzhFSTyLq7Ci5lCdgtaV3xUyePMKPXkapPZAKlCMUmZQ6o
ObCvbGHvhvJM1ppxnjV8QoNMWM15KdasAkjt0MHihgxfEz2M51O3azbe4mf+
tOj8sizZHyNsla6Y8ouRGu755jGALXfx9qqGa8FrrlPA0Dd/eDnoQF7G9Rid
TM/GXieI1PR71s6CJD6EyoHotqAdqMTlHW4lZHWUGoMLDPC7YmOeXZYWy83/
xXXrHMQ/jXcOA8/eyn3WsVJWh4LqjxHIYgylFajyQ4yF/BJWjHXYUjIfPWkO
DURBpJEOqG8hLOUHf7TuUzdgjj8SUsXw8878jcEP5YgldKCvYg5fZ0bOpBRQ
Fc0RpwqHMbqsz4KV2GeV5EUNcSnPCFYcmgpVBN9GHSS5lAPojC0Art30M86n
mkblhrtCEZTkq0FQ3MHckW3V1Y8dsGE1GiDzzUPeCBYjzaWZzMD/sVngrEdL
fO0OHW9pKGAnS4qMqWnWe2QoXb3Tg5Y6/RjUtT7laMVyleZeAydkcZsQ99rz
80mi/K8DyUhCJc1mo0pr2MDqKm2n7iH8pAGe87qGiUKKv5D5c6WXBEjyRAKW
SPkc33ZEb+fn2fItCR7Z6vooLbCZUB6ectfTtUx93U/ZzVJV6sS5g1Y9efIL
3OJgcx9R1hJAJ1gbFQG8o2hqpO1XcdRdWIoALo5X6VFWGgGo2T+aawsj+DvP
r8Ssd4nEPDDB3yd8I97Z1YQJEIndVYkAhqEdrIze0fXcgoMoQ+qmwVryxfHz
6ZyP5fapIW2Wvyh+Rb/U92jh/Re2OcI1OzpllzlfWdty3YfYu8DE0Ndjoj5u
ELMYC997gQP+hL4gy1chAO2PIVG8auHDqSBjJ/0NDWgb9PYFe4kTnh38WHqV
esodSDOLwG1X0WvxFCZijuuPi4zIPbjQKV9xV3SFz4zeH0iucRg0HlmNInwJ
kOAZ4LbSQwPrGU5wATYcqrcR+TdEE92xbK3mvRqpMX+1+KapUibEvMF9k5WH
m2rp/kKEDUbM9+7GGG6Tb01pKt9wfSCSDr1IMlKIW0WLQmWMgLcUen1AqgOE
qSvXZzrgm+YbIRCmcXpGiFDUW6Uez3kOWs+Om9GA1K9FCT+VrJGp36uaSidq
XgGQWVL2LeaEByLETnB5Q6LYW6OKKGtxM+rGTo/T/5pvlHEK98WATaSWCueD
UuJcmafgpWY5pP4p+D02LCWQ5X9MN3bT3hPUFx1qhHJu3xS8+kO+os+Yfafn
Nm/DgMywAikOTZkE/lpccnDqFy2etkHwsGQ/Vc1Ybs//WQIodw9Zhn1bXWfd
XV2FP8vlRVtyEivaPGEB43I+ePtLYg2Uc3CCLMSvbsECqil1Z55gEjb+WOTN
al7fw8cH4TB+VTqt4ZkE40CjS9DVaZy8erH96a0ioIKffONttbdjCf9cL/sQ
HoC4ZXUKQehGIPyB1EuFQ7lvY8QIDF2qppQX4wmewxvvPj+B2DUEjKFlfg7l
w8sLQKg51AdlHJ2IQCix63tsjnuGvgLudR8PB41VMPqGBbN4q1QzbhHH+GSa
4QTRQJuDO77sVZecnC1NN5LP4spD8R/AHgSqV1R0y/EyrJEou3jkD+0djv3y
xO/U8J5tIw418U7p08X4j4zFPkpJWq1s21wkCgYeyT3r49pzyxa6G7WKIPml
vLHwkXRB3bnwsP5YtPSAbQL3JRI3f6SUOOprFmV7qNS0ZqH/WO2OdnEKm8jX
zINQH5yU+20ym2vXADlmxwVfyieN7XYareWGt6LIqjn+kc1v1wox49cPcs0s
KhNWeSzTtdLCDOLwxolnvZjdKhLNVqxz0ojJcqtiFT9VecAZw7BJqwHfVAb7
QE9IRhfBwexR3S/BMeJS6km/ORIn6qnAUTG0+mHXOo8eZJSjnszlx8Fw+yVv
ibOGdtqgQyzoYRStp+rpAfL2dFsEuLI/+0eSHay+Gn+5l9Q/Alus1Lxt/u0w
L6vhRDWeQve+x8YCFewHb6RM5cbmcJJnu+7sLBeBZ/gis3utgegpNDaDBL+S
rQzW6IYd3DY+8hU4+tRJouylKh2nZw/IyIX+NgCH0sB+TIXcG0uR7DpM/GHk
sbZ3PCVsQXM/laYZFOrm2Xu3aMJ46y5fJKQNIc4r8/CU9GYo8hZrnJf4pzxq
S0viX62gID1yF8MWW2jJVqHmqbrAWC67OnqNGzXi42k2ln7E/vlWVzxetTde
bx4s65e1NEAevdgePWBKM924JObIZderOQrT3LTcdXWRXCi7jHPT/nc6wFim
m609INDi4TOo/0nVnhKeF0nQBS++SiyzF0Fhc9gJDV2nUL2QEI+SXq4PIqAg
CrdZHGemlwmJsgS0oBBVFGmwHuIUVnfbzr02HcxPiEAZFY2VBj4B2f2v9o7D
q9tzz2NOXrysiFPyXqop/lI6XiNd0+mx6TMLnG32PCVpB7MIBl1Ng9dnfD8O
qvKc9/5ubiiGZTzVGfaurSxn/qKK2/0Z4fCzHdrgM3FHDmrryAq3ULPX/Hf9
0zj5t6Tu9nP3rAF58EwcjWqp/kv4Glnnq9inRrZW09hMF5V1o6126zvwUbgM
lIem3uQe3mVecu5XRKwzb8BxdrtB9+CFeKWAM7b4rFaGmFtCFISUqKUliV5o
sigvnr0rBKIyJpouNuo/8lASIBHRG+HdFod+9HwQ7FulN7zpJ+a2HqOXmOxZ
T7svLSZ0RBykZXCB9LvJ8yY4alQ3I4FN0uSUOEYseuXB4TsFG3r4oOG9txee
ju0YW+2j1QteQIHu/au3h3ec1f8gRseCiadvCQgzt3YzHCLBYR6B5WmWmQJq
hLHy8IYHgaC1WYr0ZjbJBpDnYCYNEnLmqYtwwxSRDeBqtb0Exd4RIG8yQHJ8
mg7BGkX8XhxK3AatTZQzL/+1BYIAJGBWPkyM2R3HAteqQuAucKKpOvmABrBZ
QaJ2NPoPkl3NAdY0WXiTytD8cY/jTSd84KgTbuve2GvKnUGucny65NffrDDx
a+Z36SDHJ+N06gw2iuI8nVA6eav4XgTP3eKgbGL9s0ai0NProvo7iiNEe+jA
qjiKj6BZWQ1FnEgvElrT8FSBL0DcOEisNjpQjAY29BNq7uMj46IpcNoD0UcG
x1HombE/ottZdK/P6XFVbNibm3MX9R6tsOkjDw47A4B3ECWRwEBw5WJUofqu
hVZohiO/+nOb6X3VKeBm5419T5PuBhn65x1GAf8DO08CAOe3BjPcIQUQMUUm
FbuxmfoKyl50b6o8lQo3DYbzpyd8VyBAknmoujDe01A0c/7sdHS3CRsxg7pE
AyoKsJz1n1VzjJCYhzG8a8+/8h5z0aMWERpNxCN9h2IZF6/VYgG/oHMM+K8m
I0zBPMp9Sicz6WipjKRq9ZBonKsu3G0bTaixbqzD8smf5SPWL0bh4yjqbOHS
AylXYzcO847yPvsCYcLO3h7+10O2aJz1CfHOcFM1E952GV99HC+I7ccN51ts
6d/GpW6gw6Ipt1s8vx3nCfhf8hObSdBmCQDI/wN87FHX2YsH8vIy0AcOJyTy
TneWqJxwE522lxmKbaA+b+ZYFbw7DTl2FATo8/J1JZOqXRqyKunscTNZSJUw
969YI4asyp98La604vXCwnxjG44hLCzRvdyRlwCRULQCeImj85g/lDSgfiUy
hM2QnNP4EBVSG5/OfYRJYua4zNgRAt9Qk2GTYNA0AR5/CUCkvBsjq1i+aq9V
W0q8A0/bXw/Xno0YWKkSoMZ6fsun0AnLV9ea87ibr/qBJrI4PduCySEdWTVt
Ui6R1+rZWxxTDIEMVICWRuRbb07dGfU0+BpSWv18hK0JmNirv3DMYX2JH9xf
vc66K1KeqXWBfVUt+9LuQnNR7OUYPVL05O/+wOt+NHTgOX9krFSh78CJs9vd
4apYNfdOcBlGUM1L2Du8ikXKYcEXVtpCxEhbjNt932AHUzyPcUJpUaxFjf60
iRzGLZbaocdiXcvag0vvWPXaESNv/oTzs+Pg0bZJ5RENpax38PFTPg07GWH6
qGea6TP2UyNxixm32DirOUIa1GhrjIKPid3TSPgqTP6Yrvq0YWHcub2Qiar3
RnIJKZ7/MZcgstIGZnCbw8aJ9I9VJEnB612i5Y7JFu8DcZRyelL02RVkN5lU
CV+H08MUYZFK/CShGkq0lAPfiWcrvgKvnFYCK3BQ+VRmCFfWFM/CC3uLJkYd
4qK1HiNEQW9ihbQ6H6SGUiON3CiKBzC8AN8r0Sy6T7r/pk38BD8ouuOSU/hU
hU0cMj60EW8X2GPuwLmowgDAl2pMazjYmHkOR4WZtmu94sB//nkU6Z0TMb9t
FcKEzWD7R85Diiza5wNpd99IG0li/2uVL5w07tWXlk6fMl1QePdYtSbYZwyE
wvQsEinuLa3dkklT8objbmCrtAsSKlLTxypfCL+a7epSIxEgx2RjPRkDGtK1
kpkitVp70gby8j8WmewgdFYCS8Mokb0/Pl09qsjQ7idnSSjAfsui8V2kOG2X
mRpOKfD3lurDBEhpZbiKN7lyIVCuoWYdKl6tErUfvVCpXr9yRO9sAFgCabtP
KwLb47X+E5KQpRFWX/TST7jejA14+LQdwhYT7kx8YemWwm9jO7+TSlsWrqmW
4OZ0hpjUSHvaJGUtQWzsCR7j3r70z/LzW/YKMcUag0hfLSBcLPRR4NUmA6MK
PIuWH4ETbyiWn3wXLu4e7Sw+jVAgtBac1VPCJ3Az0sOAXG9sv6W+GwpKd/8o
DDTaNaVYHj5HrN8Fv2Mr9OxwmDxVYXmIfCZwXqnogVaMEjltfQDeydmzntyA
axAxXhpWc6PXilpGRxf7pLd8RIUgmqeF+eSfLfKzd2jvKM0vsGc8o6OHzWY+
o/OjWpMbpXM4H8Z2rF36PcwgSJZw8RS0DiZYl3VZSoxlQhJi+Eb14x8bp18U
GNNwDyG6GnDfIsyA+YQhzv7wvtGF+3DWvJBMIDUz/ag1Z622NxDcs+DNE6Ct
HQk/AGwR0Q0A6Il/pkgv623PKvkw9X8ynWN/Jmoez79Gs3BrStSses7ir/4L
AveKPdn5EojSo69lEEwiTOJ0TYZTDIuoumq1oSMpMFsGWRsXCAEA05/jvf4L
oIEA6zTTr9NkMtlXzPE5xWweqnkgGTEcKxenEd9SNkACKIutrjAWS+XkQT66
SecVD6wKLwHb824Bxg7DpT8L2QLOMcTsK/uL/SnyC2b28c36PmKXkLazJ51T
v4+R0EML+5RtZazbLrEoavuGmLsZ8wVjju2bipXpJtHfelYELLo9IIQlxqCt
mvvMglvj+FoCKMBZ/GP76IAcAdS82Vin5cQXoX+gRO7cac4zKAntH7CIrMFs
1rJgaJkxc6wdhPUxAOVwRyWWI3aYHj8TtzNeGk8S3/Jq3a6wJ2b3EpUgb5mS
ik+LMxYFhVI2y8XpSdoMr5eYjaUnJPfprFbWu8zlV9muPnyhepSqaVCpKGwx
zYGBhs1T1ryf0FawGusBYs+CtgV+GA21YmxdJVWV9XhjivYop6ECQ7mcggzo
EdZ3aeKw9XRJcNPHCv0Vk4uDo42/I62GHBugVugPMYYwTEi0QA5cv/p+IqT/
deH+Q8bLatfQ7XBSeRh+V7POdv5yRviCXfaMYs3BZDnG/y3/CW+aYwai3oNU
yNrtZVbgwbGTxGFDqwFXY3yWl14zC1IRB3fPUdlOBZGf7N3aw2bm4r6JDlxC
irBOXA/6atM5fPiAV5jiWE/YTqs5+XVTW2l4E21n8e8i9U9kQ5sEiR2c6GcP
GNS0XZqzjRcdF+6oazrw+WTn+Ef7jywAecHCtuM5Tujo4sgxWorLBJA7VOZw
k5+WtrXccTI+zy45Q5WYjXY6W931SCfjvZvPMLGBllcro0oHIHDedoIfmhYv
uqsaHy5z+TNthMP6Vn7oPSRy2ICV8bvPKSkpdnbod25mNy/U3AzcUiS1O0la
o8J5Z6w5ACzL/f+NqPxbEzSXK6rXExAVLYzxwkAq3r2jE36cKsNgKuQUCwRE
asjD6Z04qn4bDMv2oP8YE07o4yG/xgRWQ/rDiWsVTLEi+XOwnZrwnR6k6A2n
1oZWi8Sq5bNfXHdC+2dwXZnkWvCB4d/qU3Hqgl7BdOkCA/7FGoqYm/9OiYZf
ZX2T5Bf8dLv8Aq3HUqLpkAaKFsjaeHukfv0JYt+vfqUVYuI5Y60+PCnmztwc
qKpTCuwmtm7tAgmrZJr+sg/S/An+mFKbYVQWudy5MMpcbe3CHAOBk2npVner
xLH8ncCc45/Gi0yr+NfkgVCqtANhMgpbmeEPBb8t/3MKBzgLsRkDXBEMvgl4
BNsBken1U1ndGoTm+ytr/m0QpRVHrKA2HeDwfh+FAyakEYyc0vaClchhHa1l
BI34LcceGDVSCs7z89Hh/EHeDR4JK3E+mGWlpx0lmOSPlseypeWIRuvhEK1p
p+pYPoqtMroWdgkTaOKoAYKyw3d7cNezFJtURjUeqAGeD5H5sxIFBG37TK3P
GZhtEdvW2th6lzNFdux8M3BJSO8TqE/KYLXqny5/J3jJpfFNdcCcOzJ2s4Ib
0xUOb5uqj7q0FEcqCn9AbEjKq/dO60dWH5wF9+QNFATplkJEBvXEQefRyKyz
JZ2Zv9yTTIl6+UQicLCIAle9PJJbGdAtSLFcI6uASQT2NFimMjAhopj5zir+
ShEUm/farU5dx4pfvmnuvyqubwTV2drEquQMtY1a+909HrfYSqXMx2pg+Guu
n9w4FT9sm8A9ZcgGUZG8b7tJ7tPE/Hb6t3Y5e5Id5JGg7wW1I1m2NWZVlGcK
HlGn0KUIae7ZoILSa9LTYvWG/l0IjWvsRctAV51EfOYBlSAtpYoB49akCdqe
pGVw5wnW6e/9dHeMgzdFW35YNGrrh8qwsZWhixONfMEPMv+wUlFG+5dO+qY5
h8p+/MpduKfSSDuZyA2wH3O72JVY2z+LJUnOjnNZyzQjNDrOs1nnOYIsJ2WI
LePRZNRwAN7nyKMLq5NSPZ/4HILJAOjaQH6Fa0Ks0ycjt27uK0Q0SOxgAJOY
xMnvYF4j1aP/RFcjcfdaJdW61tx3i0GKeotk91mKgQqIzcJvs5cDYuWvzkIC
QJeTZwouFrEvlXoW4FQuuVJjkG5zdHDzWnVJDojBdLkGCEeKz0yaRVDhSMQe
1akz40ibSc4fYYKoQhvLa2FuTT6j6ifzE//Qr5AaKBg/0GPLwkIttQueNd9r
H4uA2EODuO0NMJWqrO09qBgVzrfJs8ET0qskWXsfFXo8bhxI5L26zADDTq0y
saMKvBe9uZNMu6a9REwGn+dp63IOMr2jM9PtCCHeHxYrE13g9260YFAceakg
qulkLxaTLxDRtgOUox4QHNMCGcu/B4QXLT53Qmol8ujo2F2UlnKXpbewdhDi
eiB/mp+alEPkxvnaE0xkVSljf9e/uxtgG6isBCtFW72z28B3mlxDABR1OPZV
coedZvxkXe3pnxhypiqvKZmzBkCFX896+gI4Gkay65fmsWaee5N7eknbsrhq
Tuez2UtkF+DzbH6XP8SeYVLzJsqZDa2G8j4GxKmcxB2BzDxA27mduYIL6YH+
apAAO/n1EnDR2/8abMAjFv9LajnBhv7lN7Is6Mecc9Syl+g31jx7oWTiHqJE
ix9ziKIiU7aZ17O9DExIJDp+ZrZbIvN2pIbgjUQDBP4TI6KVY0Zpo+3ou9Fh
pPvC02MifiByFtT40vmJCfTONR5/D3U94ZPvpe9lzoKVaiBVZ/h7zymAx/AM
5yXhR2d49/GGvSIoGCZNPviXhH8ITXYw5l1TC0Zpnrl+vu0gS3j/M+6Fv8Wb
r7RswEphfQetEF8TN7UDJrrMsCIgrSSe+Oyi5HieyJ4ZG1kT+OolcWQBCsDh
jbeop9URLtrr+eL6jyjmwjdBq2NGxyo9K9h2AiG6VGOnGKKrgcA0fUV4NzFU
c0JWyFbWGQJrSs/s+r2U/z/xtbjt2wm525EMt1RzVEFD8bvIQuVMoySg8whg
rMBVcDiVe0jL3V+wTiaemfdn4RN1nsEp8OnVLJKNixGjgTVZc7+rXb+mAh/G
rLg7cuxAQZGsdsCzTJfLK2xLU2ll3NqlEyn2x7K3Cz7Fr7eKqyIGI0jgs3TA
Zpf/CCZ3z+Qs6XAncy/4yOiE5r+Dq04GOtijqIjPf+PlXQuhxvQOrhQr+LCn
8BJ8CQilA+pWkHZuLeFTu860LRS26V0DFi7xxGZ3LetYoj7j8nO7DoXld18+
YFO75wHPNfprGKRBUd+LIHlqO0i9aPJ9uze8T2UK4pdmU9ojeANNGVpPRiks
PrP4bhumByhMVPo3rS+JU2tQCEAcP/Pf2eLt5i7KwjRxg9t2W7aSZvie0ZkT
R6fKG8z9xfFUTrSXTFJ1SS1WLZ6r1/VFvU1JKCQhTLKdabz0C6gniRBjDN8p
F3wd39sDFe2uS4E9vLWaEdLI91A0LC2jGo4SO1aCHfNgyhmb8ba9YNt8WGcH
8urpDtf/Fo2SgflitOEa7j9n/EPgNKRZb5+JkKV4rfgGHbjP3Zm3BOnrZXtX
oifTWYUSamaHlWpwqE05cNUsFy+E5n+ldWkurMo1zBHAzMYggvq71Q9S+Zzb
DMN/On81CCZ4Su+fZ0Eyz6e/7R/TxzlDQU6TY99UxU1MJ5ztHqRoHpWXMNok
J894rVynwqTisB/SqQemQESlUsKYpQbUHuMgUupyMmV3E+YXzLPUj7FtbP8S
lp1nZr1mzdZQ6Oe9iDB3fED+7cqzlM3uyZoA5ju1TuW8kgOOa+juxWEF14Vb
p5wLOcYzgdhv/aFkS7zKdJYuBtesaf5EqpszrXklaW4o9cUJisUir1jMhyeP
K1OMyde5S8imq7SYFlksz6dOaCmzo0iy9iLI1Ei8aKQ/iHd3Am0aCO//k38I
0uzkrn4FnqsIRrPYTq4u4PevFzgLkmwynm55qJNgZJJ5qAZLYLUKW8LmwWfh
Rsacu7QKBpQZISNJv/Bn8CgyIs+TObV0YheiR8sIrNeGzhoNbox6c7tTL7de
mgaQh4i2RN+DCucO147vjrw2UIH6RyMA/iRKKoZS9mAkx/s+C/YSgJRk8e3G
SBZpjdpeVbBknK2ebLJykMWqExT4zO5Uq5tnpo6GwaE1KTgi52VkEkUHdIDI
CkuGoLz/71J6Cr0Hn0RwgvI1LGr9XdN82QNKqXIHBLUn7V3SC6j/DBzqgvhk
rQwRY56yo0CPNHFTOjrg8cxo7b+YY5/6EzRk0A2R5Zextd465sZ5MCRlsP3f
MiaDklpP0OE/eTQnYlIanPrP17siZJgXRMPFDM1SMBrrvRKc505/r+Nla0dU
yCCxopEn8yVup4d42TTQoCFiaOPaw+aosYyd5Wnh5ZSh6xgZ5TZ8EX2cwg1x
t1tos3wtwniMIPkw05tdr1IrwFLd2B5moPD2j5h/4stvScygfn1gv3sdpJ5/
sXi7J2ek0QJYl39o1hlzmvz6zWb7KD0elA4jygRFoYw1gwJSFHXBsS8xNCDU
C/myeRm8A/8Ah5FUl8aa0pjevGQfaqC5n0lFfKHmcqFL9Z49C6+Rr3Qgam36
lg4/1WolJpJJEmnst9/FcsgZQXl8wHuYAX3dJlMiuuGy+4YiCOGWhyve1Vkn
ytVJOp3xiDyw/uQWcKueDJQqb1wdvFimfU/1ONyIY7R+Yc0Pg1g4BjdYVLHZ
sHXXRFMnXu9VYjIG0l2LwB3fH6n8sUD9wrmDs6C9J/v55gl0GJsW9a1aHsv+
1G+ggs7oIt0UHSdc4oKbONR7BiNYfLKcdsBAaT7W+LYAr1YLANLttavnhII8
K2O4QbpghujeGdIpwgiSoTrMSGy8sNn16UI2ITpWAfNF8C6ujnXLHzJxbu5J
aOQaatHkVueOrNHbgv3/AEoa+oG799h6/pQTzlS+V8/aLZiB89muUhjknugn
4A1880bFaVFWywi9Ud85GFU4vqWwxVR1IZr/uzpjXCn4JmWLPcoEKW6Jf/q4
ML1HKkA5WK4r9HHzt/myNPKA/RoIlG8/UCmN7dX5LYhmShitfA3d8FZPX6Pg
EnRYPgnBFa8e9RaRO6XE+//2VPB5SBsuP9E+VtoF8b4DUbOsQsfPj/RWIm/J
uHciL07bra+D6QoZZwuh9jqBsDcr+rRFbX+sHNZSOw8Qow7bYaDzpPY1XwEa
yMdD00Di40sR1eq6BxP6LhNSECoifJSDOjIIMQ5kRJWSydwO9zNnJgdB/nRj
paa4nzHONbDeXmMqvnqbLxmqOplPypkVJtSdOqnROg+1R3gk8Q0o22XMYy0T
b1iEd7Re5r0uwtbDbgAIsrHGVMuD241U+yGD8dpRqw74Gd95gAph9hxNZIET
8MVlS8H++VVWh3a6jHPgw88EojcRG6jcT7vpo4PL59qw+hQfnUHd/eIW3sNd
WCADxClKV+IASfDDirvWuDD3ckblV4bcwiC/bR0jYlkpi1+V8zGgYBihVAiH
WqMun3A8/ZbjVnznzIgvpmsBYXJXh2J2cPjlDivZIrnFe5MUWN36hwJrKOHx
yJNHwr8eRQw6LPffnzfSq8Yz4d2tq8T8grPUHw8ERXXF/WIs8oYeOr7oSyIo
HAJ7WiXncjHL7mWLg1b+zlnZuQAo87e9N1a0p+FMXmjp1vi0NXxZ6UfSSapA
GrVpnSiyJiThqq4rzNoMre/oB+tiS2Ew+oYRDBgT+TT1J5xTIYal8ttlrRem
S13jXkSQCvZAgwMnNcuGdoHqXaiTgZLJIq707DdI26drz2qMNVwd2vJaJsHL
WWYWBfrqE32uSGakdBaYGBHyVQkBomVwEQRIw7kHZTwVtLtxiWLbMqLisutO
H2clfiGVMSMqk+8EKemD0RbPht0wdEN2B4Y0QNuF+6OEpSXL0cRlSy+9sPvb
nKM5QjiFoXxx0m1X3jAQ41XcPTVxjJ/K5UM5vgU37JCTcf56Kreg300nRaZZ
L2QHRtXZcdeGTlDVqQjLIE3EobgTUQAJHKFIQK50ixf5v6z3yGk2avJn6KHs
M6ldyU1mAkjdJ5e4vhwT4Zggk/wbbje9Wi6lBXoEfeq6EDu3OvsoxnYZspJF
vbuRmU6LTLgHyOMX9AlnN7fdp2mmdq75v8x2UOd+p7M92mk/RBuxRXMaKQOT
w9fh2Suoy3rGHH9T/sb8Cx3SRnr3f9KkSErjqfChugQz+XOS3TCaOuAXoAde
Scp7NT+l84QkxzzHBPVO5C2XbcVWlabEQ5W85uAvaIXRI3hZaDDUBK3vEI85
EOFgrbiXwUcHFWl/NkjKRHzHjcq5yec9j4jV8KfYNQTG94iWuHHeHL/lq6Cw
/EgsSHnCvb8u5PdVOjwcVtxbMsX1ngpjFaNgV7n2SqJxmC0OsfcHiX7vE4wn
zTUe2vIrj+KSrpRraq1dbBY53tzoODlYuaS6u3xnWiW7MLAMTnqFQJUu0luV
xB86W4Gw+6DrKct0pKqigSfVKcBPdW0v6uUNe3h6BGu29RYw4Gqi5n+ago+u
zzQYEPh3NmWKUfPkG3JvTPlQrgWWzr3a8EMRnipmm8EMTKJ2gSoaQC8KWdvZ
nz0wu2xq8aUDEuXNjseNqosTSDPDTeyOdS3srsDimewCoVVXpRsFX031sv8G
rvWTD3M9+5ArdwN+t/v/HWZaeGCr2Rc0ZNNo+3tL6kWY7rCjyyWxHy1It+GR
i0YdLuXB2jjl+G3AHCpcIinTmIbtqdL73RenpkEFox+CiG+Jzh4QAmPIYI+h
TJCDAlALgxLMT+k6uc8163pqLbWN1uFHzEhJnBYd0Tg0oWexJFEM0QngOY2L
V4qqdwXW/iczTXDxkbihB3d2hJhf2wkFXp99WigiDsrNjY70kaahg5aJ1koM
rQzevLJ42YUY3zIvATk/+Ek6d/rIAsWZOjm2XBbsut1/rGuBIsTveKddvXwC
i8GkNdSpb117JABuFJiUKz1Qbc/6WMqJosR91UZ+njr+P4YJPtQnunt2LWbe
ONh+8Xc623bHd/khRSUledoXrz9YD+LDfCSNCIKNNY0XM3EML+4iZTytvkUu
5n6wnWQu1p4xQfgxG9vfAkGp/4RIktb8yN1FhGRiJW8XrR5CNh6LhL1gC8X3
gx/F5Jfcu752F9HgK3vOux6OkgfBHIXldVJeW81S9cGea6LEOWzwTmDxXWp7
FHGTMQZaY/B0EC2Q2mZpfaz3Vv0IUTv/CUSA8rnznRnX3faAtxoDyNkdygUW
u5ZuIHdWSOym2kqqDo6A+I4yNHIjEi8HOS6DtBq+AxlnKzgFuBb74dyh+Gvc
9ikgXrR9JhLmnA/wow4VGTZ48JZe0zIN5CxC46e0wrUzAAnQ1pufSYGqOTXA
JPC6QuilUqRFYHML8vZECnNUkj3dMFH7q0k3pDy17Bw++leOoGP7+pw5+hRy
BxgFPHUnuqRtmOTRw3Q9eDOzz2VClt7KLd+4vTx7AOmYSulaZFK0Tipq1eCf
Yqo7desBLSFYxVomvh9aSROUg8dNNhmozrL7Q/MDKAKooye1ANPDu/qT/blI
+aVKeEbkuliOHlWfYC1aF16zttiZ0YGbonoiqMd+iPjZnvbbwHEP0FqYwJ3k
VRwqtYYpOT2fJzU4sa3JLpNF03pBsKPk1sqqrxE5LILDVUnV3ZiE8EBuBydE
y+DKB5e4xupl2Db9NNrrdqD40FklITH1MvWZZmuz00t2v8h+9CF3wPM7Ytc6
QJWdnfhTUlgaiMP/A/NSinLOqRzgEZAOakLLYFDtSE4iJGgolLp8bU4NvrO4
qWMqjTUOeVdVGD07er30yt0mDZJTHLfNi5tFwm3zojBqkIAJ5zZDGJcNx8Vy
Mrg4ijG0JCDrspRWxei8eBJyg5alsbDt0S1Nb8pvhHNhYYGshmlIX88uzsxT
Z7y9xRCwooxPI8kL9zAFdGdwhVPqBWZCIVWpDxFRQYtwzahRGFejIjh6o1C8
qpdwNFtoaZgTIYwmlMhipUAF72sqO50KmiTBZbIicg07iZlNbGt6mR6xjzh9
xJUqoGUKLJOfmWjooL1gUkFRu478fPb1GzTySXFlGdYHzgBavYXEADrGLCJ7
EnjcqY4Xp7jaFvjJ2RtD1EPlUPnax5falhgJD23HQDhmjdIrA4qQoLuVKEiT
Gl+UwXXYlqslHhq2jH2iBsAyERG1bb+rEc+6cHmedbt+e0gL5c/UQyERjIa3
ex/Im96yBCNsEB5eQSSF/KkFfKTnfjs1mXI9ja9GI3WkpQ84YHwoLQCzYEgQ
V192rkNmNUXJGRrb3KjFRpq/+v2a0gjC1Th0Vhn+u5z9HhzD7vFDMT7pLh2i
M7YSDd+lrW1T4RcostuwoaTzrsPL90cdhAynDXwTV+WXxMy+NMQLB8Qs0poL
Rwyn+KuVeobITQp7CQCHT5Z4yE3CGg3VLKLhOKbGsTbB63v0Bqe2hTc0dW+L
1jbKw9MaOwsQm+tQZOZ4w1oY5ylfqcIP8ilRKxcnaZMfMvaFoE9dsNKLBcN4
vuWQVRmRK1oj2tjGwtHtZL9ttOe2AEnE2iBMNiPA52nBYya3tpHbgxNzNt5x
ToKQZcy7iXOYFDVYx2F48kciMaiOiXIn22WuYlk/qzomlU2NHcRvckt0Ago4
QeuELHsJrJPQvJ+/FECC9XEAgnGEngSimtVwC8Z5rr3slkeyuJZuZrdu11ZP
lTMi9iNLSnPgcanIO8FYzvIQTbLf0R8E18ry54tge78BkZG9mVF/5IIfj7Et
CVbNalrGhOp+WXtrODfmgFIyzEiBZc8XA5iJ5IsNFOG2eSzov/hwd0ZtkNEv
EANUy82CdudGa2C/9OZTmQdeAmemVxVdYNvgfF9LwbyzctSyjN6ehXDRyMxH
woshPP2oT2+TqLOz48oclJs51kcnthuDAi8bhknpfw0+l98NIyDIdfFrfQD6
H2KZDcwkONboB3MDnCL3AzN/FR0k9DExBiQ4hTbAf89JaxbBH39MP/LJzk66
q5MZDMXOxtft4fH5VwhYIVCSpCLDx4bOWRYikEVYaraLlYO/o8GuxKiPJnZm
dpL6JD/mf9V6k+uNcfZ2n7n4IgsfADQZwwopKnG+EMuWdnQMUe2qNa6OosFL
K10FGZn8f/39NRbR3xUJHCrO2/mYagRVI0/xcI45WDDL2eyLH0/onHfP85/p
9lSE/TukmJdYV/YCAOt14avWoB0yVRLeJu1dr56q98kM1s6Il3M9z9zRdtj+
1jWLUiFh/fMMLRBE1JZY5bVBb3XjaOIebm/fI3euTRGgAe0HOaSNOcME31vD
CfCJ8VGHg8aDDuECtR+riVbyAG+ueX0YPOruOTS5v3n6kN9U9I1L8KNXOio1
SzhRT4ag9ENsMR7LySllv4902MgznlPKLlvSq8WfNJdlgPVlqb3z6x0fzDI3
z7hU1/fNF8HgtTdI/1VAbtys9UWLeElhbZlZGKz6WIPF3vSZI3cGPCbRutcB
b+E9/D2tgBs/UDfEq1y63sg9LqJBRAJuA/OXZEv3BimSA+Ac1NIIbR55W350
nVX3p5/bBlmaMbFQUyEtwKzZ3gOdZjGXctWBwuIoNZDccRcreDaTEPqZaJPq
vCwcOsj2c3Yc+IgmJaUYWVjxaSK13gfaDXV9da4PAiYD9HJxp+mtFKoNawFa
YAm4AeMCYruwrXgZKLpkHAsdKpo2/C1HyZq4rU6N/sczi1TD4J74vOp4HStv
ERV2AKcu3scVPXd+mo8HouwpZIHnO8SnEM2/k3E4eJOCaJLgM1piBXopapEx
LLRLCH7lEFjvyHry54vQtdtYKr+5W4QHjHBOrgNkbBOIrERKI4toIh5UnlJ3
ta8wBfb31u+PFHMF1qU+td/GJNPwT3ujWgk7P8MyyHdbT8m1hNdrrJOTtbMV
/JYOTzrhcjxyQAmDJ65IGys1YD1y2ZyTblHgqUz6IBXjoCg8mEIMa1EoQH15
IDlAGrr62bp/A6vgCGurgUQPOO/Zk5xYOA/Z/C5GiyEH6NzIiyGXxqYdqF9g
UWTFUkYwMGFPj1aWtKF9gRw8Og0jsX97yhBYvOou+zWK8fG8/1yWpS0uG4Nl
2ZBTSilVM/0sqPaq3HG/XjUkB6RefUNem4ghz0ELTc2jePEGSxH5CgKG1DE3
n1ip+sRD/46hG72dyObVBXRNq5EGYwYql/6adbLqka6Xxwk95in/cEpUJHhX
IMG1ps5Pr5vAWjJzsOBXwjne0WrDS9uZ8My35eu6NWyS7gctQf2Lxii9I/gQ
kEnjFq0q3s38g6K1Ui2WQpE3R1jPeg0HekBHKq4cYtHTqUAvtM/sHm5GjQyo
JRzCRxEbbL2oKx9EH7lZUZKzLxNvbV2XDVZfawEe89tO7yVdHHnk3nS/0cqo
LFJtyOnd6dVaLAaw67nTtfBtRsppMpUNCPvLZ+ehwrE1/Hdi99Yh6SH7Bi2P
5Yb2iE/dc+dZCX8/i8o5zjZG1ndk5Ew61IQeQ1BGkVWbGt9612Fyd83OeTIo
uMeOx46+amfboNEL699xaPSS4o7zDkN4BZYUwkmsWip7s8MhiRFROrtpjjET
NxRAvCZ22dppEI4qJ4FQitD7QIVnX/rjToxGtVYWUYYVVx5zhlEWWElLFUaS
01L3mVs+2ClGCQa23UHqi17zlFy9l1+1zrNyYyUKqV1E1S3tvrBGDmNgTg0M
Gj5U5naxFGY/45akejw6Z0gjSHVbcGj6GGYs/CdfafDN3xF9WwkZl1SILTHQ
kPINemYLDZFloJDEDAz71vTM/iOY4tXPJJxFHUyWc/OH8qj+oCt9NqLl6F3u
mNT035t60GvWTNhRuEUoS3FvVEDR2g031DRPkJLf3So5qW8Fr1YnjEg6WxJy
uT4ZNsJpPDb3lFvkO18pxUP57V+NpuU3vmr9YGdcmbAWOVqJVz1lECHuPhpe
zkLp+NVU5OhlvdeYE+FKh+w0cOp7oTIRPTIWZCGqhf0SmVH9PFMGXeI1m+TZ
X2SamsNmSPFh+co354dkL1uOoHbW5amICQA/Cn0sjSOnjxXNiDT9cr0S3+YL
LEpjK5g/cEQYckP5prKXiW3mpVptnEMu2It6OQVCF+EIMVo0p2YF6pfEofXI
9V8Sf6LpXT0AIzlltaFfS7I7cq+JWDNs7rXDQQsSji+Ra5i1v3VyMeKY9P9v
ZXXYLLqcqJ/AgdLSuHMJ+PCdNBSx0ZgLoNsF0ZGbNHVTrCO5EZLyirBBJYP/
L4NsZiT4H+nsDFwN/QzntIuMFPDPOQSsGJ2kgFbxBrKUZAfEIkqzLm6nawE3
JkNfIiHp9esdv2WOugHKxtF0+m0yClXtfn+hpnt3Ew6Mw4z7n/rbXBrjQEbQ
XR0j0ITSYcn2fR2THBMDwLsHe7vJAVk6+H6TESga5r19T3BuUv4VaDFe8MrG
bjhEgQgED/uG1eXkDwDvEJcZLL2i435j+G4n0Zy4TBVP6Rx63FN3S4Zn+Mwk
QKyXzLFG5BiiId2MIA6HStkPZIjNuAOW3fHXdSHYNK0BSqnsSmAipY2rhkWB
jlwWLmlRlvl9cFoCeM+ymS/6JUWNk2f+diPBfgszP4XPlAMagQmOL2AthwpJ
bvdCPj2dVbZiSYDObUtf+edNdb4yQt02buWis0W080ZkjZSO5+Dyc2QeZsJc
F59uP9sjKNyRBDzwIS+2rc62BfFd9DXFXrPFuDEnMRxhbbnskdiERaTWxVjE
pFOAq3rummI8oeHlTFH1mM7DyMCTRvGO3pwa9mfQmCLyGVewV5ZyZxdcg5D0
MPHEi1AqwhGmgIu5wCkH2czmiH8+JksxidZgmrKjS7A2a8mQfvRKIBb1zb/j
i2pIWyCTGvnDolHZqvkrUGfss8umG/i2gwIwkUHo5ueGMFkBff2wF3qvGPzy
bufQTS7vwJE/kWiW7YUXMS02z3Pb46NStycfW7T45w1Z5lDnu1SYkFy3sU9o
rrx3naxeAi1bPAM5/OUJgpjvtd05vqMgyxFXvrcjUMvNQ/2ihY3E59jV6q8f
7+1Z5ukw3uzf02m6ZTJtJENSUA14e6zCGd9n56rH40iPZWJLV++h1gUXXSdR
s6wCMPOIGC2LY/T5xiD1INdc9a5vTpufMamqy5kXOHqvSD6i3cySt2IHeab8
kt1vsBX3ZlTZ2mbDYi+10jtyOEm2rc0u1b6ld266fXPuS0qgidTjY+qT7nfW
xaiN9A32/1wr0uYJwpIvwmXtkV0cEQQWjYRTjLePcpeCeMqShuC7a7nWKxil
7ZxwMO+zvo2LeGZwnLlmEjAp/JURtvPA7DFkdm4kCJskVcJJY6svzgzxMFbg
YhA2PDiFF5G62E2EfLjdgQ0V+gFavK1Hx2wa8ZD+ghyCwI69n349J9zKeGvn
zIbT+XAPNLp/mqP4OJ4a288DsYHrRWGzrqYSltuekk14WSfyS3jayH7+mRyb
xkB5VTC5WXImXp7GAqNIdKJO2FSyoAbqVROA2Q+OO6ebDTOAU1l1ZwV9YXJv
hjNN1Tot3NAZCwoXH15rmRnfaxJ/M36T9NhghUCNzYzW5cHU1Qg8Mk3HSpjJ
W8fz++h53EQQjhN3gOMafhoTLal89XBm5nBmFNwSnlnXiB7/rgMpOcqANn2U
Gul+XDxwvQhdsljwF54aO+lqGB79MdN1ZTCvzGivbEDxX2x5S38yS+DGqdVb
XWREsglGS/4f0+e603wBfrl2yXwh1A1MULv97DAtr+pDbgzcRSuErkiYsJXz
WiTaFI5N9MKFtR/yFfpo8dbhUXytseyXp8TJHKejb13HVv1Bdbax/xWu9yYg
r+zs2bJj8XcTmgMlHxI6IqqG8VlTwYUxAMmqz15oPAEPIYDs1ral4wjHvzMf
yS5509cCwf3rWexvsW1/NnNBABDzQFy4xrcwLeEwSeeOVjFK9TGZE/k/NK0M
3mKxPPb3J7eo1bx613UhzTa1oNSyI+O+IUNbgOxf0hpDM8tZ2l90Zrw2RJKJ
oJhp/froR2muYl8pViX4NfO49p3Zh5doUFbLMklppW7fzdtjGHRiWNr0v1co
8CnMrlQbrNwaKKON30KDQMYS3Z+NWyU/e+DFy22bJ4znVDnRWXJph3RxIUv7
7B5f+XDm5Yg2mPcECLREyM+2CCXwTXlQKl3DQ8NV8AFq3JtLcb/VVHxs9M0t
2396grn+G4gk3/jWA6zeoiJx4V2LA+tLkif0kqA0JFkLV4s5QKXsUc1WsYcK
zHFv6yJNMPiNLcy/mBAULstV5LmrMZNvGMn63q0GkzKkXpC1NYlmUvplU3Kb
PP+MeSCQC3QBQ6MgTtpB2Zd/5eHrhHWVsEMw9G/aTyULVPUfdos0F0B+o/0Z
f1mS15+RaIGh0gLE7kO1DoatfUi8hKpgtw+chwDLFoiiXIVW/CI0BZFw8x8M
pL4YPOh8zMFI8zc3/ACBBl2kpg9cn7GOW0fN5PZmsf9lQQZPuARnk2moywiZ
Gm1Y57hwRCH1hqXWeM8aulXk92L8Nvz86KPGrqMymx459oN/46EWBqVVuIWQ
U666bFWN5lgE/HuWpdxLqRdh1IEv1vZGmJNuElC8O5y1rH0B/BXURfi9lY67
estGzQtSxdojzQZMropnzR02Bu5erv+0go5OUxKOayLKQYkb7k9l7jV13gng
DjAu16ACpK/UsIrodth/zSWEbeQdUh3xxKjk5MvQE8Kus7xAi8ERJ/9mOBvi
6Xi+6wlTAE+x+AEW5yLX9UoPY3TwdAYqS0/QjgUPMBYnbKUMQh42aNlhl5QA
GsGqgi+HjZxvczarYVdAp938zW5O1ZQkSWd5inPwlq2I5XPmamKjo7zkJeHp
5Zr6D/binXjVidufNspyQxpY4RY9jx8K3577fG6/fConM4vHMajHqk3L4Gzw
uxU8bgXmSrND60b607tRbSo46o756sZybJiVHl3QcCmCBJ9HqgxKkwXil8f6
RdQdlxVCXB2hLOrPR4vYWFlx9w48hPtDfZ+LGVpVWnUfM4TP5tQZVVxu7wUb
eeiikkVSVqXP0O2JdsQ8E+C350eMWzv2iawPax2JbdorsoM7YbocpM/TmVYg
4cZOx2tA3v55lZkYULzD1MkJ1/XA9Rp5FCtSIAF+siX9I4bezNXT42eTu6+X
dVw/N2r69RA2r1Ly+THJ0XBohtPPUowqNq3KK2pqwCvQ6oQOLCOe+hj25T9y
8c0dTHMz5sAHyGjmRjm4cAFezr23zKott8oIF99DlTpIX02keQZtJdpy7kup
nkzIagxxRZ1oDIx06zuaG0sezXvkQo3XYTGzsPfvNXxs8BTmgOorltG8iMyz
RhXBhgZO/aRTUlAXcVUsYEagM5onEQOoTqEW20FPMJcAY8rXsxpF4uJNDSvY
Nn8la8Z41eHTjyvk6DAplteScnT19UjLD4g3GupYM2jvWUcpnE9gwFFDAyxQ
5wvzq0dPePpgIZtRP/5HDJrjAUx2m77ElZ45Jtudb/QN/yFD78TcH71TNNX2
n3EirnUT5eH8zXYvI6ha76pRWzWOKVnWzlp3jceDXmSrkR9frISGESMzJS2h
O616k0jSK+AfPaMozIlw/dQZDRx8U4JV0K+xXT8h1bP8FUHzSZUPWvl80w9i
IuM5hdGKzJ3EQehBKpf0Bs0n9geAc7Kb+IQBtW2xaj9KHzj8c/ON02nIZ64o
CecuvkuIth7pMDZrhBMNGW5tdfvOXgRuAwa12XIZIsFQ1e9u828u1iUC/X1+
t3aJHuvMDmEdOXxk9HT91ru4UeRwe1SeITXd8neSRrmUlyAd0AUwGGAGJ30l
0wglqjCXi/tIYyKPtXHGyxQVgdL3tCpXOlj+0VazLpi/dSTNBWXEUEG4ced4
jIyRfa3OUIrTT0Z8xB/ga8TzKmZbw4faPmNORamp/lTYgaqjygLxZ6jIO/Ou
ODdira3Tp9aS4qAWHnabiFvs5vOs+EujQ456LYNqeO4r6ODrbpMvxwAaXPUi
BZeDzhI/vqCC2qIniD/3y/szSt2MiAZaShLXj6mAk/s2iPC0qNoCjP89Ibtg
NxiA612MxHtJVt4MS5FA4Q1eFs9HZU52rH1RwpnPMlw+BcSsqEl7jYmHjnL0
tTQPgtpuxRcerRnoAE4BWPJ5sOCyc8vgsKdGOye3QgIS60lmrvyWhOwv7Qrn
Trt1UouC7zkFUs+Aek7r/ZASUgOnRGLowJzXxEWHqK5hyZ/tpnl95zIETnDA
GQJ5ZaWrKxYLzic8ZbngaRhivqIQ7+Z/ZlIj7ZeE/pQ3wLxZv51n2eCtfXUJ
8srEpP3Jh7LUdiDN0sOjHb0YnVqzX6aPVB3hetBh/T0puEsZB8z1OdNU8L+j
Zu8t23gRAvxc2r0m+kSo0M0Uak6Z2mFoVfhgIAe8CgHwCHEkCEGL6e41rhfY
ZCgBr2dN7XDm/NWJWZQNft0ZhizC4+hFIZEFAOw31/ifE0TmRy8iXQ0zyQYK
5BKMqQxcNoXnZt7Eim2qZshKW7eGevYRry1ciLy1AGcV9FMcQnZMBfvT1oQL
mHg45dN8I6EzTkzZlCXgPeEtUy5SQBonySOxcVhF3F9ScxGKjm5mUEL5uBk/
OM2Q5WkAWPUEXIRFhhEk6XinihniqpPv691HeiN/QWIchBdYsv7Xq/tIYR0w
Vu6t8Q5U76yMjVdZMhs5mJL3Z8Nf3OPlybEMEhDP9EA9jgtWW0c6Rua7Xmhw
QcLq3kXDR/Zvm6dIyxqjBLm5qyC8XORJgAPxrHuwVRPUByx7owI0qiLCOZNo
/SJy2yyraieh3RtuF71flhgbyN9riCBkGW44zfICwqfYOP69V0s3/p+yk47O
GSG5OjOJKedMGCNmAUaIkcGFNrSdRElL53Yld8mcX5PMtOu3cpWFS/beZKSd
S9xuTrBA1mq/Ra3gR3w4INq/UxswXwYOstKneJukXIDl5l9LdySEBQVidl6w
wcOlnpRguovB14oxCZbNn08IfFBP1JkLO0BQgH+ToBtVjOB6qc41n9QOErnF
Hswtq96ykR0kthG6gNw7Enw1cKqTfBidBk/IaVG/b8yrLipGm+7+cEKBJCqe
fvtap5gyN7o97UQRU8CQCA2vIGC+HNOYxVKZSoWomjCmQNf4SuT2g4lo4BrX
mDEaS5D0U6RTexuZod/R+5jV1Griqq5aDJYu5eV3jh1I3oxKbWlFgovkKOwM
1daRhXF1yIstRSVVwKikpaKdokzAszjdUTYV82F8SlQk1PUh7JdSQh1lgQTr
OiCdgB40xJSoW2jqEZGV+brR4O5Hj1+AJPR6VHBi9O6Qnfz7I+Eze25UcD5i
MENDe/IvNCVs+fa1lAe9cyvTmbWvcW7bvqHY82kc/trebC41SRu21MJIsKtC
lMVr6aCs9+N2B+sfaPOSku8CSiPjp7GEHCaGI2zchhvUw3TtFWqkgagHGnz/
7wrTU41x0xdG4WwhllALGhnE8L7z2bOAfKzO+gOJrSL1xD2nQ9Ah2V1aQsCB
xQi8++BdkUnr9O01pfgTEAnHgwjzWy16q2mz2G2B+HTd7QTILJNB6KgJD1FU
l3GWRwKeIROj76VxmoZ5inR+2bNaGsBO+HxLsbhgS9qJdqJ0Ga8niB8oKfYX
qJa+VzfBXzrDw3rVSjeyTtE0dbt+mRWkrhn06kWsV3suw7XLx6+Pap7Aszpq
BlSu6RYSmNV5FuBHU+/IuN9hPjTTPxpNRX8wi8lhGbHBLCIRQItmcLav/oK6
g14qhy9MtS1CT64gqqQ9CZDcQeBhYIpzgcAiN6YImeBQqQ+9AeJbaYGVT63U
K3ruER4zQ3NmC9TKvvXUmG7FlWidMa40rAid0swPWjBSeAXNW/Fx45CCpXMK
6N3xznY5rl0/4iJPN1eu4yrf0x+vQNh+8X2ECpJz/fg8vN3XE+J3Y0VVSAtx
VyTch6iGW5T5N6SI/DetvaZ6wHoOqk++5BWs4U6vxhSowz2pYHYCWvw7jf2m
c6cFRw2VIb9LzjI7pswIMDNj1K9hU/ppgYqXwjTy2ARZN53X3v3pcEZ7Q2ke
G0/1sc9aosr2Us/SGoYef7NDtf8RhQXyweO92/dqOqqEoAbp4m6UwFPF0ggl
5924WQ/8XRiXQX2gUqLPs0t+2UmPSIe0DCRSetJVw9UtrgsoNbHuMNUJPjfB
ovG1rHThlc08HHzS02pfntRDG2J8VE0ywUEJiwJwimo/WQhIJLX84qXfcfjA
Lxadrf6cpjGMj6QQWDTbZxl9LOV37/3NDn3RjeMBqS6M7ITBTpREhlzqCOue
eioaZ8iHagG7ak4jwIUPw4MOsEYgUerorjWt69Dpw+YWu/ldlQutvuhY/diq
5igwnyQ0argIRYAjDgOXtf3kdUOFo3awR5Bsu1XjKKgEgO0GhTKYcA9537s4
1NHbra0l8fimr9ZaYQH8+z/AW7LkpEk92sQuclnAP21I2DxvKPgA5hBeGhUe
gMF7cy3+4+pvglFkOe008fUwyeuimtdUiXPwuFwFoX7IKO0k6iGmnIR1G0EA
Dj0kbCHU7v8G0cKd/9Ru4FTGCcvkY4x8/pD0QCvAFTtjgp8kgkk0N1ga9254
d/Ko7f8Fnfqbd5raV4k5+2U93LF4B2jOkbgrzjZ89ivxFurmq2szPf42RZq1
FYdgohxeg+gSjLy1kiK1+7ZZmcxALLXHqbZx7Ty9hgvOU3At99NvawtyGunq
HhzdaMO+oHH/cp5tOXUsCfDNJSdih3uHl0U7hQ/gqUcawFNpI15djJeOIP15
Z79+/6pj+d8LsnwpCq4dJUe0UA3UYvwqH2i2fEtkePpMIDZCI+cnFhnL4xJo
h3LN3FEQQr0Fx/LGQhemtvDpNEEHF6RX9V6/swoUZ2lh2D4Ye8ry/ZIcX4+A
e++9ugnzsRillNi0Krqp8geymcQCkAyUABfg1NniIx/L2JxH0vQ7UOdvPyrZ
DbIaTgpX2Bb1WbdPb91zxgmgjJ5qUcTvjAwmtiP1kgyIwxs2/4ivfg25xYI/
puC2m0cy3mwemnpxMTqOa3n0Lt/lQYtYXYxCGDhTnUIHg9Pl4lIAksKXcGbP
NfdvDsBJ0bvf+aQyCik2PIHaVGbL86xernaiy95OLQB4EfVi02o8ALNI4aR7
PQMMS460Jfbx1D8Dy3XuU5gNaYl+QAfemabsMcFD3BqcXqdKhYUpJ8Wk6kqo
byRVRLm4knfgrlA7XcI43YtJyVJLabG5quN1SEkALwbWyGQ7cJvVoVCqjm21
OFS9nBBeFs5NOTMNTgcrcBYNNXQIGV9L+1hNOGnYU5VORbEbOiAK9mIIrLFD
mD+nMu+B5btnpHpZ5h0rlKREor/GHSVVtPpOA5PEjdzFDXDNzg5hEQ4qK6My
61uFFYNiW/dKO5WA6b8q3bnilq9adRejAQdxOyIJUjXkp5C2NzUeBFJ3wOPO
4X7ynaRTN9fuBMX/lQWqtmSKSFxknWuZOfuiqErOhx573E8weQpkR01yBMfv
gh7Repf+ALdBrIS2uMfbanmUEspkeQfAoR5WCZO2zXJLyE5mlFgz9FCG55TU
rtqKTzX42QjxnK9vZ0x7lQNIsN0K+o7jPeZwh79/w5IcGo7aHDoZQVqE80oU
quAILQWz0B2z/esAfVj1tAOgQTWKTRo0rJD/5conz45c5PSnjgZnLhX5CsWb
ZcE3T1DGvyKkji+bvmh1hCi4DR1ATPwHhTuc+TwDFwpdNTExrbzjVOOO6+pt
V4MVPUoGjQf9inliDSLO/JLHhGEehICOspiiJiF57Q0cnboqhWrQOdCHz+XI
dRWV+Z4+YLrrJtntNQUqCSa8MJ3JBt0GiFn8AnKOShdmrXmlMweiJlAHDSFE
r5vN93SOHb+mNV7A1Ry8Y8wyitk1eiONTOovKe2IYTyvIsYN3Zu0bgzM2eEY
hWhZm1GrX2vmDCghzyoutdkpmakLT/+FE9JyEd+AtpdbTSspIBlv+jBD3cjN
/vbgYZZmQP7S5ULBCCOgJ5gaHpcdJ6ghkrUcsoV2jBYOWAk9zvNMAmS25QM2
hbZlMl7fra1O2f5C18qLX7YmF1hFhjw0ZsVEnOwggafvwhqWUV879r/+584l
mkWIWdzuT4EA0LqIKUhL6fB8l3pG0IYRWPY26zwqJgCmzM27pqrW8k7iRJjM
03Bgn6UdntAaHWiHOwtLMYieaEwPYSxInwKOWPlqjv33FxHHP6b2csV2zgTd
b3FL9HPnuWGuZLklIgKQ6gG50y/aM/quMuIJ++FyeELCr5xo4+yZmq/vg1NA
VQaK5YPp/lZ94X3g1kxjNsCcg5MIjgTCqW7l8ez/vCUaDYP6KWUFOJXpsCrN
ibNUVofY+H9QiH1IRK9crU5psZvx9qEZ8XapzyuYR9MdIbB3xHj8au22HiLd
fcMwozvPSr9intubmTZlMwUPVyD/E8HMCxUqvW/xlz5tjOlL8637FA9RdWSP
aUNOnBWzTaFNyxQpn3yL74ZKXeGyUZ/CTBghNFR81G790K3i5l4phjQq9Kr3
RiQJCh9gDwj5/JylY4nb8zebj3OXc5R1YEyOsVJcNroygbwFOlrphBZcFXp6
3v1dr6cuVqC2+KKOpbLwlp8hzGeynlUcIoC7Aww/HqplNfMldxPHV34NbIMT
8k9GgN6jUrHe0nTu9eakZBbE9T+/K660N24VN1zP7FQx0OKHTmN6CXrgQYmy
gmMU/X1TpCQlEiuex26o5rSaoSXe3UWGbzo+gOTXq1CdDXfrO8SeFdGaooCu
1oVngGy/0nvuj+ey30vZESdIAU4AVAKOjX+xAdKanXdC6gO/IyPuWbcGn2wE
2RxCMF/yDr8GtfwShzVNP4qlbeAsL24KTGGxoLZoXTPPbgrtZfCMDqq0UuyZ
+OAeKxUbHc6vTbgwX+1fFHa1pfQeYUyxfcl8asV2PL9oUhmHH7Tw3MEQEHr/
fvc6RqApy4fzgCrhkFBt8o7DbuU/2K0UnIjqpXye5OXta8IwF3FPqbk8ZMnE
x0eSGX1XibClpq3sgYzKda1h/jm5BoLiNZQmyaH0BNl2BMwjdQEp6p19lErz
SGYUxdLJ6FfBosrSU5IIhHgW4d2dxNamsvIP4ge333MfRcTxBbE3PEE7fPBk
GX3HX53HDjr+fT2T6EOG64dFKIbEHuxt9Hmi4KnHOSk7lfXhZfUw3gvLYTVa
toZGJb7N/nh7WKqaF/DuRj4UqpB14mNlbFxlr5Ta06ETWUKu5tIa4otHCzOR
D/AyYIm8QjNWA7WajVsKH5wx9B8VJFClHGAHFaBPj2PbSqPNPjc4+jZPSkts
w11dodDohG2YrAAktR0MzojbnZRNU//HJaaVRS+G7vBNeT/TWo4709drsBuL
6AbOZlqhylfX+0a+Jv2WIu783pcWWlTFYoXR7q7y+ZL1kAD70NCBqZEg6adx
DckLeSnRYf7DKmvNRJTkxVft9Nn1mU8VoHxrKD1oS7jX/UHyDJObi+vE7WKg
Shl1hmUBQOFSab3DaN284NQroX08K6cDcC3mWEaZUP2viCNtS1kjCAyS34E8
Ldu8P47pQapXpiUA1IMfd+/zF/XyqguD5sL0XoQGLyQNOfkBcBQZXEaUo1C2
ZtEgGtbtf5xpRm3IlnfyOlDCfw4VB4Yols8SfFAj02NsnvlnJ7ecT/71jCZY
6z8fac2uY3jE4oOpsWEPShU8kiwCZdOngWnJefWed2F6IEF21qGyBC/P+NVn
dRz9xvH7KrL/FvxvgWB0w2E5qzatUTZb2UIipBcwVZii/k8TEcdj3aUVYBfc
Ar0N0awyJQwIEnA9GcW65NXTJ0aIUgmfd2bJt0JRHUCTXekGrBpolOD7maid
4CocG231v8EGoq2puUB0yp52wW+SividuTWSA0crcYzbutMtCxwbWPS3Jy1y
bxvM86iP7rknvsmNzy1TATqqKkTQfxdAdnJGFt4AUIaLCrnOAZfI3SUdB0H6
qssNmLmbzHstUgu9kuc1vMhy8p/YeIBZjhrt5YG+64G3IwIZhugeoXAYOmRS
yvBRcobCGLTIaQco+T4l1hRlGjtyDjBkRk2lFpDr+pWJGJ59XPw5TiWOQSN4
V0vn/QeIut+vdXHTEgc5OEIfDWPwRWjVgl8rW8rPfgAiF63A9Kq+Xydq3Kxs
EyxY88xtgnfwdV8+VCR1LbP/JxZ2DnEB+UhuEiABsYshmyfgN93MTXmevYx8
LG+l37+1cVSlbMgQwtej0azIbLTD7B3Bx5H6Ir+983Sf8z0REGsKkKQ+5WBY
kDIMbRWuLhFnyEpsXKDZjaXE7nqxxGcOVngGRLy/oaW7IQ/+rBmEdO6wil//
xA06bGmoQ78R61yp/Fa7xwJll9JdIR7m4+WfWbEvRQSYG4PX0hFr2Ff7Ouat
gJg8NIWK2E786nZlii9HpoB3e2l5mxNwvmvZckVKC7nHW+GhSbSaR0SORecF
tEqQjxbXoM5ZN/vrM7Pu6V4E7ju6Afe2a2RgyQ3sQJhY0Edbz10XEvF40crE
5YrGayg2qtbBhB/usuL3naHt2LJAxhRNyVjpbG+6QBlb7oSIUiaRnRbSOqzm
tuelP0uSiPkKCo4N2jqDHpOSVB5IFpRth//H1KiwV3WBMyJsm7DZ7j5NEej2
AcVYCNPdvBpvrGwxDsXUnbYf6LfyzYiGALbK1L45bdvuSUQb+tfxfT0sVel4
srz7AmI1nS0WaPjwIilLMo3qPb1LfCJ0G5hMeCz5rS9MdXLDeT1u3UhjQWke
7k7SQ6yn1nQbgkMM3wssFf/SgZsRAFvUtJ8pkwGG8USRccpNZs63rAftG8zR
JXcepbjbLOY8rUes03xLp57241+NsgpKJaLe4lhHgwJDzfzZm2bs2dQjsGgo
FUX2j2I5pTmZiyjfX+TGB0QDxwya7om3TdLotUT47okTsnGAjHpuvfCvoZ8c
YflgGrfLCAg8IMNTqNbprDUGtpUzAUIr1Qo9ExrjIf+xe43feVSZaOh/iEol
Jqt2YMiIWx4dydePF4rRPwwPB9UXqjHsgyHh2jG9LEvHTq7zbVoF9MBnsix+
DHMuoH2ywPcXoXLdp46Vkh8yY8WzHXbxus0NW3UHiLPbqW8BOELE2sahP2pc
vDs6T7PnY+TCJZXTmaSnZY4dYEduEkuaLbbwIE0KJmowbRs2/Z7my2FFTRUA
8AakyX29TDeio6aWuIgs0ir2bQbE/Q6qyo/KAxqVjWOVcmrmhE3p0EdtdpcN
dZs7gZUasUSoe7TLeZqe7fRTkXkiAnRbMAO/XScxSuJFpkkMP+NW9viPKC0p
DUjSoUOAzHZtr0Ct3r3oCrojaHi7PTs/aZzolwKbf1M3jOY5fl3XU1IA9Uk6
3nPdOsS4btJSd6nSFKVPprftP5gGdAhNlnotQufnuhoPThfHK5ibDQTrhCfa
uEH0mkMkNJ74CvJyC/+WnzJwWGienvbjafkaLHykK/1+DW5EKaSU03TEvj/l
bFATmLxH8uGBy1tJrQJ4WF+Ibz5WVUKxOLpEA53510vWdN10PWJEEsI877Gp
itVglaCAR+KHmIkBANkC8YDDGbyzq1MPeunTl91rNun6cBXKZUPfr+o3tkmc
FzcWV/uGpUgIpb+LBHEvUKz7JstHy+3NalPap+t31fGUIv9GihOFBEcKEW4Z
fYnlEePdGG2SLwEPSEME4kkSaCPojTem/wU0ZEFvl2q+EvwmhcnHkjJM1cY6
U1LviPlCJxYiwIrQUcKpqtmp3zH0+HKw8BIgDE7Jeu2QZAauLmCCccSoqatT
p0omUMWvCYLWtkk77GJUfH3KpLyOVlMefxEUoqQVkyy0QgNeyogQsukspV70
qS+8Q7IDcLeyqNztetYhUP9Anm770pc3nsnFGbUsIM7iUK+U5Ens0t1YGrlq
j5Tu/QRJhH7jroY+Xv0rPKq8iQRgHbSu8sV8JNd8rIMCs69RsPrezaMVF1Zj
wQgAoRv9ajnS7yZpWxo5c1flf6sbDfZYHsfs6oRsVH8CTNPsSX+c4mCNiN8n
APNPklyNBTLukSHpsIzDPceUBtYL/CCGHAJh2njD7NsuqHUuGDTZE490W19p
9tSbApEmpMFf2Q8VnZmf361iDkLyn6WuxajTSvQiD0sp9+myz2dcH3IOcC9M
Jge9w259kQOjcOD8oy33ENIKxRiPRSSA8Msnuu6dcL9wEMnEOiHaL3wSfOjY
ok5qyAloV8AI7CaeZ2t++2RA0UstLgQ+zKQiJKewKb3NCDoQAQHC8SxQyApD
5O+8bWqYkM0+3R6xOUoDZYlYivpnyptsajLR6YBI8J6N7tFwHbdCJSQbcCyL
oxOPR9YUrB2rYCsclCbOdKm8TTYNhe2iEtBHSMCgctEw6XYTsRzl2DdJFDAN
WPRfBwpfEWhjxINljQmaE7gmvDUyut61QAS0putzQWImYMI2GDPO66JJSIh4
wPvNydXtcFEc0IMQDZqWqlwZ9hvd0K2xHAoedW/TCArxeoPIN23i6oAyaMG4
6QyDO99B6psHx2iftXnHXtupvMtBNWirvS6kblN+koLLHVbJtc8ofRyia7nO
dnyms/6MDCtzpbKM7Ggu1mTzkNdM4kQiu6/q51zbHF9wj2VOPilaxFcIczM1
K/ZTqMqBkVaX7pk3n9JkRvK4s2vmUOsTCjfE3NpoPObrDJ03L55LxKSi2K5E
Wl6cRgPh2SeCaz3/jH0EUKx0vOhV0MV9By0ZB3iASYhLvKLLsQgf6BJ4Cefm
W5RAXPTLP1lKiufEfFE3iyjnT/K2YAwAgQNb6F9zE69cDdY+cFxsTpmvw8WW
nDEnwKFrm5paH+gMysqlsdfgoS3sYsFB7VeFwVc1yi3PUNE2j2hCGHh1THU+
gAzadIdB9MIZkEw1ceOjCNJL/feFz/hGlhvM2HTRh3InTN4WmMrzs4AXBZ0d
ETWRVMl0cfazHQqmg7cyHAbEm3OTqpN5lRh9P229GnQrMp7owTVxbcBEthPl
jfzDivDZe0kz9brR/Vmcu92MtOxfT3ArUMNz3lHfrDAVbUvwybJf+FUvkYGB
VyivDmUEGXDIVdMlWkfgZzD25PpobNv34x1/0s7rdvHOjx9XiNEO9A6d1EDN
J7I+kUWTutpUa+YGxC8SYcep9n9F7zTy37cDnA1yyLR0Ajzm9aykwuoKnI80
TaUAPGYHwgdbvcHHdgvCdEeVieMWyMYzSn2x0Oy2dDjE0NJoIt9j4GOJYLoT
O0fdjabPyVWQbkwcYs4pNn1acWxTcSjr2IwYoiU1m2BgTSqtY5G+9UIMlSjZ
179Hfrkd4NersHtAQBkG/dpA+VnnKvBDy8u7B0Bxr2ir8pewXLOsDAOgwCvn
LMGR6axLCL3tyTdfhr9jsXxwj2CdW7abBG8uF1yBBj84/egeQP9KmHbyKQuz
7TYV52LUhLaYnkAW8RBICIvMDaYyRkgdnrjtWN3i+Vn9/yNKQDc+9D9Ynptl
t4Plc6PehIQ57eeCSh37eofXjWISXVDSI2P7uPxT4HLId5aarrmlTARNhUN+
8hwiWxwrbpCogYzwi4X3MmFA2SM5Z0If86ODolOPAHcVjbfc5jIAvXeQOHNd
faxOfte8ifosJ2KI7Qop3VslEBfzoW66bdZUySda2aYw8D/ITKSMgoXQetq5
BPgEVmf5TJcUdC3hzRBoBRjpjXXqf/j1TF8KSCTmUzjHP4ojFg1KitDEfrqJ
Pf+k1hJMlCF2AZUpzD6e0BPJa6+rWvpKCWz+pYWA43Tb490bJ869tL23sLI7
bV2l4Z5TGAykYP7+fG+hF50K6HYEvC3ZYuOTNWgVZ0fB3eyhT9WCD7SMGUo7
QXhnU+8x4stYA6/JRUSlCeT7Kr6LJZ2lU/TekhL5FN28MO2t+tYhazdNjhZX
Qs2Rn/LJE2FwTUnqI64+DWyCkzF6dbnI1wYNaIaurHw0fuzTxdlFN1OhFusC
pMCcZ4xKRQIGvv+iQc/rP6JNxHSdhLMIaFGpUQZjOuPj1KB3euxlTsGHfPyz
sGpPGKBcwBVdDHBDdDK5anCfAPZbN4Oo5dEzhzuUyWrDny50higRLJuGN9HF
y12nG2FkeAySO8r4nTfZ7+nc0L/1B17+6j+nFaORCgJyLVar5USABLOC0io1
ae2poxJ6wPN6p5qwx9MwR1nYvzPTVgmX2HX8+vbmaMnq+Zti5dPXe//ucz0F
mneCulfiHTQjwaibzTdz8QF/QM6zaVubggwhr3NUKWEVmjECHF514B5fmfEM
rHe6dno6+GP4W24mAoYiedkai8PdSmNI1RSM45nDFztNKtKLvEf8CUXnl3ED
RIs/2FI9ykdBz5LthPJXEUoSExoj/owdxXy+xHnUuGdEFsJEDA42I2xeB0PS
p4dBn7bhF2dn041XnrGm674W48BGaHU2tlm+qNviFFf/LyxFMeOWDe6hZ7YT
EVNYrq7VuWsKIOzYDun8kecr91MGTWu//eRjfhwrLZCjtHZLD5tbprZiy3MS
zyKr70/h7D0HItN7e8hm0xDb1HwXaZKgLpSop3vXTiFLNHkST5QVwd3eV8UT
6WYJDqxDQnX3E3hfAWrNOn3ELxZYioITQq8wMIoY/NrdPGXU+HnwOHA691W0
T0T39gkBBN2XOf3yhG+0RKCI/XOfA3KO4LAIjHsgPUDuVbzghJc+csjql/Pw
mDLHdUq0O8GEWZQjXF/9a3/+9VNsCXI0B36E63a2N6X2+xLvksEg3XTROO4a
anzMN/J69Cy1Yc30K82O5gOr/igwkNg8Ppj2+73tLe3LwJUOXPuO0RmBXtbV
EL5wIdlUt60KBx6O5rnCu41cvChLA85oEIZ6urXBjJfA9VY/931E7oOfX9Gs
BdiinN/2/JoXzijt+b/EuLsafAuOjCvsOXdUymWcac0L6/jgMwu7TVIQ5v6U
q3ciVmLiXt4tZEB5UHAFWwFkn47CB4r+/LkugB1TlDSgFndE1mRgC+hkmFpV
/39YfKx2IyZ35GG7LNp7DBomTDXgK0e6s7zD2jiWjjquYhLTBntaz52hwASl
09p3mvqILV/N1VwUatmLnyVWWPubQ34smSl42aoksX0T6QxI4w2luCnF4X78
VxiYP8rmXziIWmEfe9tVPpz0lUbtQtkoCsOqHpG2feJPe9x/vglZbszlmBv5
adR6Lm9I02MoDiWu8YHFdYxwgSc1bD0P7pG0s2A7SM+WiciwAfM1/mTDOn6A
Z2c74OscqPji2YWRFpNbeEK1Z9KeQK0m/oRs0WxRH31ZBEqdmVb+HNfUHL2o
i/IEJ3ngGejXldq9EasjwyUwZEjMG/Qn81ugJW39YVsHhJ287W2I0TUYF2Mk
sb+QDAadUkFdDT0Twjnmgd3KX379tVfCWcYdUh6c9cOIGo6PZGMRfPihPxgr
wuhdX1C4NOwAFa6wHD7JrIaJYGnbLvT/YcImGcOTgtl62ohShmUtWtjYxpVu
YASKQzN1QoVe9LtnOD8c87cV48imHp2b8dm+w1xF75YqYtYj/twXDbi/dI95
jZkCpBsnadHi7sNjYPU9vvx70ixzo8MFTSXKKsaQhDZiiJBkwZne+HhNUP5B
Ua6VJx6Yzqw35PbcrG9PXoq4aZmE6EuTEByRPdDElaBh5vKPMAJF9BnCJuwK
v/jtVekX1niOF5z1OVzp1CQcrxV4HZY9+6+uYwM2YAcnERD0Jsh0FTe7obBK
JqbnvLBxtyLOWH9IpncYW5NPEHE4n2BCNHoA9VYdKMLby6owoCnX2IkBt3uz
/oCHkw/rO4LY/ECrOl7AGnPz+tuPbajv5yTwTb1VU0VjL6TA71v/nnKSXspZ
Hhv8OTmaHkNUBNw4JOqUpy8kWZU/KPVDE7UigccVhfnCyLlov29kD1nhsTmD
yZBRQNj7AZWZgGDFxEzqQWX5IYf2zKe4U2LAgejXfMiGQC8MJz2mTPsAu2w8
Us7ov07+feqadi9D0ylJGR3QzcCVf+Qci5UZ2qH2DfVh3jDpn9d+zddzxo8N
Gk9TKAzBSNmXwIdkyVBSQ2SIkc/5KYQk/+lAVcml2kN/OTR547tVXnPimxaD
j9NuSt+Jqdqs8mQHhjfeeeU1XKDa6gYKMLADzWuwFMG1WHRs7k6BFceX2SKM
2/bb1OD/I8SA5btu+4/z6HdO9BTxe+gHDnJmvZm66VctB27eZVSYMejWx5LC
AWf3bKA2QmNIHpdlvIif/JmGL12Glhekr/XJMDBoxuEFw7giJZrzItA0rd7P
4xH4nZMcr+jE176oaJAJ0u9DKHXhB3iUUW23OGvnFmm0UoN5O2q5iihUc8vG
xhZZ+eRoATLr2oXROtXy+vCqYQKS/xpKzmZyR8FFqiih/lVT3e06urEwVy05
DAof8n5reP/KDqmCiq01hOzKxLBFW1r6VyG47LEagQRq9Mfi2hPK3KX14z83
I2+XCdbX9J2sKMeGxcW61H0ECjq8Hrz245oU4JkHAM/5MG3bEuk9zz5r6/rK
LxeOFPneULjN1IuqjSLO1fKQFFF1rYoXSweCB4RcYAAUllNqbYR2gG9zqs6r
AOWXMY8BDIjZ0yht/TO7VwXxPXWBSJKHwnXpOzb/v3m0/K7ouCYc6gX9N2+W
xURvoy+mDQTEBVva98lUySY+hvIpdLYxVEOP3BAcb3M1vvE7Kkml29tsqI2K
FGVBVTQjgxMtnwnBUhah8ZFrdQdbdvf37/FDfMLPrL/2qj7FijarFXK2h+BZ
2Jovjt/6/Wj7XyOhDZePSFF4UCWiWooRaBFU0MbgM07+tkdF0eNqDCpxAmqX
hr9Wx2Hfy0PgKh5YwfzrBqzqswRwFkhwmV293OMXUJt2f/p6iB/YFno/zB1F
mEJzU3BX60qrPkhGGeenTgHfOLty3JhBQTFnkaC/OQ1OmxD015zRrV5jKEcR
huN3wKagemJ/EaiHoDt7InGyZGEoqBVtsc2Mvz7gCPcuFgWcV/6U5e7cp4Uw
Od/YEKUwdXyaEu5lee1YOXTof8CnaESSUSd63GM7QHAkvnym31iW7tvn6QYG
MKJBPqZzWYDxHXgxPuIEijRm1fiogsjcxwAJjMPYdOeskuKwIiFXgFeZPUf9
GD2bcfWDHiezjBZMLpCJPm+UsC25x+k+XbvzhFSDCGEouu46najNLiEki/t9
QpZgeZ6wQLmqQFWD6qQUfpNIHJwqqM89BgbHegUwLlQpruy/rHedunGVFayQ
9/ok9cDLBrUbEAhvuwz6Dxmc1CtJNLREymLBh+jSxmDZhYdZxh3GrLFKWZm9
B4j2tW7rvAEWnETFeSB0JATEf9vC6bWh1JyVrY3h0G3v7sIBOc7w1GCVVJXj
FZhb3A6w65xoOOWDFLELlOTzVeTh0roITppOvpGhT9F1Bou2Mxyd72xbN8O2
NrUX4K0L+x0Ps4OJK7C3iSK02WKDAi1W2+P+q1rpQ1mhGBSO2zLBua+W2sqt
n0Uc7Lu3rMR5Qin8qxPHSOzno24iHf8wVGMOlNZP2eegEVoLtl5EjOaVEqbk
jcGNhQVERtLlQOaBvS3mbjmyVme9YL8z3363BALhnFyAjrnA5vak+L/w1M/P
FCb+5qw9NPN+/MbF8W4FR/PIGCFXFczzWU66BhL0sRFue91gTu8q2MrpUEEL
E3zdRN9NFTfrdbl/gRODvlks0hB+qHR81nC8+LpvlBQ8vUjTrYcrbnkCaeVx
1l01aDjtcypOUO7m7110tHsT0h7X9bKk2kimAYS54PXETYc5zdUleRzIMVok
hPALlkaajMM+vvs5FwnEwXLZXANQ3x+3/FRX/Xm67RYA/FPy3iR3d5OFbS1a
E89vO4YDRifSZMkaZ8AhTRqKW3qcMjSiIZCSfPK7u5E47ypHzp0ZZIVSFTmN
ILXDj0JODzXc7dYHe4v2Pl3IdC55Pv2MKXJuO1VMmobwSQO3QmRgSdbG+9MQ
fqmpDs0ZfSfMueWRKeChag72lkTGnVp1zevi8idm0umRdAQRaMUis3pftENh
nEurbEBjA6Ovks9bj7AjlQjZ0llA1V96CAUp6gHlELjE1E0iu1+cavjDnh8u
0u0c2U1ZEu8C9iMF06MBS6Swpev5l2ywero5MsUjXeTJqBSkO1cSWsumDjGD
luYTXPbTPGRE0HzclXJMe1jz1GkSLm68YiBnJczeb02v0m48wgoQJQQY32RI
+1mdFRw6PFtHDBAH5IgBXedovQm24immAL51D3YSv7ogLPq6AKEMB6XUthXd
foQm6Q/+Df92ivGa/uH70HWFbgunsWjPhU/ff9BiwRKwI7uuv0xMCySfudZi
xqp77sd2xo03BkDAtM2sRMIo9dlpdJixNuwX9Q0/1ee8zUz/8Kavfp38Xuzr
9fK3fNJJ8osOeJYB7Cy8h68g9hr3uO0cAUZoY29z+nToVSY2Yx9v3yll7wAJ
4tE5BizL/wDS9yuCCEY07zmc0lI2v9ig+y9Haq4y9Z+gL//s6PGYrRf11BXS
wxVXMxN3XuRNAZBTdWRoL6HOuPzNAfZ1fO0+ODzo4EXbOLgxk4wjW7fJVIjk
SrOAOCUjElouMD5wK1Q8R6RI8ghsXS57RsFfS14apPSJubJXAzsVpht5M0fD
JzKDnYp4btduYbBxRZ0074QjBpo2cPVTFORxpYP2EUfOVWidyVjjqzrb81wd
6TZACWM3EMux6/wqHJ3e9/uXQdBBLaA2W07HaxwmNoxYaMElrZbZdGDgwARL
EIKCLMuMRy4aVumBed+CFw6Con77HrHP8BI/5NfdRTUxtTQRLQR34hIvJFqB
PmnwKlxXNkiZxBtTF2vqj3/8Dk6kmp5EDQB1fIueUqRYCxS5HVwI03kzbWUH
GEBw229gtDYgHcexCf5MsobEoa+MZcgNhDWi5xD9djr/U1jGgySgnWuGDMac
P1LSskWl0ecnyluVujgCBZxX1TVEY1sfVoSPYRVaQrQqGET6ClWCaTayxLFI
c4rGzaCfgYttzqh1eBejl8louzydJvzIc1q4zs51v460LY2v7vV9PS9kVze0
ouSVeSz8CwzKGsTk2m4TaWe5aedCagmaIFo7njK16SXGjafEIjO6yn0h19ph
P6G7a1khrxM3X2/JOEwIjAooGYYGcKFMfvPTK1uo9hPEElRLpWv0bUo8S1Gf
Jsl9n1nsZNwFSrYy7WhsWNoGoNBpKJqP3Ifu2vLzl3TAAyvk+jyuaMnut5d1
rcqBCqTaCApMejrsDWfY6LJNpGWqZufu0Z5js4WSlYDuN7mcavKiREW7C+ga
7HkWCgCllsJgZQJ9dJ+q8atIvDZNf6NQ3I6v5mWrDUEZkCQtT9axyn/4GfLP
mGAhWWzbiSXHqq8o2Y2BBMJkIlvXtLn67mtPkU0TmU/oGbVMtfcqKzv+8S/e
KpGXo/SOORRfi3DXo11mOLA7QPsLqDJ1Cy3w0R6F42RTBdnCzWw+vzt5bHZo
at43JvvEntqz3JLe6TUzicNdaLp05hMZ+W8txMxyQn4/TRBdT7/eyRLeWbdf
YiENRhXR4TkTqFtm55kKA6Pm/EmyolScpch/ug/xETFaJs6UeSJgFOFWH9+m
w52tIOeCYZyVhgaT0PvmDYkFVFEvn7/xEO9VtArVqq5cntWP6jX8Esdrs40O
IQj5CwA/S6hUWVS294D0+UgmsW11JCknHRr36LjA/HmpuosaRBaVQ2yn299z
v2ZfcsKmMCFtWKBZpMUOmX9VjvwEVuEq+PvPxBUAaLKdVF5SrlKqAKpPTYkJ
h2vUvs/sUmVqJDvwMAAeuGYrP0s6UJzt/NSMZaMZE18CSDIUKvoNHCfbq7CS
cltUFARBlp6SxnatTjnKJcQaK9eyAVm3CfkM2iNbVtbCaBgSIEapDwCQXuMN
Pw9Xb3Wn9KsK52mcz6HFvmfLEmeJ4P1fgF4vxDHoQQD5jvKJMfKsDa6xrJAN
9O3oRFc+kq/sWVcG3D5klsH5Jn5B3SJxqbkme+KqcJumMSfj6WIiykluHEyH
OH5LQnFIIKdSw/Ypd7hnqa9+jF1OOWnwTvkLlgGrxlcW1Aal7MeuLP8FXkwd
qmt/VGXbX1XYcvSwLjUX+MyoV+rG2n1G7AbZbGFR4q5yvR3MYUVCIcp/I7KF
IfktF4bpxCB5TvDmArZwJR4UaFEvsDv4osHo/3RUuln05mpA4orNdCbSOhgs
S2JF77syffHMuWDYOoFW8RRpy+/SPhzrNMOTXWdQqvgKGdwjiDdwEVVyZ0We
JUpGPBrSpPluEP8+gimEq7y3x+Cus/iVUFkX32vPEZhFUfGmsgdVNdSp+2le
Ts2UvQ88vc5LIPbmRt7eHAL3oCM4STQWlehn2NEZy4v+ZaszE19biEmyIh0V
dW5b/+/jpQWjvemxW/j7XX1PVSiC9qoxEDAdMbujx7SNgVtFAZN81p0znCte
5t636l7Iu78sNGHntmOHtOCAyOmr56fqSP+rd6xETvguIiEqCnh3cxMlkhfF
upnJsNqRTmbpTE0+2U0a/5lRRZnBk+OkZibchKVJtEpm4W4LGqgXSfOCERja
B87uZuo/CHoYJGQ/eMpUsWA+4uEIZJ37Xv+md6vLuRoGc+mlimrc9lwrS2Ew
/84p6NA2yArhXHau5T/wsbff+dLswoysgBTP3PskM7tq1U1xIT4EpTxTBl12
3uxGUTFyu+XwRd+DO/+lo1FiHZ5V/xByq3KEMd2UtFtc9fCkWvQps7nSAO94
EmQX/rB/VeecgKclqaTp46/F4ukdl4kzPvxfJRU6YM99H5CNO/MHkUDC9ogT
khfA1rntU1SoSb6kZOD4upchvUOx/XGy2yQWEXAWSJOjtPyCkprLNZzppy5a
od+XUjlZhkA6OLYZElOiHMeyL17u4hOy580A1+y11GTHJSBikJ5C0lU9sU7C
Hm935m/o96OYl2NBqzL+CRbf5Giddm/g+XSY0D+MX6phPXmE5Ezv54BQmetu
55iO4I1fgSg6G66ZT5pTp3BOv4Vl/79qj7SuKNzfK3TeJoqmGbNyV2LNSt+4
ioPCE3OBpBY8sqwJvGKT6CV2I8d+djRC/yp3vALljFs6nquwGA8jkhpLM/Ve
qWfCaZsZaCZ+xxrxkmm0SMUkXdYwzGYT1ciwrUD5x3eNc7N4Tm41bDJhPVNb
IvlaCH/aSbpc3pg3xwSEHfUzFLh49418PD5gVQWdMxGLKwK/X+BwHl29rxIL
T4sZUGiUwKq+RTSeEIlZAGSjxyD6k0ssGL4D3qU6I/Ep/CN2noTL/ULtjxjs
+vOjo7PrPYOgJS0wfT4+mIM5aea70zhqAyp8c39Q85pNZuF1dya9/ep4GRXU
dPQOQS54qvXzOapQj6/mVDrzbD4UvWP1j6L92JDa62emUxnCmVuFvxYVIgiZ
DmiXugd+UCi8VXxEo/kxyscMwtsQQ6WDDvGzLtlfOJc6LqjEp+nJAnRyw4dt
HTSZC1+cmhxKgDGL+tyOrmVxF6kyOA4Mra91V582UJh08MrgCpc2QlzPojWF
SXCf6DgLfgRWgq5Gi05Y/Nu7T5m2ecxRNWRXlFxam9hBnrSLI7aUSB4M5LED
hO/2Fx+8FJCTz82k3uADuZa+PrhBF1HOWo3/trQKC0cRWhlLez7368zJuDpc
LRWBjMv2Ijt4kYUmv+AJdzZe/ZvepJ1K4L3DoydvKSLCQdQVX1nwiQqrTOsg
s9Y2kBCI7crmld2NhpMMz4apLYZ08OHPq4LVTu2mKesurAdqTA4rIlo6r1TA
NDGbIepXvvxmWfY4WfXNr/+cyxOVpyL3MCEafTBWqYW0OVCm3a2BinzvFEU6
PJ0lic2QkWb63Mokvd7DIR9XPnD5Vr5mh71cgjPZzLdb/by38SI0A4ewl5s7
/v5VJeEYufAW3vVLSHXMLUAZhJdxGc7wHkvreF17JsFs7PLMVsbkWeCBRgA2
JCoA9QfeoxlVTrH4vS7q5G6Tuwq3NKo/0byEquhSpGhdSB1tGQuEZ28cDd+H
YNUWAm836QyqDczmu6dtbHxxHe4VP+wzXDlfqzugjbCgh3zqFBNNecj9iHeV
5Y7MTYGeXrLhlq1tKfqs5Xp0SMwfmJijfEeU3SpxIwpxWogYBzwgZQgG3yCO
DISGq6jn53CpYWqXl9HBU/8GAkMknqghxCer07F4f8GfTNZ/x3flziz7iOWH
tIXHDPtKBv9D8xMzgCyeY2t5reDANt4TzSs1dJd6IxidMdtzd+RfdYT3HMpD
VPDAdtriwo5qqnwnnqaTPVIULUqasmeN78riZ10j2dP07Iw1tOQJ+4RPgpUf
ddy0+b9k6z4ZKZFkNziW8J3ZLWqAlDay8LuBx1dv+jkViwxj3Av1YTC+SMmk
rM0z9Wd+n2qs5m42Uq12nxkTPBZiFWqHeqlpCttC+LAJOD4l3im3W56PpKac
7XLOnSVAm18/FDJL+GQ+dYldw/4yn62BGW77ivZt6tWaMQUCF4Ic18N0yjrd
JI+vf0gET7qxyG7+Gbk2Rzgxo9oFbVtCTo0t7uQ4pSRRC5LlYW7/TOg3KTbC
7xfjyhK5zWyMFpL9gM+Py1ef9vt3xGT5HDlnIY6dSGpXCdhM/UnWKQyckPan
lCMAHKl89con7N+9r8GeMoP+dlK/R1p3V+QCdw/123w/AYAxcmQViES5y5zY
y8R1v1I+HZJLgUO11I6G8/2sKPbNeZJgN0IqsU6/N92692CRcnmRLu9fw59r
mQ21x2grM5r6eCBUOq5QVTMdRVKWEfH3R6ufstM1LAaWA4dfUJvz2pvTL6OJ
qiIbjNY6X0kCc6ArZ8rwbAY/kobEhipp6T6ryeyorQlV7BRTXMIFOhLybR3v
0TpyXSohHy5jZfDxOiZArbRbqpGcIRNuX0kXW69THgcalrSGNKAM2UOPTgGn
hQtvNAsMelPEqK66TLATc+no/fyNAXjkN2K5K++7bX/bQuQwpvgZZ+bIJafq
oN+7Ixqx/qKnQL2fDIbx2V/oeSXsGwgRfcnA8x45oY3mkEPIDK67z8ln1UGT
HpBQYRuC7eMw7U7nsY5rD8s6WbtiKwvhGhQKsDqDSgMITpjqb8YKoQPkPjb4
WZ4jTeCmXCp9D2faE8qki4bNn1norzH1UQkmfYSf32Oiyqfl9YuwD/RnB/1/
2q8c919xwI72fKy8MkTi0fPB+ZM/s2jscJvIAXoCbSRcmyhNHKjwv4gHanfl
1/pCt7rI/cOJTlpcQbD8G/tkiDpUxa9kOsDOvGMBIhHEXGSxoAz0HPXxz8dW
2tZ3lF2mwLmQz84NRyq3Cq511J5mU+NBS3glCB3zjz1jX6F++0ZE7zy8VVMw
lUXJzK/xKm4QZq1tGIpBxgcZA+WoJ+Z6Cy0Ay5rYe9jicKxNi6wIVZqjLcUO
H/I5PL9fPgg9xxPilev0Tit88s7e25qKxYNS2s5PmMaQq4uKdO6mn6u3Njxr
K5Z2sJQWWvLvUsBYcTYcFCiAfoPKMNv44RHaOw/6I8sy38x+bIkw2wgji90A
teNwufb37ncXDg2Rh14tdwVBpv+/Ugxl8d6qQjNaeKXgnDixP2xc4MxahnF8
9M/OO0yKbITgvP00IDEyTMDPxI6/h+XPNpg3D46XqukLePOlGGLNIgaJ1yyW
YioYuwXBWLiB/OpZoXI9MDQxQs887ae6e7S/Xm5yHHYMg52YNSHUsp9qnGZm
dsaMZbQxvE+jOMXoe67hj5blyHyt+osePoNkSGvUxVSN2HORR6XbK5JSIHsq
LzOhglhSbGImVyPtdbnWBaCMOLNPRoUHAYMu8sDtkQamyUVIVdNFUoz7y3ro
pp+HrTtDyv0qA16mX2AhIxRQ68+id46UGIPOS5RUn5CsQpd/CSEHBQpZLncx
bvNgQe/+8pR0KVKherX77TyPIv9ApE1U6u6Y4IFlhGfezFr8/1TWpCaYdG7m
8mf6HMiKseyOIAlpOPIYd28yXh1GJEPK84PwfXCFO4BDjKcOoGjMHcCcNmXk
gC8mJGnbgcXlIrdLV6azlfMRuSom60pcHtl+Bs3+t475H4YW+UIJzmXXEkb9
Pe55u1qcb6Oj60Y6ECTIpD7gmlrRNMiVwqHgWD52S692q1FkL3+IXZA0qnVW
FyzJv17/JsiQ2T9nO4G/yLGnCWq3MRVv9C+OHqqB82NgJM4rBlNTfx531CSv
nY9ypNK3Y0xPgWGCj7PvitJjhOp7NON65elidxBuyfitd2F0Q6b+kD35lbIE
QN8Kcr7IN9hQMv5UqR/0Nw6gTbFAhF9plD/lrhDxihbhIxgECC806PGim+dT
eABCRcnLqz7NtIImZ2TyHQyoM3giredUTXVC/vryadeeScs2nXIrgiyrF0+m
W1Nn/9L3mP5hERFOGJ2hTAYSt0Sk4wONXZX58uBrUad8iYrcOuVELdWiYiJD
gRzqaX+qq8KHPRkvk+/1RjBQ7bGetVi9vp011BeFCS9s1AMZqUDm5oRvEpZ0
fiLe6pvK6++GSL9igX62R5ZmHn7C0SFIANT+ZMYp+ZWHXV9j61vkzkdoNDZx
5i85G/tzVV5W7Q97nBHmqFU92zOz9GCZMHxgQFQxSvh/gz3ta+lew63f+Pkp
Wvyvi1vcDp4LgIu3HGuJV4rl/QghhN3X8woPKjKbVPCQVaZfG/eglKb0BtA5
Jl2CSwXnixMAwi4Ra9MnWdtUSWyghgP2Hn6a78BNrJhpIJufQN0ndndizUqW
wEUbpUGId6SCV4jtt0LWl+UQGARAXem/jGXycBuyM8y6B7/tDOT831vCwPIj
C9/e0FCsfRwhoWXvcSZJEVCU3vPBMOUDQtHku7aVZlZEBoOvWpJJ1gHwZJZ7
u14QtWFdjw3zNPCU5GAqtLVWlh1gyqrP4N1vIa+Hx5fjqir2ydl7ZFoBXdUB
Gz2wDLAuPK+JmANaxv8E9HEAFKY6auPEyGoLVCVXT+/xv11ZkO4Nr5Nd+Vfe
5XG604wPjthqOUysmoj6v2Ts8OQkf+L7er37gKJeB9Q6qy3XfZgJoZPPLSN2
XhACJ1TUCyVjb8FvwB97yv3PI/qTzkjSwQcpR8gxG+l0hrYMbKkxF+Of9OpI
WybX00ehfBy3GF9cW+T3XP7Z19EUoCHoUI2y0aMWKiHIAVmd5lRCfsw+tPki
HTEK5QHs78wTskmxTjZXMtI38nvpPn+vDZ62dos5KimAYV6gD3MPKiSppChE
hg3pYrynUkTa9XUNVuOHwRIHgEjNTuxpqvFp5yvjGg7nydr4nl2szpYUlew2
uiY1KXdi3ahHvGkBhB0B/qKxbsRbmjkRJcPG7cnMdZfVs4nP+MshpcqwgflG
4sYX9uk5I37BwXx4Qv532DfzI0bmfHGeOZsK8IcxFcw2oYLBkh2mIgzlRdad
okTeMJuPvEhvvt/VgVb8FNTfxwCmux5Abb5UarvBJ7gYto260CJ0Su8oHnw3
bWyprynYBgnzwaKx4shTLqtvr9JD0J+z4EJUMAIZOXjvCM1unIz5lGWLDmbh
Ec/kJ2IPXNhQpenJUWAwc0SxvHrKmEpIOEh63c/LyGr60N8rZbFh4KfgGH+t
vHJcDPHh8fNPiC3culW8mJBqFy0HI+fGekTC+yQgHlMrh8FrE8m/QuOF/PvC
CUxdCb9nUNRMZO3ye+Xu2ViFXlspSypbDvD+rekAjUyIM4w1CJGvG22w4KdP
y2ksINyHTyuCxdB2/E7UVbDqNNnIrKfk9wgg15NjWYUdviPWYIHa7gRXwkFt
4lJD0dzdrvU0lUqFi4+eJ3i/zjvcFrCqhauVxd2bOxYrbbtpzFxudwJnQxO4
g+7RtiivNOIrNyOvd5BJB5mkcbebInxaDKNwBOEfnCnYO0OcY+dNx1Sm5/Y1
+9DXPz1ujXVYBo2twT95GNqN//WFPggFhtRvsYHt6FOcRnfjOo1m/JBF7EGJ
8CERtz59iLmkpMmgLAxlxBt7+0sDwDOhuDdScglNoihSQgVUuQQohlUIEqz9
+KxTEvbVped1cauI/l2HvGhGI79wixB6jhOg/dF5BWDuCC0IbRWWxngRM0QR
H3L/zFb67McMiFz3PtNRi9icmt2x84DmmdEEA3z8DcdeeVicsZaPhUpp5tWP
SLuZMNO+8r3J3+FXORaCO0R4piIVZgSOI0tEmpoMs+sYrXAICpSNeiC5k/oy
eDeKMjckVAKDye+hqf6Ddlgk6CYQqPFx2yOi1id7NO+4AVLItSHGRcpXFwl6
emildZaJo6JrkcQQpHXhFOnwDnbLnxO+vDiYERhvwCCMtuvzB80bk5BqZbOK
AFkPWMWYNbkfE54fOL7krpr6AB0QKCHhXRECm3ExToYqd7d3Gk6YUtn8QoFJ
mldifsqC0w6ZiYnZzWm0PSxfvHM4uMfWyUuNkubIv6kZB6p9sIkGBwPKZKMI
2/Z4Fdhj0d+FgpvMf89ryPKLaCaHdoLFek1bt96bzleQb6baC2ZhX6RPdEjw
goUwcWBvfPCS1kcm0ITgG2s8qlvq7/zguW7iI7vQEZqdsuE9ad6xTjTI+B7W
s8LV3wC4/5jtYyWlRlmMBtLLU/MUIQnfwd5+9IiVSvCppSnDaF64RXagMwGF
MupcBFRDRInHO99bwuj2m8LcLbuug/uW24pXQAZ+PuGjqqp6/6NZ3/b+CqlS
EgdxRDtmWj9El62nAfcY/3jOOVchcEvtfFZxUbO5lq4mvjpZH60cn/2N3n9t
6Xqe5JKo2TJ2WEdHR/f4szJxaWikMsIvwDq7d8vZFJ8K6uUoXQFQu//CU7dy
teK4iTJblsY9CHYALaUoc9wreVGXb8K1IbPpzeSry5Ug9N/arkGQL/bBBeLJ
bN/oGfrVDuJUxKaDfxm0A2OylPPnr6FfxnPZxxAExRfKH7vm9rr7PHXoFzmv
O+JtyFH+Aozbj2gNZHyHR3w7UCr4jNr1lhimAat3iSya6x5i/HYK0DuokUs0
UHCVOP0q8WVJD8hJhk+B4GBssLUHkqGGxDsSkuZ0TMVbcguRdJX6aJnbcB8i
hxZzHWQHZjc1JG861Ac22536JvJuiDmfNntq0akyvZ8TLprHxh2AWv9s9iYX
YUhIxJjSkL0M66byPFbVBfbuoNlkvlHvXpFmH5v7HyNUYzC4+iQliTyOGulQ
CoqeaIK5P4QrCiqxInntcCMGvVTKesLAOkPfXHw+01qY7TL6Vk0hGnlPQWI+
GJcHfUYdmH0ivnQfomr/q62TuSXFjzb8gyitY8Vle1IhM3Ww0W39OGT6jrBu
OaIz6xPT0zc5A4p7AgQwlv91k5hN9ngG3Zk51EtWCBvbbvdWNlKC2bhIPEq3
8h74/ekrOnlo8q7l349+XQECaLsvbo00w7UGCClV8q5vT1bWeiW6WEH7FdnK
UV7RHCF3ger+9eBG73Z5b5ozSxuorsbxLVw1SwJLNn10CzqpWaqipHk/j7tZ
JmjdMEN/6KEHhdbcgAqLWeguQ6zgIc7DR0l/xjwN7ZsYl5gpkxLjk8vBkiL+
M0+W+OCKao1XqO8p+n7MjXYfypQmeHFlst4ILIuHQcp4UUOUutX8i+qpnkNv
g/vl6D2olgf6NJP/Lg1Kf9tGHhFYxnf4QD/CboF5hWUMj49k0GpPwjOPPz7z
GVuGwOv0B5bjJlteqwTgT008QnZKWrw/l9uzldcujJcNlk4lCuXb1uGf1xZq
nYtCvfwqw+hK8hlztClibbDPO/M7+nhD5f0u588U+Kn70XNltcNZXly2vkMH
xN5EpmqbIGRVLHUHdMDdEYeMav/+0K7Dx1xQ0SZh45BJr+fZNRHebtCk7ueC
XAKZ8R1yhl+DmKuKHP0vMAp4j2nYiPM/Gol2MZHNq6DScqkG/KgK4SPtMoeM
QBj3+iXuQTeWZ2vBIbLvORkBgdnvdTtlr/OHrfGmtxp98l7LpSNdCgXVxGNX
73orOsk1KsY9AsnsHMjWjjsU2xiUptmjM15wedfQ3a0FIzYkaf2zvAJzQU0x
bSVBI+VLaqs1NSEOzmWzZ9O0FgsAVBeqhy8ye406pk+Uc73jTdagtgNwpsBo
JsRMFi9z8XMrl4EXJkSQiYfxpbj4lcSJC95LZiQcdlN679mCA7lRzpI4/MWh
8ZkA95R2yzHDi0vhicr+zQ8EMgnDtee3F5F4k8C7ja/NBO/xjVNO++kRlz7k
pd2bbgtMSovq18JoBj3Mq5BnO4APFl7GtyhgowlVa66EdlWD5FCxOxjQLmqs
vcPWPDWOmEo8tbpBEymM324nQw1gWkjwNwdhHi/3nPbYQp56YezWZjdlCNlR
9aUelKjZBIqapEE6iTAmGy6L5Lsd+7Q2g2HNNJYda9l8oBx0GNgDiQ1KycUn
ccUl+8l2MSa/hEKiuTuKB30S6FJeDfwgns6yOnkkyLwvfgeHxR3q6I68B6Cy
FIQCs6rlWklZcQYPp3aJCoxW3yRPKOKN7pnSZxjmfHkZNSP9XqsFAaqfum4y
VvmNL9iOFQTJ6NKn2sHRck3YITEm4DR03g0x7dz3xeZKuuTvssFKrrkB0xvP
WIjkOluy/ueEicD1GBVSirmO+D3rYzx23+odIMECKvsU6GvLBVGGRsD/1bkm
fhM0k2j4nJ9DBruQtUbzAfWO8qpuSE4rZPX+O6HCUpiyz66UvlYoRyvrA4O2
t4yzCJ1cT5dy+alh9iikD5z4dzPOnBjdYRpomW3rPtnxjNB4qIKCIKIc9GMW
9Zyw6YJ98sczFltcJp/tSz6Ki9/CDrjxtrJeKOgOBHUfj2v33/izNMHI7SuI
poC4Kbf2V4tfzcgNgMPlYHRICP4Mg7TuQVeBImr1zX4XKG5q3W1XNvOtSiUm
E3sO6Q8I+qsc/9q/A1Te3kFP16OR4x/5nlORoqQGsMgJivjjTwrjMUkZYcBo
cYpY7dNAebdlUxerOk534uzmGyL1jnxkqdX/qVFb76XKEj/7fEiZVNZR2GIB
5qELIvdinz1wTv+LW52h7YtZRmgXJoTIm2FwpktEK+0SYgut7gIibB5R3Ida
2/PdhGtYacoY2reBRzQYL3dxM/H23PqF5HcDEYSaBiu4WgcQlzrWl1UF0h3e
wc35KGR/Ytp867Kk6Zrk23oKJYqezoB6BWlzpS84/mAICsYtBRkkQ7I8yChK
PAfsNqo1yk+gk3RqUyvc4tr3x03flMtrkPdIkqpt//IJQhjqCCPLsIPgEGin
RpNkpVyfKhhGDnxGU/YLtnPWVwdXvQoVyYjZTqw0gEaZ+tAVYsA5ryU9AOhI
0xeehAQdg430aAARYGO5gL79CT09fDwF8Hwl9qy3QSIxLpYDvrT9sXKHuGYL
hpm3M6Xu5BNffcEPVAx5eY0RXz9CPqswYH+xfxZ/RiSkHfUFUPA4QAAWEhDh
eA1CUiRXXIqY57AxfwvrLZN7IUf227o58RhHwGiOIencMnC9SuqwUBp4EU9I
fM2B5XqOpsH/99dBieoMfvZ84d/Gs6gj2+IAoO1c7fDZAfqcgEVRl6SItVm7
MpnE6MaNPVaWmke3fABTNwisTx6IDUBKnvj93A4OQi34b+ss1C1MOz4WALkl
P01memwSszuYIlH9jn3Q8O2zr0+Tb9CaEsPN3hTSzkdeoizKh2XYDFEBXoFl
dLsCnRPoXF3HavuneR8NXeAAXOFvNng1+lVm6Uw9C8LcXy31htB2zdoE2hlz
iCL4eZxNjm/nL3C3IaBT1sgoqJMJcVvnaU4DZOtmKSAz2KucJFZ/mX9KJzD2
OD4KfcM7NjL9lN1Sb5KQfgOdmJmgLXgXleXhDiyRKi/fHCpnZyRlTgATa8aS
4BZDzdsVYvaPfLdWvi4OpbWxjx/qS90uUQ9lG1egYrZHQzlI9+x62D+Ovjdw
BHbp8Khqd8jDOyhZQQpxXaxq+ufqUipYzZTg3MLSubTm2ei1LbhZuQ93jYc4
5CCv7kYFEsFltlkJocBhPh3f3C9T7mKXnArlYHFcG+YyXqXRo+w1cP0KdaaO
mj2bUT+QJadLmWUIkTzP3cEauYs82O9VvhHH1NxLQbMN7vsIXLtja3EimHip
lkf/gX79GN6xLRcttvecjBzQ96fozDVT7gDkVWUspicCALiBvgusf0ZRW05W
d6aQB3Z+vby52LrO6HMnqzwg0FxGwvuarO5XwDM8ECLMOZkma6uVYogYFztu
MMtRbB1SytpOgef8yu4TLqo11/M7/CJCnBICOgVX8e6rlDFPtXceqd0W8kKT
nrloXBSxLmcMGgz0n4iak1mtdH8IM8MpU5lJs7S1oWzi19lyv/jMN6GI5gK+
cZGxhkzJxJn/LCBK25zKpqhRXcAcMj+waW3iQVB4PD7szdNCo07n032sOieV
5Pq6Ov6dd+otsyt2CZtUx7aA8qP0CVQI/1ACMJRSzr9o00bOxXFEKh0eRpad
5gQDRfoxsgxFv96mouGPJOhZHoObAxua5qWZuicyqeeXJHUKDXrUKfwjokVZ
sO3sqVpmIma9WrqUIJ/89j0LwLxeq72f63CRwIUXTpStWkpAgvBZYMgVPcmn
Szpvhq37UnB1gc6kZ345gH4HBcs/cRBXmFaWI2YUCe17cOLSPzb380I9ITTI
vKCmQBZC3ZV49fR/9tCh9oTgv3y7ut7I5MYXO7I9GOuW5KevzJrcbtpOnZjJ
jjX5RoGQy0bLj+QMHKiekrojcn23L9FyQ8mizqNns1KeG+0Tv41KbwzR82Dm
odr9/3xoeWUYC0JPWUI70lQMc9QMMlM4KhqJQOMTF949SHBt+ermf4K94ci4
DaPuqt3SIc7JQMHsWlDJLPf47a4BsKcdYzjMl4IYT/SfoJymhOfQeO2p/7ds
IbORJuzVGfcwbtx5vYu8Ov+GIqVsB7KI4qo/GhMdpHytgSLZHl+1tKjxCltV
2E1uOkesqgiR9+A58hu98HUE2HdkVQgT1hcVrQk1NReNYA6oVzYsJF/pTfa2
qne/1rq44vf1AgPUzMCTSAfXv/OteR3X7GrdK86cXwfWHWzoACEM8Hyj0tTP
x3zYSs7o52wwHL8Ge9QNWl8YNt7YoSNYstlGk3V3YnRomxZOeqV0ytvA8XDb
kLoQm1PZLoZwVGo0uozclIjc7ssGv1PKG55zsgUEK95it1PdyGrMz0W1pcfX
UI5UAZcJ0eBSC0hIL72blKbZvWqv2VTi691zuLhKQAQ394u5H3S+myvHFn25
rQfWJr+jQCzjTtfwmTCHIE/jkHQ0WbJHkYeIroFAS4Yyu/NV5TGVU6TnFmLw
/Y1czMGm39VzmuX0RJGwNyUYH+tBjR7zcUogAXYorFRm/mgCFKtC5wbOCX/u
26ZSv/nYf7HwIrmVwrgOCBSX2QGfXPS9sSlmRwXJxDr6lmQgDlKgMothjf+r
dooEAH82HbZ0Si7vOm+tAor3MX9hnbmv2fKkHR8ed/A6YpgHT7Z/1g4o2Hyi
VEJIoXu5Nl8wMLUqyX5xMeK1TAVBLKb0AatJU0JbNKZemLyctr9GMWP0wJ2h
8JXafdmz9Im0/mhuQ5tLlhfOBId1Qxc7+Ecn0cXDu9Y898FZFiR+MF0o69NY
Bu+LlD7llP7Rt/BhlB5tGORGyGdAW/x6dN75ng/dFX6P1frThQ3ms4fkfgqN
Ktv8pIxrV+4HlyOPIa7ARBk81/ZV6nYIekX5jhcvODJryaXz+LBVYZ9YiWsA
cskX/WNytSmCyroHRBgMl/hg3VJO/VGv//PJBioGKqAE5+q5H5orxpnptyK2
1I6rFf6ikuD9lCW8c831TDidiV1SR+S4va5kKfyfungnjjGmqy+aoJve+hvT
ukfsMHNKAB8kS1KXg50pBUuPkQ6Hhg1qrZFBHoVgS8L9x0AVY3mLOCo/lLbB
Ws7qqGGYsSAH4kHjXvoDzTbf4nf5j0bhvEw6r47KYZQ7nPboqRE80RJYjNlW
yUTsmtymuuF2accMgsKy6NG2DJJLLGrYcqby7ZRTg6ejwA43Ao9bkFDQ22Bs
I3hIQUUqkGrXb4fJRMEjPJmcppyNEKzKLwBCw2DpzdgHyngwpe+XKeik12hq
zsmV0263nnul18rTFw5KOzwLtJJCFatmsVUJoStJGypVBacKgJgQKg7wLYQN
J2aoHiyEMqbRdhgnVjMPR+oA2Jedqij4fkGAV2BqPDkd5J1lmP2bsVPHzMLY
J2eJp6WBo3hp20Vw0J+UQGGThqSj0aI7IU+SmwdoHiUJkHUUtgg4k492kXvc
zjHrclhsLoIbSKpea2K4gGYCVfH4L8Gm0WTW2t/rw+kIB3t6v0UOfaKPIMw1
y5fYrJ4lhcm0JoBZWvO/BYNi0ytv2e4r57nG02s3iTNe2qBZduazXTW00zCb
aTEehrDmsQXA8e8Bb23rpFPYOWxom3iJ1mCOzA45Q7AD13Z219n4HOvVEJRS
nUMgssmQf6CgJFNv1KjrLX2DmjWBkYgQiTtzbWjEzJRFwVU5zar1iNVr7CIA
CSpvjt0oHDHNgEMkzbkWDilmwEtGi8PQ7LErByQ13PI/5I3i0B8dbYKZYD5w
g2SpIbMEXu3PcmnLV1eZWTH/U/3ZSbXbzQg/VWtf7YGfUOp8YbGaOExRhs7S
RE6XSctf+7LS9FPGwRAaLuh3DojKuLJqQ67DEA0nYDPWnxf+p1hVDEYDKbMv
4mjc8Ym4r3lP5oJ5qDF1WYZ2mmiXUD2uwZe3QrdTCbQ/EXlANPUbrp/PY2iV
Ppqxb2dIO7RQsFVE/fcm8qQnbbdxe9irKNBEmMy6ih7k9662V1HaK+FSndJT
9qGF4A7VNNT5DegQMwLKO7w15LD1R7trqE5RYx1iItynfwuZlcjrghml2DGP
rL3SZWVukvTHCou4cSbpocuqwIHDnz9wjSc0pKfvGhkdSok15G9CSUY55q0g
KGNAJ455gsgY7bUDrNIeNEr+pKmZLn9uZoMDAo4xAp1Pva9YsgmZxtVX6qrf
Kou/2oF7EjArK0FTgUG39UoUc8JiOI0AsNJktbZg5NP9kyMsByHMvj3sn3h4
y9uckDGdZ1do+L0+HZhivLXJG0EuaLAhidgbfBlkxORnWjPz9qFUZgMHj+ro
Vbmr2mtsuT5MQsqiFVtwGzapGvHXKkuhSqkV1pFgBOochZvZz9ZOnohFkOhF
RLEAnvYtYyMO+mTfa8Tf9BsU4LbgpJ/2/J3wzLAFuA1j/4kK9ME6oUQYU1oD
zHDC1UJv/XOlxOwgxESMu3DGScVdL6MV+9qIMMULH85xX7VWeH26xyCHKRUB
btepyLFGhNz6KQOpo6FVpeoPYC9XcprVL+58Nk0YYkpb51FGJgCgZUqyYvAq
h4YLGmn+Tp4jezD7cY1K4myjfI9OrYIz/e1WFbHA34PRL0+HehAEL5RDgrC4
AX0+9cd6hojHq9T1rCwbos1fNrUvz188szro82vwY7OAItMHxp5aiA7GZZGU
YwMF49DAsj95s+uXn9/7hiLMAZKo0CO8AdwTuC/TRbNzI9oC0wBy/P4+IfRL
Gu0SWP808Wh/az+/uAAEj5rdoeaiPtCkRaPWiEaGI4BLMu+F072Wdlj60mGL
f2xro6UoEq4gX4pKb5UOlN2gLvrciqQ7wLizlq6gWOQW+8ttpcOtnzf0h0AI
IeN29S9d3EB893Rm+3wn21psanPcmKiAMsU6t16/Tu53IHxRqNVMZhvNviJ1
669nFQHKF98jufqpz/F3rApFVLsIUr525OjTVwjTbxBeZr5508c0DDBz50Rs
BJMkUEjOau1tZrwckFV6S0nB4/Q/njyXQ1XtWHApEOrHXJlA57oqDc6CXXNK
6XPQTiE9ACQHUQllRahxwxtWLxKcmPp/6+1GIQvl+H4Qfr87cZX8YcmMbGjK
w7kVDrBdHp9jMdw0Nz/HcXG6zGyoEzSRVQTGsZLYiKuqQzGBg0+sO9R9IrDp
EEKCHBCdC3SGDZO041ct9dgxf8Ti5Sfc3pbR7Dy2ku9Vd+E8CikHxKwr50HQ
if0E0X+672mUNo9PcigJIRTUWEtL8CozNMZqd9H89j2ivCMUa6MqRVTPu56e
TwZRFoYFS5TgKZIYvvAIBXY/1vQSk+BtD42YftATTwBaweoVZkmGmu4kw7ib
zXTE6cQQiuTfwQyF+b9gJGAIOrfVfFcTp06v7BXpTk22DT+K3jZa3oZzcVu/
yAmzYZ/0q+odal2293Flhch7mtilUJfDrS8sPv1fDOtbuYjDqANWFJeA4XTP
MQaZllPh+OfbLxbMsuKADZ0n7sKvHNSXa1nneYwpLlefqtqUYNpo65flA/C5
v87pp2tLyxEXKtoVJJlIhuVxTCh79M5FJxTl9CkjMD6WNQ8KUe7kQ3OHvSgt
HcXLa0Au9ct4WT+V1+2e+58hqm9i9QdWqh02QKWuYAs0MFvu3NOMKqcqT5y+
Lk1T7iO+LZSkN5SvbWYVGJYiDwob4DrXVJXo6Xgqk+QgBPyen5yiFM3MTuPf
hI/mZpp/ATrDYFOsdlnzeqmcVHWQhSyTN7GczOna5zWuQbQVMtNs8opxuDjA
Cq4bXRFQ8YR5lNv5VgpeLtgbEUIMgmUdDJvemSDH4KXfruKmK6SGJIyki/CU
v7OmhfnOSAS3UQkpR/3bxqe+r4VR9yC3/4fvkj68/y88sjybGXqPLKZp5CxQ
KZwhI49x+yA0PXzXjYGb2xZfSze0QaFWIOzHVCni6foj1HhENsZz2O9wneZc
2l2xvEdYzMHrGNOqH0+RYrXAMst7g4kuM2RHh/9AU1b8smNxAjD/3sPm3KCM
xfE4gzu3POS8zfTZi9eeAOlhWvPaXDklyB/UgV+ofWLhWJFNjr1FwyymluAd
jVmew+pggBbBQjBMPRdpWtv8tk5US4G9RXwZT4GeYOky/w4QxTrWuGsT8rXA
t1m2tLw4xNRZ+fBtovf7n+xLPwKbKmYHYCV4Zf+FTO4sMD3sFwLzzdbrsoLY
cfPi/eU1E/oq2E9XOcITAXy0iSbzP+TXbcuvj8Rzx0qJI+E5FgqqIlp8eofH
2FI3SA37Bt5gyYILo0203U3q+F+AzRwJ78EWDN6rAw2EPXKsIddNSE8IY7zg
YSaT02U6oZnqAXU3bfEHKJO9Mt6wfoiBvKRRM3bRwBd+yXwa1dYfgipMx++9
nOtS6jZdsH2RBKsVN3MOuAPRH1bOYi5zy1azyIlUuxb6uurI2xsaJ35nkZTp
W/3TZaxTsG54QldHJVhbSvX7qUQvYr2PXuN/or7R25A2D1x/h82Aybqm8bjC
kZEl309u4tgVArY5NvU1ZSjdDSjIFFn9/VDOAXoh8tKSiPG8jSTfo9XFrILv
6O6V1PU30uPE7T8lZMFsxrMB4GssSQh96dyUJQjnTuW0oFkl1Px0dVj/+7Ta
pUTvqxxp5ZZR8v/vi6VWWFcG862Kd8fCVaFCF1DEMjXqePxWTInsOBptk9ry
hvwTlD8HOSnceRJ/hukXLyPrwMe0O+c9qado7m5PIj3qb7e72w9zTsUVVseY
avBthNk+ou3ni2OZLfkxzNTLXmjmDsiZNskzoO02kpQMt6KuS3zkIMw8+s+m
ReyYpNx1ix9bfL3nS8mXGin4WEwwCd6oL86jDZ2NZOxNK1ckniHmaIZiZpup
5hyMzJrgahgfTOxLhyx98QayJAGd0wpTDqyozMpMuQL/C43bcr+cGb/8isy8
4NA9SqwXXAOyL8XUKa5gGEcdJtlt3bJd3U3Lzy6HA/DuYujdXAD0Cs8pW97k
vilEhG97z/kyKju1JG5ULPNtNoG1K3vxy+xk13TDaW37gEbehKyF6p6NwVPL
DBaeZcej/FyTrn9ZRVppFfMtM4aBZrg8q+DingdTkwlM5sbjBUXXmzKG0MDg
0y4D5MtqHecEmC4CkM4hjKcoCZhB5+REIwP+1EUbalqmRophy8vosrkno97/
lbVcQHnwiYBTlceXQopQkARA7X3O4zk2VdqWA3SP3d5QHqCwHdcLc2dgaiwz
hB6Af1P32+qWZMEtbbmDiBcjN2HwTv/qg6Lbgba8GoBZuMPArshFjOgntwNd
LL/u2Ck1U6ephRPQvqv/wz67dKSE569r6Jrri1V/HM07ffnC6Ng/jSbPp53F
mOhyjgF9a8AvQ6ZzVADdjiSE2lgCGa8xoy1Ha+YmKZ/yTrUe7TzAXLNN413d
ehW7hpovNXqZ3IkrxeiGO8dX4oJnfhAcKUohsUJn/scsf6EXrZROkI7grTcf
K6c6M4m/c7u9leIe5qdITKuIePAerc2Vn94562wilBpnk3mPVp2S0LrOpvYh
wE+9HL2EOdIJO9vsZf/9/ik+G2RL4rzeeYtZAGJRWTEtgtRqEwoRiUA8vj68
fP8WjYdCfHKaUQjZwfJVix1de88TVucgKvuVXIFInGmRh1lLvjhtZp4FaXkR
ePf+zcuErygtb7odSRtolbGl1QTK2LJwLX78/jTXewwkoOOG4AQ0krAaAVTs
SedR+OXlCDv8aTzpScvY51G2CkYMqMaFaqm0JqQ9fce0rQif9Sosi7gvOVen
ffJCdjY3iCPHNgkstqkkfsC1JZOixSHys4N7nc2ld5hBecG5fWAHDMaAa36u
HYdtOwcou7iMT+IWhjiC53s7jYQAnSai37b3DabeT3GoDlyWJb2PKuCnh0Gx
p2HHXolWb1v3QCpQ2RQqUi/WPhoOme3PyrUi1TmnFYCgnGjFpCLwIpVL4ElA
3IvzrPncrl8cxnCdlvxxowWjPqFfp2fPLARpESaEGAiCT9/wNgr220ssEFlX
ABjc8zRczyA0isyEf8+k6uafhyfyTKD/OJsFHoldDNFQuhBr4QQ3myTl5eoe
6kqpZk/rja15AQwyea1hoGHY3xf/7TYsXXu+gM7uwognzP2unkphL+wo06al
dXraq6iA8RiEsn2L7f6FTcjCTPwMSX8spAzqrkqLPfdZrJpuNpEzOIWAfXSz
gPkYtfgSwhtslRGR7BJn3MaTWdR1aF1rJA2QkXg7qTE1TZKtB2WqWc4ewPgn
9PCnHQuNJsvA16tocVjHpERy0EBmHhOezZXEZhGxL0i9CTow/GwPDR+WkoKV
TpSxB/ocaZMcBXsWukmSbP4qLOHeOVqW+S59yaaImEI5aKePxb9/mBxrE/3L
PsjwO5S20nMOMP18wVOeBbCDvcvgidSIzwDrre9mbi6kTUkNYtj1ItuLIWG4
s2MbMlTH8A1txRFeAF2Di8zYY5XXz9Mvct/nKQkfWDPj5OvZUqv2QRvCrX5M
cHGRM5LcNu43V1mXqtKlX6SC2mNEEVH9imPzXvCw44ApZv/61hWEbxJXGB4A
rpTay6b8awqddAWnqrs0dI+FyJWh5et+49UjYryGsIBanQaGHrb5/pyI+Eui
TZjV/1SvQ25Zjtg6vzAuXFzbr94rnrMoFR+g1FtUvPe4mRUQ6f5kiJeJpDs1
5w8llzUbGrCReZUtGcY0mwQCpH9xSe7zZ8QT7bkMtV1okPwb1uKd/l61pKi0
tIAngBbe3UMUjq8qrztgWSZo+V6l+qOhIVHUomV4i/EEj/+m90YGciTuBpSb
taiuchqtvVNt86C3ivsutP2YNMIhFIee3W0dWrLoW9J7T21JuQ6rZuHvr5cN
cle/PfDRDR3RAwEr26skqprFbYmmhhdZ+ZhQuWYXYNucL+rthhh3r1lDvGVQ
6kfqeHkSRC1WC8SOaZ8h5bp4Lv8pHTe1Ps5EkaebcSOHHnPjakVES6P+mnv3
n7dFp50fIZ7g4fQxtYuiMHrUvmX2v7qhXdH358DEbbfKfiArmeiBdpqrjFQv
ZqBdKGqye93A1rE9y+rlmr5rfncBQE1IhneXhUFJYZGDQO4doM4w+xEp+Bwn
NwzPjU8ClW/pE8WNUkdWG02ue7cDL8918kToGI07Ao8XJNUZvnXozMmIdnH6
9RS2RgsokXURrkXyFbFfOJkYCC94kpmVsgzX7h+O7Rj3X+Or6A4Z24E4RY4X
cVv7WVifNUvu7DSCcVuRU4a4WP7JoYh1wudmBmdoq/rfy2RCc8+qqkpehNI0
KLBmArSzFxjo61eILlJ2AuxmuFw1by4IgNp1ZGtrrymk9NdlQnnqFLJT5Tmg
kj78vQkfkgwy7arBGKk92Er+KxwyaNkTpOL3fO1yEgRU6t2jHrHdNI8gknDJ
k+Fb0uCHRIvZA3+SMXPzPw3IZAamo5kzyWjWzhttyeUgFgGe/aPPDEkGBIg0
S3rnu+wJ9uIUg9HyWKhCLAmKSF6lXoF5JjKD5ImrS20P2MFZUSQz+yB0GeNp
H5RDlGxBxkdGu4HKo+z0Ag96HqUhwBTMLkRfmnC4XuNSwCGa3um3tuvAfc2j
fxIbVduiYn8nqsoy0dS3z+JI97LEIy1dSa5hFl/aJI98CeB3Mhdr16I7tG8L
XNXAjkWJyE4jNiDnI+FNOuFHjDZN7/TUqxbjD6mvZQeHTXlYSoIL4IQcZ9on
J2jwOE4cfmlOId6QY4A/kIsa5um+HZZpDae9NL7liB9EJqW6icNGjX6az46K
YV6U/9xLqqxVrRQZV29tGBoHlE06cLWRcL5qCPlNPbM7ia4AbYht60uOdMNB
nR2lpmlnCo22GzNh4guZoMrk4VfDFtZdbSVqGZmjlTbcSpKp+bfHq0Ss+8xf
dIUVYGNY4sL0Wci4pFCZg3Zjca0C4unqz5W5Q1UsDXVN7KSY3ld8e4JfdlBG
F5y+q+zYYaoCnqRpdss6OnsD6KzqoOZRDHsBFTZ2+xnZVgN2rDhoe0OQyH83
u7Ze+LHgv9qn1TMwmN9hKog0xX0si7gimlmIBe+SxKF1dD3Z5Mlt44G+JF9h
hYfgzp2x5tuiL/Ctemk6qtjWU8Y6vJcRLjd+xbY1KoUIap0RI7oXH2EFImXE
Y6brfmK/dT2nF8TnOnFbyC+vHslgOYqePpOuQOGl82zGuIRxPDZ7UNQ00o9l
Q707QZgnd2j1P0GQvs9A1dBx8vAXigDrJT9tiQsATtru50tzxpEvCZ85W/2F
ZQ/ix21ryq+oxQUWWY7lfS41VmU27VjzfRRg9gkycYhBMh4bI3LpA28db9Oq
21kCN0imuNqfR2SHDuOWInyJx/rE9Q/ZmlB8PeC4DQGCf5wL91tsxI7aijOF
RUhf872o8gDOBfbq3yuwNLLnRLhgGp/6+metrMBY7TOPhgZdZRVyO7wda4xY
NxyWXli58uqL0FRlA37i/c705SbD3ALGnIChMr3Qbxn1EKyBnJBVV+Md/ae+
pMyoY7icYgEihf4RD9IFBSv/FA3hWBfWeIOvFWXreXd3OBMV1BtQ7tjDamsH
72ivW0Y2j4TPfIIEi4E0dRwLxytscAmHaB/Fqmi8Dp8acumhedy1AXtnbW0B
ORiB8Rpy9idw60+stcbGRFi3p5mzUF4j1ioZXe8fD5rn0Ny+oe+WUHIgbo3I
tA10mpMoaPenuH9vkim1O3RJ+SxzRhKekssFitlIXZ/BXRftHtJRwGak25le
2aWcMbBRz4uOs+N3UwfdKoW8M/lW6kVooFQP9Xt/yj/0q07ZV8o54q2BlHM4
k8w0Nl6IyqhyNMW/Fyb+KhUaw4GUVxrE10c2WEd/kWMlOuNtFWFZ7JsmW0A8
ek/ZF5oPVm/5Y3Kf+82a+/fbYI2DTKHCIFWl1NglbArG7L44xUqnqopPVmqB
vOwdjJYlUNRL+Qzrm1hJpXy5qgKAFKDvTHOXVx5QYqSFmLgINdbKzsExLoxH
5D920hEM7JLxR6BjQ7M3Wiq30yZk/tXis8pqx29C3YJUw/87kZOkKkewuCkd
ehUc2zsPala+xaftHmKlFzX626gPa+k3GGLxHJ4tlMWoyiuTzK2Iyc1f2wvn
ipbHXeyAa/F3/6hEwi5l18mbzI6RxZ3THA3xljmsclLFtC0OpGzptHKHWSgg
cyB5mDCZrmSA0k2nvQKi/EujduuG2yi8WQ+c/UBhCatuNkVPFw3RHNS1q4eH
T8ebGw3ogL8F3fFOHxdX26Vtc0QlZ+xe27qrMKG9/jumKScXVeKxppNZuAHB
sa7fH5wEM77/aJsviO3V/3pQnNFDZnVI/EoZh9MhFZP/+eARNkR12zEM0Me3
OGOuoNgF5uypsuwgMRB0PN6thQseg2fqTkdH9YNDhXPNO8KJFWAoEPyF/PXs
Rec1AzNklHzrIvY6zHNzx96jVSNFi5nTwOwnLRLbT3PHGkZ6Vmf0kB7bNMen
z8COmDqPSLABTGXW69LMbprknWF6wReCKYr+9IjujBQsNIQY2whnH/mxlnFJ
a54c19OY+xR/eEOHHSPWxzD6gkCbtJFl7pBz/roFL4DfpX+fqoUQvUPEpK2o
YSnmI+NZSOwczxZ36mfwCZgZS+xQpwMozoQ8RMXhKRc6yzuGhIGy7d8eGhvw
cefx734pYWNQoJjF13Ktk1k/k3p3ZImRkKtXse1G1Y4sfUutQ4UJV9SOrd66
poVvQa6WkXsfEGfAP2WWO5VVvqr8x4uu0jF+KGHnjWit2V/KweoYmv1K5oKw
a97jAO2MkwEq2zGHFlqDQzVhD2yMgQJLpjFQbc2hGSNtEYxxacUIGA99NYEG
UsMUArbnpc8aqEXRPNlNWEqTcIx/RMu9dFCXz3YkUvPcEqP5y2I3cZh7mWlt
NEXL220z0M9ZnmVbkCryb0VSFBZ5a6E3nuQOsSn5WLOdKu+3xjkulkLjnURU
TiClLj3WXbiWgOksya/4Oq+U2DtARoiQj4FQvJ+b60bwjZhDJaP5a1YstEzi
SQ/61IvUHWaoPETvy0KdDHcqyOVgGCfxEQOlo5uKnCnxNKl39Er5FkjCSr9u
taMo5bcOCZbkDZcCicWGadYYfdAedcGoM6jUos3esl9htVg45xTNCf2Hc771
pge+xKrv2wrTPPzxdII7skKEppoJ5+A4SLl0hdtQzmBUvmtGUkY2dcsQE11e
Le2WphwXPkMBsLpvbpQBcRC6Vut+c+6qbwcE/aR/X1gOrLav5LFSTYlIKpoE
BryQ1PayWWmdwCPLWOzFjAQ1QGk2pzXOTRDu6+DAZbdtK4BpXnQiUdw3RUJT
i9i5OB4qfV/4o8WnPKqKPktkZSFJVKadSvzuq1MqyL0bsKuoYGu6G2ih6FPP
S8Cvn6Y1DU1GpyvF+Ne0t+KrI6j1VSmf2fldZtp8HkYcnCSIKT/MLPZzqIOs
2xI+3bjJs+TufUPii/3grjnHXWKLikBxgLC2+YJaO0D50npRSLjUDdmfB/ge
6KALhX5zlUa63FL10dIpuNmzH/2AE1qNWCndDR3OjrdDhUL4dId7TpyAFi6N
ViB8LcjzcRcOMVT1QRI+KvmQKFmsl4uV6c/9dk5o2z4Vq4jZ89fHQfkldbPY
JXBioDYFwQKxHynYSc6huogJ1yIshzu1pBrfK11yn2Nu/x0o9sRZnFzh+T/0
/7oQNTpvE5HBMii+ou7kcnjfYqxSpbFtdaZzAPmxoS/3NL7GaEl5u7z0musT
1Donz9wRj9KgYBIAFkPf8ekyflpPyFufWPhgmZB+m6Ak1DUmVNOm5ixGUfsG
NO53gDOgTy1F9ydla2+WBm6cdm52VtQKdsRVhHw2gsWyNxNmBmZvj0G/4ojP
tfACtk9WOgDt3AvmjDClCSl0vf/A/iWNRtph2V0v0i9OZt0teSdHtIUjvCOr
M6Eq3ReMqNZ0fWHPwai7N8/vVisj3BWx8g2ieJooAXAohz96xMVfQizL+XMX
H/Yly4ewdOlOTruHYLyU4qMnrdOFoQH6+WOBEAfdsMbE5rNZqcbkrzmEZ+q3
pLZNNBvyKYR7eSQhy2EXUmSV2XvUidyAzmiWXdcYo+edHARAYHc5VcEWyYeX
f3TeID5KyTz0jQ1ztnThwD0AbFAatRHemR6wMUFU8bywYhVK1jkUfzLNLV9E
84Z1oUCDRb52o12x9J+Y4YWfQn3xRi7uy53WB7HCd3/6zWyC+yRavPFHUgWb
ONDW5Qo8oFgQR4UXJ9MxK0iRgvkUcH8dMszdVz6VOoC7as3SWYW0GAjvEPps
frjJzF6VQOvUHix6QKgu/PRAxDzXHBGdYPbM5bz5JxpZl4Xi8OmG082Kp46p
o7IVTbLW4FX+XrqPHxU0R2vqbspV/JzJ+027vmorXUTMZs7tvfmXhrYSsala
jEgaWx4NEB60ufAhbgt67XVaDUbR5qJBKAIMdtmXgFHgNvzqAgN4YQI1TbxG
z4Bwlq+EogxBh64pL/frnAaBnes7E510nwK3wFWGOx9ngnjfMZRlbsAgxb0A
C45TlTcSMJYV1qU/vrS2L1VR3RGOGCLfhK7No1gO66HOjp+jfOaYOKRrvWpX
63+Wm6X7D/uXMlHTaJGpix/Vw7BVL3dILuncb+FIK59sZbaf8yX8ChtsvjUL
gSkIZzwbRTIwv1Wri/+ePrnCmXmFtSy7BnVhipgZP1NcVA2HfnOtht3I/qWF
uC7348pI3DSBY1wrcs0uHN45AX+NKgDYZYlVB1VTyPpRBCn4yjDacN2icRVf
ZJs2ZRcEx5ycMW6FuVm4drvRgpS+IFd5ViDjkLVy5gOS8lNZeAkQDXiVRccg
R7UFk8HTPAI7pBG86PW+mXH2e6kIxt/psazy0hD+o6V8R4ZyZu/ZuPdqDGga
bDcWKOoxe86M8T2Vnz7EYrbK5zM40ZZg307yWhG9yyYdeen5ihnW6kpsqcKu
v4ZX8wtwf0USSVxGr+5PokRd/f4tvZCIO5HFGFnfCkO5B0J0i26nFIb4VxK+
PUFltqAZeIdBAxE47Dx7dvBKAwbkQEWlWCxwfYxs7YqWtWQ5csQDXUPag4n4
sa1OCKM2BwSuJB502zWJCSNEVxZPIA2AJGbqRqJ/mbtt/twWT+NzgPrJd7Mo
gMEcoAMezXc8zCfVn+Z4JT5oD9YeWdVhKZjiUebxckCw/35jzH8JjOyK9S6H
0bOor8+/mOistSKsBlDJ9jyfhC8GEJh/H0QWJlqsBPO5n4erfSyCpWv7cBFC
T/s189ZBU4r9YOboCmqYA2d305t9bwC6nvlekLsVeAUGSnTANKHX6b9z6KMJ
8GbHQy4M9yVXFGMoEN5PlGvFoxS9BZXaSohLWbBk/WP74+xWraIRIneRX2E8
8RorMVJIiKR1aFEB6jrupnd8CWQ8FO2RyzGr87bskZRDy13iT6B7Vp6Rer2H
GgbhoBighEJAv7jbXWwKO0lnv2x9xUudUC1S/FCiuIISrnBWd11GXrHmSKH1
6sZ2RrsIzG9ODfNskVMJ/DQRSpfFzV/egpXVyHoyJAU/WoKvOhgBayEHrECP
vE/slUcjUGHcRT0xH/olgKrQoBFjOGSw8vKKDPinFCkAi4UfsgqiR8qMy8TO
0RFGQ7vz+1pNbHz1c+eq0CpCjvHEwMdEDv4+iWzwtxoAkNv/oxDledHfoPva
WNlj86e1d8yVNCr9HqLWK67kLnGrnYYkk60R0JxCfdmxE4Lk9LDVXQ/iyke5
MzfrtYrDYxtG4/7GdVS/8TPzfx9Memdel4pIcNqw70OhTwh4LSNLTO4siUCe
RrcnfSAytdc85NvY5Rhx8wDsWX51WcEwZfGlRj6OLZwsE5PYZqsu+ZNL62gd
4VrVJPNGj0JHoKZVcCflBrSWUu63QHgatrDio1LSqqJboNHJhZIR38iUfJxz
CEkPPAnya0pWoRNb8MYVoUr2FkpqJnvRpcxj/FZQHS+mB7pM8Xxcjoyt5Q/y
xYH8E+TyxhIn8Hb3IUZT55eF2E1UwYQm4zKRkM58Ou2zWQtb4f8W0ECWVBTD
UECbtHlEyVoHgvd7psnSh+Nf9q+TbjsRCwk3viG/v3ipxBPzxwXFXIJObyQg
QPcJaBGsYtbTihpUFESvPgyIuFqs8bw4PrZSPXa8mMLUEQ0xklUs4dN9T4sj
qKLu/QAaGsuCE9pkq0gzpjAWhpIZGJR+QNxhiqFPfMJ3T1N9gYVyDiZ3NOhW
5kK8g7LRG/a3EVRmsMhBSIiQuoDkCsYFoQBSm4oLkkjhLkdGwPXpJuf3UDWF
VeIA0bRWunIlJkPz/I3iScH/UIEIi2WdA/7C8uC+Y5aJ2dIJvXBRlqLipAPK
5S/2mse9TZTgNpoX3Chb16571DNTSXuxRwY54f1RiA9TZ0cygth6agj9ydz6
qynKZLxFo4uQ8OIRbxilIsP/XdXOi8kfyiBaJw5tCZlNSIEMnUEWZg7bm3Os
whvEpW44OpxnPyZH0WLvoSJTC/IsGDyKP1I8HIXp1TukiwVfiWafeTNnFjHx
bq9bsgeR/2tddmBFpiHfVfTkbDUw4x+HiDw1ftrZqnsCWs+BitzEU2Dguc4a
T890z6auFiEKIsNuFIrc568lOlYNYjX3qRcb2ti8PpQjXSqXFvVz7erXNRZK
WaIV2PwO1rMdJUPjB/ct/VYDW4tp04Ac8AvL2mgMdfEtEY/XL7Kul+hYkzd/
oseF5eMSJTYpGuxTmIPUG56eTC5YfTt3tEHN9ifxWm1dG+k+af2o3ht4ECH4
ineLdVjzY8vj/4M2CeRo3aeB/nfgchInzND5NlgI8vhBoZ0YUJO7hPpdoWsR
q/2Ubix5693x9dWEHbtbx6NPTGV5wddfzGxRJILNkWuxK5V3gKGmfC+u0b7m
snYnDS/IDuDlIMWIFA10/8Jv8SGT1rIYL0VCC4cVrya2RJRnZZFRZQJRoZIS
Ne9XlRh/oN4rGjskSX7L3Z7eGreIhKS8RZ/9uj5GTKDFEtQzOA0psSLAInRO
dD/M/xzarqVm33S0YMu5I+HoJVPUcfj2P9IILi8uFy4uZzBx+y6mSJIQyLXP
zGdmYW+zrCSZ+XOFa7gWSFYyQo1ey+h3Zu5Dqjjdk0ozK0Xs6FgVouLycaP3
wEI7gPYPs1LUMExE6Dx9BUX9Hf3o/5BErrBo7rdE8kMHBMVFKI4KQ8C4Zc/a
ItrgxDh+pSa69PYnqrpnacKoTX5EStr8fymWXncnwl+jGmLb9O/PEi8AH2wY
Vg4/vZ8kxIql6vHX4bhPw8ZZ02oYdbQUU/7BOpKz/05Jl2ffzhnRv1KmMWzD
uH3Erxb8I68D3cuG/MmDJ5H3Qc0nR1HgHRCyDJqfXc1Sj+NxVov6ssCCwyGd
ZrSrWdX2UVp9cSHsDjpaBlEp17putQrZsyOkPfxYp5Z0deWbijrW+OjziB9/
upbWLJ5JVpqjBaeqJutL/2DY/EhHMGi4QAN9zw3FfRfjdjPEq7VP0vu4a1QX
JvpVqvO89G10VmXCygAdoldJRfJMB/dMivSiCLPgsiQgSMvJmwoaBkNUnDBP
CflUpZVBkgzwsQZeiux4KULQgCYrfU/K+psx2G30LL9GOv242rhkCg39oAde
WPQ3WXZDKQ+OeRBj9s5OSi0uEXBZvf2TjpklrigmsGbTVEdwo8c3W0rDRCeu
DMNwhX/RJVVY5brQm3tIPFTBqzCCzUk+tGidGz8ydaDxbHTShYRoauKV6GBb
2odbO/SR9XvHn0y4jlDZ9u5xqxBesRQ8PflSCfvpmsW1vk5Gi6S1nPS5AzmP
GS1ieqfe98hueWpWtM78FIdrKjgrmRVmE3Y8c5Z7cl+4uMEERVjH0WD6uW5v
caoWp4C1ui5Xeav0cItkIWhAv2rUCVzwxu1HC7lluYsZRdL/5zagDk+uV2NL
tTewkGNTY2YL2Zw9qztzgzJdCg7WCjwa/gPl1/UZfpB1ciHI+hT/Hl/vAdXH
lLZYm7uR4y5lFC1F8eidr7UkWLyXb92rgHyDP/NP8iQQilLBK1rjDrMvSeYp
rJcJ2/vIF5m2RyO8h3tcrq/dITcApAIU5VexujeBUzIe7vDl8E7LH9z27Cmf
QiiJHBQaSI/Dzzj0EVDPY/1yBz9B4yfcmsGrE9V2pgiTj5CmRcw+n8bMPvei
wR/fb96YTGg8N1vrDV1LOIC6dOpRZPwFCM99aNu7P0LrE2ca+n0BMdSc7pXp
TxZiirIkK3KYs+DLSMGO7BZCM7yWtBhGnXUpMSPmRZjoBEjYwGparI4y95mf
+iSW6eJv3XFRhL17O92r4PbdgFLIsVYxqMpFfFFVaObwbDH6bLbjPGZ+C8Lb
0IFYztCLl5CtDZfzjkG2zRpPQQnkVUxUO9CQIBVxPEfZNgR/DMIW0OecluFw
3ShEzCptoOZ8ZmQjjAbLShm2PedAqOjjCttnakrphAQHin+c025l45D1cZ41
wFM3MgmaYP4ppg+MUUW+uHHlF3TNDGnkIAIp1iu+UkOxvnzgatJlz6YYRBLi
muzNOxYfXWFyzu28wqPqrybplJAE1CysoS8OkDQ8bsF9qzNEIpxXWNNZEQJW
v8FntQ9eZTSHGl4WKjdaj/23XmeQm7JTfhoDNU0dZ1V1bbJ+TC69Iq3uFvav
mfjsKy8bPEta0XNgArDFDiGv6xO6pO2irhshXizXjLeTfCQc3Y+z2p8IvROE
QNUDB5JXRAR2iGKQSsQOBf0G/KKtgL89LBigIpKitqeK6AaDZcaFkP8JSWPP
NcCX2hf/0LWxWwuE2J7iBTW+91DUHCfz3adZw51MCvdPbt4PWCA5HKHopTAN
yjLtaxm3KM9mXavy2Alk7Gp4klMZzxqhm2LNyoifU38bt2KbM7/0EjnddntY
T1X5KugnLcvht0SWkQ77CP3hgYzLcB+zMAKl2T3I7yBWQyt+O8axbrKcN63k
nDwRk8q/Z3EcPXaWcWOqi3HxsXeGmzSaKFnYIlOHkBfz5NjLmTG2ddRCpEq7
JY7TbimD80vJvY0zP8UZUzIimi6qQcvVm5+ADJxyaJdo8oSRH4bBI8WOKFWR
/DjQ96GsEbD0hRBflji7zNQnfjOH2EF8oJWyUxjHyMr3ywjsDXB1xzm2YBmM
xyysMRP5cvFnosekTyp0sD4wTdgv9L2fjXeOpQwSR0eQXfriitRc6oneJpb6
671CrfQp3eIWwnkfnZqeo0ISMbp4kWkoZyZDZy5cPwureD0CDECL5+EcDAEp
bCL197o/cyz0Pzs4m38kNutzywp0DHN+44/z9gS0q6EiZQah9q7Pps8bWiFK
00kHZEX4PzsWTdmDIr3ABbvzu1PsxrrhpDbQxRVCIGY7qPr8V8y1wHZFSu18
DU4Wb+SGExmMoD0sbyPYFUGNH9pe5y/xwMVbdrX3lAsUCIrs1bxrqzF6r8Tq
j85nkVb5xGhtM02qjDu+8po60rmU7PSyMoNaht5YSpL8kh18G+fi/nFLL3Wy
xPzSFT/aQ3TyRo0KwxuovAOElPFXeu/WiyBuQimMhOONjLxTaBOfpnbITf93
DIWLMlXGEAgMdrmV73ktdMZ8dNKB1dGLjKO/WR8cbvR0ENRvSWKr7U3fFxrW
MjLZBMN/hZxcwcXTE27a7F7Ni7KkLXkmkhbNhqfA1d6NULzat/hRGBLfQQxo
Dr2fN3cBJxA1gOLckcrB5hWVqmictQnitUpdPID1AYTsowRLGT3up4kJyo5D
9ZPAjRQKTfj+Qdsp0mtaw8Sl63bl5B0Fm2f7hMn+Qgv2VgVWiakzab2hpd+p
9w0Z4oEfjT/Wv2EM6YIZZEnFMSHCK0Qj6o0+PN29HlFXy2kSY2B8drfWjBKX
vfagaYTWoGFZPK6cZXk7gmpd46cwLJTWkBpEm91TEWu1umCqgN3uhDZ5oZ+V
H9JrJr4I4Qb/uqb/j3yMoQNh8a2iJjb+w+IwRY0QmcQYQHiQzxvmRrPDQC5R
meajeYq9pT2pvUWwjbuWICKrW+jDxKe4vbX1v7Gm8oh5sfIbD4FskXSwfUEd
lD++gKB1IXHerNngBqQosv3HA3CWPCrb8KvY3unqQdrsiYjnQCPDbSO2/8JS
e+jnTCzg5qKfmvV5VB1q7oTwEvrpEe5ZKUaKNd6G3WzdmNfgzEC0yAloXIKT
mhBz/qB5tkf2SFPo8iqSlLIIkW+6PB/O4x1XXvnZEJqcQGQlOHR4vCCRBezI
qi91m+feLbKK/Dw2fv/jvBUrPD6rjpWPdVUyo7S5ARAL7aBgPPba8jypfTOS
YAudXwdBtYxm3UMP0q+SeCf/hisNrQy9IkHV986bOeBwUS/yJt3QAgAIJMZy
CsPU4atCzXsW+EoEzp6/wWTXdy5jIR8t+g+xG4SZTHAxUz41h/P621awUbyJ
bQ0Paji+9VFjHyKhexjld2TDKioWn8en2lLdjOA7WT6byG2/pJ63ycmUCWik
jK5W5hNAQ5DSzpxu+qn7GALKPxGBXgFL3031b06vK5ESHz6SwAPn4v+DHCzQ
hN1sboDP29R1pVuDiUQ/wt3jNPKq+uet2Ch2DffokWlOWeoTie8PO6hdjzME
hQ1oFaDTrA5JY80HzW19ADEr+ssFV1g7tpjhdBYLjrTqVAILN+kfW85I3qZ2
DQTWeW6gEALs0VAM1o4BaWTjlyGPsfyLqp6zdojhitliIcX08U1Ge2t52RZW
+QixCp4pdL8BW4v0XY66Y0VpstVX/83xURnCcN7QRCUbKflp64AXy0/552FF
dFaFv78ND6snASJFlQKjMghvbQv08SJuT3p5CyHZwesIcJriPEd51CaRrrqu
7ulMs9ZmX4mnaOleSg8TJU1b1bmUNbHScJq0dhhBlm9p7UZ7+6N3Pouzanob
FMWzlYPRwwcXHJGGnaWpS8+DjdmPKVm0h6YnPKYCYh3mVe3A2oVfB9i5uzc1
5Lav9VnmMmk470LCTZOSxRGviDzRVWML2lUwE+8Kq3zYKhe2Aa7LBUYO7wyt
yWsB6Fv+xSMs+Bk7cDEAXZEHaj2UHCsNve3rXhal8Sh1wqzc2C9mbq10dzl6
a23SyegJ+DQI1eWTmAy7zcYnG7CV9hHrs4QCcLuj35sljCnI4cK4iUnWOQUc
ofxL8JnHwF1nXksXl6SECnvLjONVRibDjhvnkFVjHnDHmbKgiWlBj3DFCinE
FhSVyOOwMl52rHlEhMaAgXWQoCnaAgr+xqkyFugKdi+3Zs/vKSvFXX5mK/8l
kaRZs7w4ouMUuBS8dv6YTzXMqy5/SjJzx4FQ2ON/fGmbEjs1VuhEkw4jf6aS
7bZk5G9E0Krr0NLk2EQApyIMB6kqLH73WZvxTd4lOifgQ5BTknAr1Tr37VdV
kNbxA022o6T/Bry4EsqKO09ykL1Sfk3E2xPoLTC9Z3nNbXHVpIkqYc8c0q/+
9oODmMBMZMZ/oIFIeP1ZWdJV9i9y6BDwZ+/VXou0K/4dm+lZe+kRDdIBP47r
nLekJZgj1zO8uDhwlintJ/hpkeplzJlq/twj1acAGWLSNoCF9Gwyk0MNzmp5
V1h9HKCEMeXcmU4Byo7Ey2dVpfLdlFH8xMEsCojt/8mexUlSGwgoxcXLGvGB
NtKfmOy5OZ2FYT5rWe5poK8IDxvonZfjwIEXSV0FyNhTha4wD8tNNRjTXmNc
BNX94lv66UiTEy6LBj5y2uxBme3x4eX4yWmkl18hW8shXbgEwmtV9pQRb7Ao
foZIj/E7aYcbRPT4Fkg27O70fpyJokTrw9Qu5Un5Th8QCcPgzHYZdY6Szmiv
SLS+Klk9990SxbolGUwaRaPuT3wfOOoDrhyWwfHXz0UBus2B8QekQSF+TD7u
iw0jpi/PzQokCPIXzTOdgwXWLR9PNRgfODvjIpQOYToe4yQzXPCva1JPRTu6
7LDg2PTG4QaFbFctrK1EuVDtOTBhu4+5Is+l14py4QPd7opSlC9ImH6RlFvp
r09Uw6QHhhb3iTTJSAR0sdwLpoVtS2icmAMbcqfCRvQ25fefRygj9z2P42wD
1rmblRokjQwdZfLHdl7OJqiydK+kqN7CBEqWYTdDfUWaxGk4m4niI+t5ru3b
xSesQ3cZgEAAjmcS6dBodHcH+CDsYTRli+exWbVOypOtO6WxMoe12qdpR3jt
RkW9olpBpumS9PAHkRYBgb/flQhqnh5T924fatS2G56x1dgu0FCSWF0szo0Q
UiV73nfapjVI/8DsR2pfcqma7F+E4VVO1hB3C0T+NWGeLDCtmp88mqrrptCZ
nGkbzCwOvcW8Fzb7F8yJk3IVZXcF5aJzGiW+3MbQL8E54O9tS1W30+eKjBGK
sm/eyE85pUfAloVVpT2e8cHeQHRyrSk4iV7JfHcABdNsxVGUfNdb98LgDn0O
TkMCV8XFajhIzs2+2fANCnSR52ZBAxLSReWVt5a/DzE17DjF/JUW3BATpsCr
13A4szHmhwjhts6o1/jkWjvyXrkkmJNx9BDf1mA0hzRHwOeOeefPzOGWHgcp
NqO+wn88hJt/HYg2wgBDdFn5mjfl17lddKv7XJO9NxJuDSv6QQmgEZyUDjG7
udtlHDHV/Iz1o1x+yMLG/tuTwFX07snAGZ+vNQmWM+RgWnHzPzhRgTYIoReI
1okJyQEY5OlC39UKkK5FYBGpQ4TzTQfIhRAEgxFIEhSliShtHMJsZZ67ornP
JRLQCeZwT61Cgjktspc5t77SFsHOYjGBCf9QfmYmHAZn7Fw/mf1tZYX4tJCE
AIIQh4ar4cBEX5A3Kr0NCFMTjbWnEvdXG/6KUs9TuS2fa2x1xPEQNobWRi47
rmoqAnMMh0uH67wahjfXyP2LmfS6xgAtgVsHVUf8aara5PusjWMbLIY+wuSq
7sF47Yg7Drk8PnQ6daaTu/N/SkU0tQNTI8zON4tV7o7Un2TLTBdV7eCf917C
8Vaycyy/KywZpviEZxT81TnLhzM7Xvyv2OA1DtP1yzdqq+cCJ9KBRdi6S4iW
hNtcFOUqIJjQ3idKKonBEu7OTaQRa4bVeeIxWjWdEgDJ+mMeQmQfgtFbcda9
zB2WsR/BIzE/W11HVbxnvSs551GV68QHKhkZwL0ZL3stqEOESD7AlpsU7uXm
4fhGi+OPsqQ4ssVsMLPyNeu17mtKhjI6Fh8olEV+VaANrZZ9ZcOBM2w3m6qU
w16n8ncfOI0zSD7IJelu211fKc9T3KULlDKzFp/R69wOVn8NKTNJkxyi3IJV
kDOWNcYHtyaiqfcxfMU5f+PTywoBCubGDZqDp5v4JGlGm8B/P51L00quTkGl
c5sDzXz7/kDeMl6luKdtv9SCWF3a0V6akAphqZ77AOt+2SzNKI06927xxQqQ
beadZ2wNtjZ0wJVbVBjqbhx8VsoARbpNDKUt2pNGcSKbanVlyOibtwYIh6Dz
CcqsPj/z0GWCCQ7FPrE0Nbjj8KnzTWWbucuHimDIsUr+adkEsHIllQzscBJv
E0lE+hONyz0bALK6p3uqr+lgHKBye/u8eKuxeX7kORiVOgPaXMJlqILO7Zsx
i54GeJh5sFnJUkb70Oy8VCjN6yYSaUPQvkxSnv678yDefG446VObvr7ynkCp
1Ju7x4Jx0GyH7C89fiLvyo2iCGju1x2gKuEDrbriEqmSJ0ya5nnqLe/WDn7w
2eOs81+DGfJC0sRjNXRNMKSXqU6BQnStNuqIAxopMeQ9h1lnAMdUhlJCFflq
kNhAcDfdgufef84Gc5+LGQ8O8hAyByzZUA/6xay5ZlDoG6I4Mb4gtAV01Spz
poGfOAVDdsujaPrI2pO1dH+I+HzynJ1vqKJpw+1COue8N30LS5t0fQfmhAZJ
c1KVMksrFbiLo3+etgJ/ooQB7s5uEXVqEs6urFOzOUF2MsYjOz5W7CbKAT9I
x51JCmIHPrT2x+TO36lHB0WE4uYYgry1+KvKWX5DsCiLkdH62fVuBHZreSPK
zvhKzQxEOeGp3+9Jg1QIAiDwuEffuLDzW59dG/PP2YjLWN9egphXUvTP2mLy
TSudwJZFKXNsxTbdWuXmzFqH5qcaa/W3Ra0/EHu6NfFw+/tEUwp0As8TO+lN
/O9TlCY54VNg2QKIswVzTpIt2u9/v1ki+i57UcUkGFpyVmQvmCuMsKlc/N6d
aIURCltpnuTui2K5sx3PS/j9NXSi1us7OTB0MJuMHLSWLrpAIQMZrOHsZ/KC
ws1rfj2NOJ8UZN7NNmtc4MpzQSM9jTeyfhao6CEN28kdf8ELy858kZPK8AiO
yW+fqoiMpxnobfWSeti/dFeOew2Ig3FVObEvuY9aUvykV6+Qzp95rfZ2LP6B
5rl4YTr8umRVXvYrU1Gdij3DZ+WrBCSVzmTFSd0ekBN5I5XFMMaD6/rSf7cU
SwH4Sj494DcrtiWKsUzToDnb8tAtAriQXZ7jv866USpp4+jM1iJdgATbhs72
FwVe9JBRiKrZmpFQdKxL64WCT5te4I4bjUXjzKJfXLlaOFxUQOCJjjtEEbeZ
mKiwo0AS5P5pG1QM0NsodAXrkiGDiS86GqSo9O3m3ITqp+Bja9DyB+K8N6Pv
OAKzHXxDhCPRreTX50+KpKV2xkmlOSkOXE+0HVbICYB5B8/KYsC1T9Th0PZc
sRNtnQ7mSUBSPfgVC2QM5N+5x5FAy/J3uW+zRkD/l0DYOtIdttaf8Kvj1FWz
OJ0kOE9hJ2r4UMchn0gyq5ZShMI+0ERO6fWBFLock+XJVaUyPauOxDXklGY6
yBw9lTVM+706DrBAMslrnqCobLY+riwbKL5i8njL3QjqwOE0LPX/ACQoDVnB
AisGEgaC1Qh3gElyo2OX4rdkMSUy/pSiSoxDNbQSTZFv9+cdmPMP1OX5IuvS
ZgCffnqVbX1KtUW5g7VPdJ5bG6+lmKl1y86RdwyvxvuJmywHeXLp7nIH47OG
pfSEBgED6pSwd/HS2IgFlH1Z9Pyk6sLcPIQc46193AIOu/tSaRa1O2TusxU8
VtkFxT+k3p3d6dlljnmBmphDYASo8nCZIjwWQbZmhw+m0pAguiwF1UGACWR+
B529SaDUmpp3jnbLPWj1TkzHmVTtVBdNU/a2V1E8KwIGDkv+Af1XZVl45i1Y
9Yb/c8H/5G9ysJrZSmxFXkl+7cCgWVABwrbOGWnSOHQPvf+hac6+x8/qFjBZ
GBGeY1GX37pMssQkbLsGcZyRqjLa9oDPFEAd3tpVd+fQDR3Se7qFiWo8yMqy
UQA39sqGP+9jSs59VfEVq61tqARGZB4w+fb50JxOVQ+d7aOlDFpzBHVazLkz
LPOUMcS7Sjf6nXtd9lsjJEGLrqRt9A4uqORSPwrlczzg6qmG2PQ+K2xPElqT
7Ny3jlRRvEDKZGvHTRTpgTx1Fs0fHkJ2q8wkHUj+FuBxYEzU

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+Eqrn3673P1ACJ7jtPx4zd5TDkaQ2M+qYL6QJ4dROS2PvprtKDcxnO+KiTfVbY5jm2v6GyrNYR7qrKL+hg+n26+qoldH4hOh7pBJoUsqMa1AB5GJQU/wofimMAxWr9CyJOkRSjrSggcGC9YPrcmgJ/BaKTlkx8YmX0lDpNwmrCs3qWoW6A39KPcGdwpC5oNfPzPKj0xf0YufHQDqWI1tHl4s0sM7ZV8KZbDq3oBrrFLpMu8nLEnDHJgWH/uJUHv+4vSst+zA0kbSJMY4zp5dmeDYvQzZCOhecQzE5P5If25YZijvjgIYSK5eofvFViEMYsnAI2qHCWbe8rqZtveUdZC+6bOrr0pd6ywu2Hlc87YtXCMSjWoZz4zn4FFgWEycMmH8W8SOK+x9x1eZKAVxh64gYXIqlBfRbwLsJrCHsGHPkwuTYPVmWCgVU+8mMvX3BBlTlO9zRwksf157zfvHaeHNKc6MHN8AByejv1V6/T+AChyvUUsvBPAuXSJ+J8327T46Cd19H6sk4ko6LgIqvbyHrU65I2hI79nYHB098Jab6g6NGHgdVp8xaMgUyy6Fe3Z7Nh8uHHn6gMU/Jrh2VarZXS7Y62jXfWzUbiMrYXqVFVIzx3ejknvDEv6LJQb2gb1qhlvf06CEhonviLYwZti4RLaeuXXfrdQw8+uRoNjX7xn/JIY7PMOSLiQ9XZCxo4V2wxK3k7xfxv3Zsy8N7us5IKqtH/vHoYYhBDKWJ0YSPTGfIHPqQqVG1og2kt+92U1R8Av9Woyrglpx6+wAJOPT"
`endif