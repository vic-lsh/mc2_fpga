// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KWxMogBRkHV9QY6k0BIEJq+jtnwgJfFrVATsUgYMVAFgG0mnGyAOeo/02/Xs
6fVe7uzhotA9PmRTCQdWRaoBU/1cZ4iqH2lYMzZhRutUSpG6goIWaYrrJgUf
SxY8MNs3pZffk1alZX1nBZeGeYoJvRHfkYqD7xJT+Sohj6TTkqkCJOPkkBck
EMriimt2jZ46J43Hc6TzbGgABQdAuyDiSclZcUhCp2ljYLhHSwRpEpVMIioa
5Dehbdc4IfTiROMR8oTV5TuCugQGhlJsYbk+E6LWziKg2boQOW2S8CYLCSd9
Tb+PuqeWjNYbGWoIwx2igtRtFgC2LGB8rxq0MH0FRQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cWNOXu4TkEna7iR8VeccScovDjQIfO2IXS3GZpFhu4LrwX5+mjbazrdS8kdg
yQ94+vdvFmoGrmcYaoRo/TEF7QR6LIvcGPUVfpbHqpjjzFa3Oj1IShpTHStN
FoDVw1KCHLoT9pfWelV+deARGM96uHDt0EegJQCX5B7BARv69Q/1ocKyB66G
Bk8UC50H65VFamC1a8BmzLkljTxseq9RUuV1ia5VHqpbUSrmb5mXs3Ufzp3k
3pw2LY7mvDiA9UkK7qX+a5md56igL4WiXGD7qE8g5bA+JP0GME8b0udOUYbp
bfp2FDpHcqUax6+83Q81CLpAs5J8f81tEMNL9zqCAQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rFcJa1XmM9XFHvz34H/jRE/8/wxtCx/P6WPsIbGfI5/lTsXTlng+WfOTSLDn
ZUq5yrDY/28yiSQWKI72KQTWu6Tj0vGV96o6Enaz3W+SMmJK68D292e5+Wg6
ORNkir4mjYbLx5CLjRFRr/INlX5CE9m2NSAYLAcYLumTgASra9Jss4ZzqYI0
DScwR6FVfLnaw9sig9XXJk37q+ATme4+aHP4c4nmj+CCTGDIf2OQw5B2RrC/
ms6JJGG1uNcuW4Z/ZTAogVqJ2JQmy1B8qzDi59G/hXhNF1oEJXc9ZziOMwPg
UxHh7qx9v5N5b/LcL4FInKqbEw6HrqeU/9xRQruQXg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OzvzZSBzXpMMCIcWcYu/KtgD9DlHIeiM17MougzS4oQhW+X1Ssmw+hl6Vrhr
QDcmiA9wh238O5U7xx6c8iTMVnOZV7AEYD5bLAl+fhiOBscTbI6/FO4okgrA
wNcnN/lzB8zZSstmFAwMlRDm9NWP2gHza0GwzbmyuVPDu7z11ZKDlfZ8n+X/
LFa4PPu9QO+YaozURFiaAdjwqHfsy5lYgNB96P5FGovbFYxCPVF7trzSjRhu
VSMrehbMl4m13qECd3v3cakWcZtNiuz/ZMC+WT2UumVa7Rp7qkp6u7hq6Ub8
WrUWQzhgKAGRkSCFSM5ntODKFIiNzOYBEaX/ntHNFw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
g40NKDH0uEC30AkEfNOxWRXnXWLjtesuHthLVt+bZzL/14GDDIOPrWU4MB7r
2p/DWttVJYxwcg64rKvgdgGvF5axFlVjZcOyxtXOCdcaO/Xp5CJwmt8dfvax
EWohga8O77/faLHi/lXd7vtmIQTFtMltcKbrmvsY3nqoHBWwTII=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
MqCNf4UeFbVgW/lH0DQYpRoTNv5J7+30azgQwcO5Gqw9iFPAdTY18OtWKygi
pauswJejTncFqJcWae4EwqO8Z8vnmiOIxHBIYAx6sH7l4bdaIO2idgVCjLFz
WZr3zAhGTb97Qovp9y8V+Ti1w9zgRr7jmzLFpfPN/fJCNvgJiVylAPP5IMKJ
XcHaDE3Ar7X6M/ZyrZrf5N8yQa023tVa/PBMNahLo8jIDRjdZyXCmOfUME6A
5ooeNor0ZVgPkksgllnE+rDk1aORNNTLMYS3VbraQNS48UF5d4KOQYahssRE
YFYZmZhmYb4iChD2IBucJuIZdxvQcFSJtaUavwrYFzg7L7HUoWm+nSI1XkYE
9tRGcOctG4lSfmuZ4pbTyqPYSh1MEpJr1XcXGWpe3gCTZFklxm+65IYRLIYt
E/O86NpqMrzWnN05896CwN42TnFeDKPa1h8qcWO8fA2MK32Y5a0db20KNDXN
wz/Wn5JqEV9dWRQ3O3rus15LqWZyTi1r


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Pp/jW5w95R15Y85HJF3NTlQftjiVPSB4OrOL2urKksQoBGpEVxCkYEAAFGXI
siUnGWuMLhDA+7cN46SM++YleAI8jzj7cZ+6Ux+wWWq95UcOxurOq4jYMWO7
q3U2tY0rafDwaUnvPUvkE2iKDJNolm5liERygwHCbFY9v2udLfk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qPOp0y753ik4e4QkgLmNIH0mlauVfHjhDmD24MfgAVXHL+K6X84ikgjqNm7n
agcL4Z/h+pnH0PoRsFzU0B2JcE0R/mWqu1fRQefZI38v2513q3dhi5hyqCeK
c4e8Hb5wi2+h4fJbINVcvZrOSH1WTOjZzbXOK792zQB/db0tHh4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4368)
`pragma protect data_block
3VlleV6K4XuSx+SzrhvQMSyZ6wJrE8UKQPKQPMI/HVzKC/kQfc5Rwd6MWRPY
ZfTBJBBIwN3cjUUY3hbxDrmGUomS82p3a//ZLBamYpXb9scm8B07pAa9cwfr
PVMh4rGUtygT73YaK4zePWSHM99dZa44YmyQIaL1sYIRiZe8yV2GiVFE/ABX
vJz6WIr7oTRwz8rU4+vhzZuYna7VUiWKmvCRmwnMjGBqpe+kzC/uThTp16BX
lx0AScNuLrXGHCFtQHvl96UVyNUpn76PgYEyNmOKrjTy9hxCZiHC/uNa4mve
R68U0k9wPCI5nq5KI9+6GadiHZrPIkSapMTRiuoEoEFqPXL3WNfM1rUAFKxB
MOE9Lb6RurrEOsQUWord5BYzpoTbyJhB7eFHKsWsv+s/A18aBUUcdpSdtmKo
RskzQptEImh7y62ZPOEj7RM8044Z00UJRU3QUm7fcbCGxyeQ+0GRh85wvj47
6G1fNhulP7b5LG6eNIOknORrfGEA6Ll9icJWWyBnu0queKZupMwAeFnTKzyp
qxfsLlx3i2AmdwIRqZwGprFXfQei+0rSjbEGbBpni0LScJAlabXrPU9jWAYw
qBsJQ8HM7P+copfaldr1yzv0OthecmrBh4B5v3HOpVjZM5TVtfpLYGFG8nHr
NpSO4fQ5wxl4OFxeYeTnoftjSnTb9+k4XFoc+UMGEm9ensS5DlCvbqhtkNZv
OGiSgdxqCERkvpQwjOdECYthjelf6WwnHRtnMaWj+8tg0N8bmJrH4N/qg8A7
C3z2JTTVs48uvkzbewzk2FD3ozk7OlstCKwCmXvBdO7v/L2IXhN9/0vef0fb
3r/oz7qQPGANmEIpwhKnRksAHM3P5qIIcNhBLPXys7rwjKIsQbNupgVdwxeT
CXfwgvpp0FlXEJatcADmnxHs5pApPAbBJnZTZtD1u6wHkoK4XESx78zBz+pE
aFz/iVyNRCPagy3vqGttEB9qvzM7uhgm78YT8EnriQgfiJYfjPrbPQSCk/qG
LWVg1EFx0lkNKSMSG+kobgqzdPJoX7NJZUdodz6fmcIOrHrx2kYywpcgGjn/
GB8nfPIvbjxg4ZWHI19r+KMB9fvUMy/Kf2+PGagaazqr7ooxdxxJq8uWVcht
Slnkb7qfAWL6FrkJE+ls1HFmZuw9IGxJaWOmtE7rvJcB9SPMYAeCfUM1zSkL
/fES8UQ7k2lCeaMOA0SuwT1brJv55iCAZGWAiD5WvWCVOAq1Fd8WXoWC66D9
GVGYYcRNhG2FDmbpswSAfGTbAvkg9rNkDYj8bIzFe6Pbu+WTPfi3kpW0+3oi
nE61nylJrOYB7BBmQ2FmGo9OmCS+jgaMD8ykHhKw2axVb0V/ROQDIp5CYfiq
zleyXnTJG8Hz0zkjd1MjbklcQ139TLIFuKC7ZWhZ3IhNFF0NRi6vu64OMnao
gt6B4eU9/ABYKe05b9vONhY17DFPd9aS1EoyTPp5zAU2cfveuT4qyn35yPWB
bbgMVrGABF/fQz5aYddLJzjyH90GKS0ggKnZpNud/jLkR+uUiRNebaXkOHFY
KRP/JOMaLoNB755tDd6dUTPYJjlK+fRgfCMkXj4XILEHD9oH099gt1Q15IMI
Z7vToIbTkxOU1zYaM6PMGLWEVT77Qvne/MxpX7Vzxmirjr4BkSsFSgth/nCn
OTWEmi5LhaXKZWscdMjkJS0EDlvuwu2uvqx7b7J8mkMXu+Cuod4Je2sPevu6
gHipxDztKRf2fcaetNF1tm42wpmG0kNyNs3iMEO8jaP3elM6Sw7jn/D568IA
bZms2iXNyilr1fLr2MwEzaWXsL9/91rFQk6qHe3viP+b9higuCbAI87hRl4J
EjVjDYd9uBFPf6qw4eKpKXc3oI7JITF33MjPdEev4Kpxo6iGV3zGe5PNVPlg
QMxN2FKX5BmC5zH6p/mhuVbvLg/G8B6zuEvEABCwB5UB7oHCchfUF1aOU3o8
36wj2zWr7g6C0yzP80IB6Edqq/vcQEjj9I6HUlDRLaA2of0mfh+mKh1BQpV1
DLt0xSUmD10xJCUi3TgKgyvwIzs/sUAFv//yMXQkfNNvEt2amH8JtEaX4TSB
XCCcCYjpiuiMLqGBoBBJtSs2pMMvE750bTm2xLBUbFzRwoGJR6By58779rsH
g3ViKv2+1otw7qMumjxBo8Dw4TNvBs/9apUy2DwCQa8zmnUL13wUUtp7fA9D
22I5F/6F1r1SUV0Sb+Q73xl/oCnSgIaDAm6+5MMWZ1C/B5hSyXUgLeDBPHBF
ZJ7AsSiRYgDnNULyMkEZortYeO7whReWjKnF1dQrZQJb24jJH3ppqlMfyPIF
8F6X3zOvRD6I4VWUhiJCCFOanCJynJpJxj16ECYn+QRnEP7aZ2OpBbuszcQI
DhfNQTgD/43coG96U2K55IlY/oxSCJZ4ZGV7W9O9TNbD+UCCVObZA48aIKKK
GdxHkrhSD8wOiMKX/FzLaUoEoSSxRH0e2qzg7wb9mVUBy2Mb4rSggoVsOdD4
Xl41J6qfWV5FH3tWYdtIYVtcilfD6bJ7n3uAQvJDlgNwf3bobpq7LpKRdt4f
uK2Mp098+I6oSUGZzxzwZpdjKEQ2HsQKDq4Cgxt4dddtLf9dEq4V4ac6MJZr
X2ox8F/8CMYToQxqNUHP7kXLIGIyQEP7f1CHCqEFzmtW4SLkUHSTt49/ng4I
QMxfGveJ0pfxflr4HaVx30IxdJIGZFZ75jU9Tpz6lbG6+B/Of1Yz+9sx+K4k
jRyycLY6AhlumdsgdyT93T9Q+R+Yp+CvkMWqPGceAdgG71YNr0vLZ6sEqD11
llX/xoOftAIDLJ1sBC/2sTTr8lR6XOmsLl8UY/s3S44kXKDZIiUthqyF60KZ
xXqxpDrbiZBYQBxG1QqZtjC89g8ciGQtlXbTq9qdGd/2yNH0IHbqGD/WcW+d
mzOw2ndlVFWd2KojExS1XoiT368zLB/4tBjZFcd/+IDFNQM7SVy8cRJj+5IW
ohlyOC9t44UJ13wcIoNV1/tO+aI9T1CwsGP1bcVOEZajNxhGJwfTmzBtY8k8
8tO+HVw3Q+iF4bd8nnel3vSskId83BazZPN436JrlVvoM/QpWewzg56omkpQ
m56TE11LukIAvPL9J1l6w1TS5+q5vq86qzSbeCopSLqxwRXSOzs/crwu5bT8
ZSc3NTQ13YDDIXpYd33NrPbrsJSvtlja3z9mlwUCrSgOgPQMNDMijn+hDJv2
mppz/2kTFt7QSivg7XZT/LqjqvT9Yv5eqSE5GOUiXWGORSYAWnf8R+Oq+vXm
Xy8mkhAclo2get/uxqqZalQAUIk3MYdW8HnctBrjhpXAh+G3e99Y1cn1dPvi
OCukL7DttDigigwX1f2RhQYMG2gQM/9528VLTbv5EH6fnDaX0ehXEg0iU7HQ
AWJ2+7Ravoo1JBePB3NNaUAD/KCSrKzMwT1B30CA3F3DV0cMv7GgGk8CD2XJ
0hmARHHo4A4sBSGrXueQWKBWnauCBFAuBt2se3aQjdPGIIusM7V5fCG17Tz8
fQ6EBqUO48ybKGoZKzV1mEzNLW2fTgqcYs1dKqhpEDB6uD7ghvqJgYPkG0aR
glU2IZEepUAggQdX1weizABdZpJqOo67CFOGE09LUY0pyCuBrHuQUCloWCCy
jQKScWfE9BBxymJJxgXAO4bt/pRhohkBszAwf/fq4gG1+Qzhl+NaIr7Rwp+9
C2ASUQydw6XFx7AFg+/yIaBQVuUQyHMQUjBw7JU+ehcRIGycqsrXth78Texi
GMuu4+EnWnA5ZtEVzy2bIoge8szU9MxEk3RoOElesk7TS5pN+hjHV7Denfyc
rDCJPUy1avy70v+C4XyGstOmtbEawXxF74Kj2jYJt/Fdm0g2QNqX/1zxfEpi
srhu2eLG4rjy17qvhn/agvNGHAq5FNtPxZPkndMyiqkeNSRG59zEo9yi0em5
i0QCVCYATpI/BQyRTBYbfl+WspLL2YZZAbDFVz0cL2NQAYRLj5vGPCYRCs3L
pVzsvXUNtbJua09k1sAz1inu3Cu1GFI0V2WWfnawAAuxxlqUggxJBFdTF7OF
UWmYsl8sE2Jca1h2422eyYEPtkvVYKblj34rVj+gDG+hNafXNZenbg7r3DQU
xLIQMVhqGpn5eLHlMkz4ycV2eIloTrpDQfUhHjmrbmYZ+AlXDcwYfzejUn5w
ld2S2Umw+kr71RIjgR6OVWbX2sT2dGvMF8tw4bGogQxgLyjrMdFLWVfqI9XH
2TA9nQDe8+zhODeTWx14llHJ2wKJmuIg0evGz/mtYsSsbk6FyYGpqbADGvRm
BxlBHH4nBtH64M37NmMGR2u+5cSdkD42bi7h04MQLXClZg/3iuNIT05i3Uz2
xl8AySyb7VzSkGFcWeHhd1/s6DrU2kpCn620keN7nCLT/8qBhMhx8ttQNeuE
BMUXfZcz56vDwxnEJ6URA5xA/oLH7xPi2uoV56xqr3813ygLfZM0x9AK98wH
FQgq4QoFfsyrrAr1wgjV5RzudQVNRjb5oVWNtMr0m3dKKzZyWu1vTks1MrPz
pmnLqehQPxFEKM4hWuzdcQTT2/R/prEJfdEYXYwIZy40IyJVXk7V8kcVF9oF
NlpAQRxJJNBQ/iHv/TNUJo51yuG5pjFekQImeJ9K2YOdskn/eofroJyy+7IW
IHw3iXP/t8aNsqlgDmYKGP/oaj/BVgahgi/DJOy28g1HTKCvlCj9zAxVYdgv
nG91UfH0pYgYXH+L+VUzAXxJrTVxzEfpuK70T40+1SuggEPitx/nhWMcm37K
IwioJsFdhppuFW3rImoafOXSx5A2Hb//qD6m6Okg2NXZsqgLPxEREuk5NDCZ
kalkkAiksIA+hvnWjVaJlpk6bAzrb3OqFhGar5qfdkeAwG4OYCJ2FBc1WhkY
FO1g7MlahkJKYi3wHnalFR88U03Tj8I1ttDzgM5NG+OWzdoEPL2GuQHlWLWn
38tRBc4M6+fWOKp3x1vwDtmSCBaqo19ZWxbKoP90unr07jBgNBJiVKgCg6Qf
PvTxuMosvRl83AWuwMXc2csbYwdJr1+ly2j5yghi+YIura6ONrctTNBIa1Ih
bVjEwFEVjpg/YcAu1J3Js8pccSoRSX1qSIX+fkw3agNlkjIf+9Jxut5rOL3R
Z+dHHCXk/X0skfZsnx7XgN3EwBdpqWbGBOWXGYyYOz07mihE+sBes87Bpxiv
fFPI6s0BqCrPO54W0i8+3mar5tP0FBhFfzo/G65EUJhYxuQr5QRMV2d0igFk
HSeBh7BVyL+G3gc2ym3ZBtKkWDcsinYomBCc67aH246Tlvh23kI8J72giH+H
APMciqMzDxUFBqeSytbGJNBQ0qfUty5PKUPWK4OXqR8v05efPPahxD+eUjbj
pPD34VvwrBz0jX/+gca3vhcHC9LKlSa4tRds9CAAUCeKUBYTcGSjDb55rOwl
t09lM/iRlcCUKpF67JJ+FFDwGH/zp44aCxhTaYh8E5F6DP8yKl1f2zYRZs2a
qJRHSyp+W+6Yr0HR4Dcfj5RkdFBt7noNg10Tw9uPPGvidpKYsjd+TMxy0WTP
aLkrEJKy3C9gBSaYu5gCQAo0zU837fsOVfXtyG0zMPe++rg9W3RrPof+RURd
EM3EsBmqDm1lYncvL+/z9hOHfe6CBF6Vhx8hTSXRdlmLBBxEOAVeel5LpCh3
n7oly5FDmYgMUH4rgURd8fktyObztEagN9Z8NzZMAKylP0UdbZQa2NN0bWMy
/xuiatnBoYMO5drZrjlpsi4FBOG5X20PIEmP8A7bPz+am5flDi17XADKaBFu
HwgI

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyIJETCcZMh6YEmVUSvSoLnTDguCqb996Tc3YKGlzPmd/6E4J0Rrm3xMc84tyIrxj/camZMkMls8pEQhbyATy+gbYtav1UYy/Tj4yulBWwYDYMXrBEh81HVlbGnU94IslA+cdBUrJeNunWqqkU4X3Xyx6ZwwBNAnN9Y/dafVDtp0w2XWdAKvr1nd20he6K9IhdKR5qV0iHjtkRWyQbN9vjWwEMWsfhbyQXP3773Ot6JdSQTBhkCMlZ10+zhaRzy7xSyGuZ9jQ/MfM+j8wxe1QkkXYl/IPXWdaua7oamaUhE8FW/1Cero/CHmheLeJATPkR18PAKMOMhpEp8ITo3xNiwJJ4pIPq6LCDRhlG2no+YcoIpmyx+NawsM73YPYM7OpZY7MwnXtT+HyGHseL5pTh+5l8BAghsPSteNICJ2dlXs8R8SikJeCjmrQ9CejLPL4zQFXYYuYvBdOmiVSAeavjT+xoIH1QqHnwL1AmqWDIwt6kgmaV7Pg72aFmRISNawh5xL8DP6UExvssofu/hJU53gmwNMm7ZhOs3jZIldVA/Unto5rfnv0bruGryJCueg6HYNO7ZyJu9fKstf6kGKCg5HET1Huoiv8vhd27XYduB7lIkX+r7P4aNQnlmShqeXSNYXacgRz1G/DEq7uZtku13rfRft7YEfJv1/8+HMJbNVgCVFvHxhq36hz1LSlEyGDF+lqtMLQB9/l9upXCSblUmXs/Q2lUt7MZut5VLRsRT06CEOnF6OEeZVXM4djdnHijPOGxGizgF8VgFCKmjOQDEc"
`endif