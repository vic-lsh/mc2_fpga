// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BcZJOCrJhemYbSou0fsjE8YlNQQOKqHx9GdunCvpm+OIZ1pE9DZO8JKiuco+
JMsUYIIj2om/EMBfx1av70Ruvv+yBwXmTTXV3Z1Yc1eF62GB5UMyTsdiXXrg
ev/R/5s8pRCL3VNKcAgRay0LzcXrifizCBzM712iTAb96i6I1rKabi5xV3bf
2BnvH5HaI8vzjzg0S8NUzjxwCrwPMaTUgzdOnPal8GkJihK/gteUb1le3w7P
c4QsVM5+0aYDqkzBT4muCQmbF4av5m8Qc8RTwZOfxw5+2K6RJgPiToKBXCzq
QL7MOpqaWIigYbXT4zgF/wTuaTyNRionyHuajVfLmQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mndzUPwNriMsQexMzu6IqrLqcNkuErfpkwCE4YnskPbJVEPev4/GdeAXlcGb
RFJuLQqlc9W+HLXmwgDWp4+1Au1FpAeqA627ANR0txEM1T/IFTcGJn6G7W6S
bl9AaVktavwqFVtypCZ5As71E7GeZZtnmjKXFhyB/ivGOgR7J4uPnNC6F+j+
ZH4h6dlsZML3DFP+3Ihw3UyQrJTs3GztebUrB7HAv9OFXjgdAYq+/srHyz8T
ZVMuHsNWQYxfFbv29leuVp18T1sKYkvCekaY5UQWsvy4ZJUmfrlporLvJpgW
n6WMIlN06QaHFg5zIxpD5OxIJqwgIb5DmEJcBXq2wg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Xelq+1nuuHpfaqyOl3OaP2mpGlmb8BiuQTX8iE0rFiyiPcR4JMYWEu0crnkH
FRAXpuJlRHwzXqGGeOHEzsOuUm3vlyWmNuVsyWQ8mPezEG6kj0EluaLfyxhC
ocBA4lXNxZy0hDsk0/nntY3PvUxxJQu2QUv/WzIXttDU6Xz7E3Alg12nwdTt
/oou9wlbZ/vYwlRToCrZ3QUzY/ESp7xG5CWokmXk0y3SsOnDVT2AzkaL3kfl
aVmyIdBH4pKYYo9XWKFlE2xqxgEnbvQmqi+2d3Xt0TWaYgRrSr+OOvBtObf7
KxPqDrLMcQ7a90U9SLtymMmm+UG3nGYvMAMB4mVPhg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
acRgh9ZLdjLWKZfLWhjiQJFKX0P3HbRgzz/57Si5kV41GmbyWXbX7pejkun6
nO+XCE34fP020jGZm/LlE//ruugS749WuUbnTdHlwm6ol/SzlA9oKvkWpniz
oEfRgetNiYCjmsk4ZFCVvH/+lhx0ppDqMGEeCuqoQnSG5XW0AGMG9xmZd/NH
eBN2VF447SPrN3zms0+Iinou4PGTFgHsGXub/us7S1L9x0u8Hv2ZCHfNsyio
/xhyIRj6vxGpUrO1XT68X6mfDh0va8HuqAiMgGGlN38zbOTKTvlSfRZm15MA
HDMp/Ka6Cn27stOmcuqMRHBaZlrng3AqfDF7pI5ljA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dGMwM1i56kaXntAYslP/StTejizoxjqQMWZ/oDelcpMSfCqmMn1kijybg4Zz
S4TG7P2qGEqiQGefBteCueXn7h6gQrCQYyOuWLN5KsTRIvfsgKVvgdJL0Kfo
MyFM4ZOVyQsNzObyIYTYxT1fItz3RZG0rGyW7EP3SCFzDSqwOWw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
T/hJ3DVyycrbwpx02nm11Ms29T/1r5JMfC1ycO9xEiXC7KACiw00g5eLQq0X
ZnUR/CidvxBIIUHM4DvJXqEJp2e8pYKUKaEhl5+sKYy5t5yF/4RuSmSPEvwu
K7xx77oeuSN0aD1q8cdobA7Qmy6HvYov3MjUW2h46FNCr3+q2Od9DW5GKx85
hTGyhoGAIZBvluGZ4QTUUbGD2japbjz/uOyJaueiMW8J1vAqSILXIRqHRQbP
i1Xf99c0NwsOh8rsmWmnN86tX0sypcqxO1YhOLfefD9hoVttAuumW+/bqtA4
K5dEftoVoD5cCySILqTBbsyfO+xtL9UD1eE+SE5N7U5JiMjeJVaC9n4x5UBm
wjJBTZIGJDbKTAlgPQOeesUHYu+wFpoLV/H98lsV9Bb+bd+54S9N2L1Z+Nu8
XamI1xRxPyyetFeedjT4QXRCUko+sjr5+LMZdfdisFzuVctVv83ZL75B1QTw
tOZE4LYSX40f7UYXGJPR9yXjBiOj4pQw


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PsXTIDrStPfqT4ip4uR6EWAuGMT4q6wd99rlG1ujjtofrdHJjiAIgQnfTXIZ
1/ypH8HACZ9MBSq08OyO30T1RjDE/GpMgbrmBRlMsIE9pnsJr8CTYzVYXNY1
9luzJdE9V8Dg/epY6h6+N+RZcep33wf/0VQMCbzo/f8H5LPRXmc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Pe43WIoxhyvBiC2QepFp/xIbvbvWHBjGoIe0f64HH/r49BOVLze3gwx3FDvz
XE3l1U7Wkd+W55VMlx/kHStvjgYSFwbnW58tX6wHjwzdpVCQxg418H7Zp9v7
K3zz2igMvL67ddlY413mQzh4b2m6/Wjoar0NW8dcapcLzz9SkDo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13040)
`pragma protect data_block
TttoKEw7DVbCjjfsIQDVZfnYvj9MtuhxHAwP9W3RpxMC9K92FIKQN/gDliu/
gzmpU5MemEO0A417KadE7KOYQdW2ZHA7Hba3OCxbRloyZypII3WGsBTOBVWv
2eo74oLNkmWnLoIXCf+Ou0Ow/vW9XeYino+mDlFqqqXQ5P3t9SkpiAfgEu11
DuZkR0DGH6mxLx1nDTETPSFQVpnehixeof+S+/dcO4n1OHWQ9Ng8/jxwDIGL
dd83/0qvkx8TFZ8fFzsHQ0c5Fcpxly81QARh7TB4t9NQOgeQBRvqXX2UOkO4
KAg97WFxE15+oc3GAUhFc4mLCXT2LnpD7zAyvJ1lr4goD8hQPqh1QkOgmYQY
bhX5HTavut+1B0+pONdEK098/ymaAN/g5mgG3dtxQmMeh5BVkykpizutE26E
t9w34HPmzTcmnX2bKL7mBJQ6IFet3q8Xznx0Znqy0+KzVTHc4xUZlT4lU3YH
ZK0ywxrSD1yvcC1gKXPdrAv8vMMRp70AX1p50wIdRThTxjIMyin3wbObxNXO
9vu2Mo8ILJT6TZm+R4aVq5DPka4LCgBTy59GvnPiftpA+wRJjUcVR8aMQ3xl
08WtISufa1j5oq0M2bbr6W7pZ4yNt5wrqihjBJuKod9ov6NQHJLyI+DuyxW7
ECXpm1MmWPExIhYHyuEMdpR/+EqQRkxR2gWjKw/tCFoOVQWHJmaJCqkyuR2Q
LZiPvF9oRYW7Y2+zSUb/QKE64BIkGtZwAiBEmhi3U1zBAfoNUzdhfz5freld
EzsMQBo8Uj94ZEijT+giHUQuEuSKmbQ/C6AHY9op/7/Gn5zY1s6zXsdeYKdS
vgwyVxWCxe1wapdq6vS0Lea03pAGlbiKxb3bfWjQHC6kBGVCW6c43n1wTYWy
YKTO+lAHugvUeNruqaaFev7tSbJYESvzuEjTR6jr4jxDUtEqCy2uJA71s0Km
deiB/UY9v/viKdEi3jlKj4BPW82W0DfVqawYTUXUJKV7fzHXodcM8M1DYcTq
KxL1UwhrZLydgiyNYtD++VOPwTM/x6geKmGzM3XLtIOzNZ0HXjcs6sUhj+Rg
NbUdx4Xypwr9LUItgsvbyUwvdiJ2uyAEJ1IT8J6bxiZtdFX2hB5Sw13oYnR2
UZLqMJpTJFPqU/tqi1KX4/tzvJ1XvljAgFWDgLyjFW/Vq64f/Lh8+8OYIbeX
jBFdBQUBS5rwTJDI0yBNj1TYFp5rca26TT1P0rH1BvRQD1/IEew8/TvzsN66
Ejf/YU6MNE+PMqEaJcKkTJR+rN94TGc5744zRZU5rcv6H42TdwevgiXNQxIq
kRI9RqSrmAHa0020Kw7ENwjVs6nZGkwtP6k4qXbfWJZJwqkVyiFmD5pmNo8V
fmIJYI/8ofgvqukNE1BbX5j4LNtQ2BvD6In9ygalGXbbVeHOYYarlUS6ducW
fO9pgGhxhCb0/so0Swj3Y3kSXRKOFLTLtZZUL3i68oJLPQ7Y6Cjt9/6GpkK3
3GCvbIxaKf0yOPX77zRLxJPqd1J24f+E7DngEeGomn9/mfOI/b+eONgTs1Wc
U0sJvXBNMlmzx5P+eK41A8QD56SkHFd41ZkqS0DD+eDpqx4n4creWIo1GWPO
JQAcbMq2nf1DfyaJ2hJYrS5ZJmlJirxRROwsKSDpe7Whl2CGvnK/U2gfLbqJ
MAnfvWXpzn8vbX/6lhZuPXJn9MP0PxwQYLchpPQT9sTFbemBQddixTJm+BOM
1ADMmxbb6cKiCH2a1FGa8gUKy9Kj+m9BKiFojbJBrIc5wPQaHBV9rV/8vDPs
PL6A38Hm/+M7xSBN3YO2ACV0Cq7oI1r2awgXaACbf7ZPwKNLRBpgwLBpFNf0
yIqKoHvdIwDIL33RwOxWhPATPPcfpDYSmjdmafJcP4VnqUWpXjAGlZQ6KU6e
VTVueijRibbYrHGRebiWwFkaV2M0YUJCsOGFCNYksxdJ8k68igLkpMR8XC4J
mNHSlv2Ctqf71TU60DZzGiBk3Q/NjLWBJ8dzA5rUpkwJ972b+N+u8MK8W5/5
zDYgoDp1RnIWxGJ1tIdu3D6c0I8v2MTSkqXE9v6xzp+QpE4lIRAmYc5cu37x
0QrIoEEy2Y4L3k6PDa+B2iwLaavoNfF7PFG6OHnsqRVQTocoUznkL9+ITc9Q
GikwkYMjOAsCDIrtUx1RDc0lLR9J+NMF8Tz9ioNjLGYzP4ZlgRKnZqW/xHIF
lMp2yrs/1Nri0K2i3DaPNeg0uzx6N/844FTHnusP2KrPWK3yIiUinPGoBBlQ
FjPBtebVufQERPXrWtLUsUPzEZrcoUJESbNPZB6MylT5zogmw6lO15VM94VC
vhZppp8E0WNHZMyvTp2ZtgvHg05ekyKIgl7bdZClApmc9OPuBsFtvr9E9yAT
2Kj9YI7RiXATHzMJrkTeM92qcSMsTwZnpv1yLORpmBLSyLZwT3Z6eIsupSdg
X3poZXCaMYqugG002nXGLNOPluFo/mpwQFI424/3AE2UMxo7oHI8v4Nt9sew
3/R3jWf1biQ3GKZHrOREXEd13ee2Y6NdBDZB8IyuuaZKoOJS5K2fJg54U8Ey
hlpJvLa7/pRFJYWJ1fHyKRZrlJOMCqGSRbrsBo2OvgL8aiwsO1oEuRJE4IiJ
EMXlJwWLjmLp+RE3ogwHbnp74FglSd5MU1yDYBV/JeGtlIyleYE8syLqUzwC
yyrFedyxaWJ0yl7atySvgUyPnIPK/aYWoBn/6hDK476W/TxmqMRdM3A8YfQS
PbPezIc4dgi2GLJiiLBo3yNjaPitruYEyYIByZsX6cQPtWsMUhYzxqyU6kZW
hOIHzyr5s5s8jr9n9H0oY05c521an6qN2qEXB/hwDfqFIMxOmECKu69lryBU
f4b+uUMlguXbFiHyboed/XDOyhuhP8+AnHFt91ND59m4lUOXR908H/RZZGhp
0h8LvNgRAkJAuwfuqW02swT8d2dU3YpoEu4t3KKgXF5VY5MGoF8v4mCP9oWI
VpDuqyunSSksspXrBXNVPx25YRlAEEIcnT+gqbrYZp2jcc4CiGThLWlWtIiU
HQIxs709iy525z3QMTIi28t5rm0HmnvvbMNMl4almYVS92lL1cnGynGwF90z
OnJjoK/aLBBLGndz9EiCYAcuFsDWKrQc4NEUkVPYkHkNDBigL8NrT6azJmWG
4J2p/fWLBzMlv7r1zaG0Xw0KrUS5D9B4IE0WSctj2mZQbp/H7DlCV0ZPRbti
SBwog83gWaE+mpCPGeJDVoNPOaVb0VHVImzsIredJqhCdgY6v6/PmdfsT70J
FP+4aDLDh2+lWRcCEod4s6/qQx0kqnd6urM2E1V8Xpk3K+bvIxLRqGzodpOf
lTYhuEruOyRaEheEJlQ9hz9QCOzGwDUaLjNPfBGgr04JJVuCJfHszMk87q5I
g9fVCWrP7pPyP5F7H6Tt2v9KkOiH5fGowNU1d/qJ2jPWxDAhgYlO9UFvl2Fa
ReBIHtsMtj7FyXPXIY7ryS/7qZHTLZI5hlostxpgQK3TxFds9dss90KeLkjA
euVU4QHuARRFp7BhC2wOaj9oUjWHQmfcxJjY5hR3k677eYE4Ywqi+EK3RVWP
8vL/XkdOXsjfN8YCAnLeT0ri//aBCwN9d73cr+QdJd+wOb5KG3Wioldg4hsI
Pl07VWXUaurzn9l+GvOY+GOy3u0Zr2Rgq8d+3O34d7teh4gTyCgRl5dGKXa6
6igExw0+9rSRQgXbXepLsHvCtbHL3CUET37hfOChNkaurXfVMSgglx9ZVFsb
dgwccmzY/ZzOkZmN7VMIvog0wTBIs2hbGae2b9Au7H1P1QPtdMwLkLy84LTL
kEXF5R26zU4Ajvm6WSY5z1SUpdRWi4pPBmtUVYvk/itsKCYKYKkSB8jqlmHv
dct/6iavMAg1koRANBuCcuDnkIQmapKpDI7TdRsLzfva5rs/tAv7FeSyP8F8
zHhQCioL8AWdC+m0/I48PdoX2fjKGr5nkTveBxpJlEX+hZc3Z9LsEzJRs1S5
Kj+FmBEV+5W/0yLFEItDfnYV/q2za6x28vkVMUK9kLYAOEg4SrbHjKbioEwt
9JK04YuuWZ/wTm6mOBm09gbBVZr6bVlHeLga5cy9AuO5OispbwKMj6Y/t1U5
EahGlstPdJXaUIBoySJlSElJr8t1zCW1qKdNYqjbZu+Hwr4Y092eyEYAeduG
+bugZLz5b+wjhczBBU0AVu3YEQOBFoQ+aPRrHsWMfTSbPUzOONkuKMmrr+VQ
9egfQ2e3rJ38KmmBiQyRbdNn40lX2ru0KXdh2FZpPMYDA2L9W5OAaF2ZjU6y
AHO4Aotxu2dlpm51w8tTBLhXP3HtEdhQaTscBagmrHDhE+hbWSvLA7noEJAg
UCnHTyo5rH1P3ScKipi1ELLa9z0S1UMKnC3gQlHdAq9hZ1Lgrd6pXua6o1vZ
88YmQ8XhFOo6VyZvp4LbKjPA58tqkS7Cb5VVYIo9cd988k3DcOZuMsL0a06u
i7wTTWTYz0qmd8u3p5gsPA/tUHnoy1JEVTFIWoBRIpTf7myv4UEJoUGReH1P
3mkExh+PZ3VOO2csmK2n2+Mu/tdjkSJ3sQ6vh36p2ARJEXk12ipbRRPIH6Fq
3Idz0wSbDqENqj6BjOeY/IGFkize8NJT/+gFgCrC+NjtjrJyw7EEJ0Kld8o3
CntgP9gznafbs5PVWUEaqp92wZ4Tf0sRw/e4GZj7JIh5b5BtwH6jWj75gmXm
kVHNJ9bL4aWaWn1pPFeda/Ii9DHVWDuzLHX52RhdTdLeYdD+AdTTAnwKRGkh
VvXINdaJVc3/dIszJvvpJYjhmNxMjdEFvhZ0gQtfTLLbbn5H86dY4C51eyd/
NTemZ6rLGGuomg+8cvzfm6zN65EBk2N0T3NWQbXZ9jIACY/aqZBE6FpK+5Wy
8xrVcXbVm4F4wbmx/LW6mAKZz8THQZWSmm5ngzoApK69ntVGrhzSd+NWetjG
U9fcs+ra5bVNO+FObdZfZj0FKSbdmzDBKAaDTRk/kEDsK2PNexR6fkWVz0qt
yibyqu196a9/HmEu9XgRRIeJ/OdlJhjCowkxkTvBKlN+NVDnojZ4/+qAspvI
9UGyop5YIt3x8DHu5lvSP5cZSjpP7gWn1kW3JXN1J0TOVKbLFMXG84xP0vpm
DGziSHdDuUVm5aXadvkmINz39qjBvkdruW/+biw4Uz2xFxV5QUWO/O0e4uV/
ihGTheJWNfcwvmioOVE8vUcn+oYX7H+Dh9qqCFw4retazPkgjORrX+f8V3X/
hIUck2nXxdXdg8t6lOvijyZzTCjGcF32gcVY+XRdPZUEF/OJfz7S5n9mQOVV
jVb1/TMKmvv4o5Dga0FdlDDrHOdiZ7LyHkQQNqSRL946CuVcHLZ7WUYGKiar
ckOb5GFn73ruQ4a+ixzxX9UN0AZ2vPnl+kqiy2J3CK6up+111wd+xLS5+8l1
kAGVAE1SEdmbwTaDmXN2r6jYFoB3mc2S3EN0dGjA8RBLu1JkLpPXgCVopMKw
X0Mq8AYlzjiO/fMtLLCxiUn57gh5XbN0xBf4iQVFXdX0IScSUlfX6EiYBBhq
rJ5IQBgi8wYA3qICh6xMkwr/djSIPWSMUnx+8XdjpFLd/B6zfjsWdy+rUPKe
19c4gRx/l0p8yBmob0pHWp74qlMEmmlbiFZwOp6NDRlVScckZy1NLJzyDFsg
FkH2hePWPukBbNYVf+q4kliteVECnQHnWN2/5giAOMm2ve3LFPr+izT8DjQf
tJIG1LF7woBkY74Py7pK4cs/gnHH9D2IAYC8tIw1nwsnH4RoC1IEzZk1oz4U
FxfOIBfHhXhG+fmFLlrXLR4x0VK/qxwCP+1HTZk0LIDEZqjsswPeInZcYdmP
d3oTtfRbpXEgl1IWagbYysQqMvQaVsw7aejc4AvmdOX3xLNGNfyvLNLSW7KB
th1f+oOnhWrPryxX7C6WYjmU5gP8u3F9aoJQOc5iXIo5WzxoFLuobO4W1w06
azJ5ztj8AoVDncQUgVm34YX+kpiJgcRoImf6B8hRxNzo4s4e3j6HOlZG/+NU
1KG6dAyLeNEeXB8kV3SKHNSotn4HtPU/fnPbzFShg6Vi4aIz16uirqkjfoLm
LjZudYgOuIWA4Pu+Hgzz3alh7tRfS+uXpO8XVcAbHP96KPMoD1+DlFEvXo/o
5XD3n6j+RPhMmAUt5cHsXlFO3mcEcOq/x4jfeYnsw5s3u/QCPlU5UJnoT0cA
CR0z4ilT1BXI25q14TDZb+ui3fo1iCRETO+/zi/5TXR8mQH3HzNVFQ9EYQJo
ehC+2ooUL+JGeZqYM/oekzRwLhXxTzwGychzj7Kl1DitNk1/jr4hnjon9aA2
Rv174nflVhvUYrqCBxpVFsstHRzsetDcama5QbcVlA37G+wyef9cZv6pubzL
+7XTh7/4YbdHL4AuNlbS/GpwgI7i2Tb0o4mIoBpHUciCuv1ufGWOrocG3zuh
gYOWeTu4vPzOEWOdDzgmdBBDN7yczpuk/mD1xHG6WRn0i67wmjTv9lOMvKgE
J/XaxQhs1cMGyzttR2LgN2JYWb8XmViIr1/oXq4ZftUl4jj5GMLaQH6smAuX
2wt0viJzYrm7OwZY+gBK975F92h8LgLqd6Ih6qqn7RHcLwZhPuCZXv/Bm1t2
P34e7QJJzuNhtQNzjtpzvdeXFxSXRnDxLofPFlmawHhAgEIKRuFnaIaRm4au
tJ+y8GAodprBQsx1e1MZPmrqkZ+V9auXvNET3/v8g9YfS1vjL8GMTEVVoQYT
h2fF5/uKI75BQ1A3ayZehVnum2g3zx6GgzBn/As1/pNPIJ/gBWKbRElYKd74
d6leZbuOfgcBdcrQiJjsL7uVsXodJyvOym04RlStiR2TYYBz9bMdytC/r+3t
u+rVbBlv7y4MTyWbCYFFj27VJp7NOrJL/2+qRKZWomW1i1QYdD5tretTKcdw
/Dmjbn9mG9B5MGWrJR1un/EXul0XGSUxxo3WiKKhIeyvWc0NLfcioUQzZ6s+
Xf593noxbwe5eUW6Gf2uoWlsSlA8SyYo9JmJjGJ6YtfBah53MgqkonwDY0iW
xh5ey6WTzLyyyUoVa+KlNODA/cgISpDS6fv5KJnuxQissGAcu9n6ZVDzWi+z
FuDFXAu9P/XVtZ/4iaGk2thyu+A1EEfVkYXhPuhLnZ6sJpBKRxGmPsiN4S90
AbxRqbWoc7c/CqhZOOIloD8b9g3nCtp9qyZcModPJadyZA/xHMz6H2zojju0
PvJrn2DSqWEx6uvDotR6RlwKSUD2Uqa6/nfhjHybYHyXuxVU4KM1eCQR1Agj
QYUlpbkOFzg4hc4wjOPvEi1OOoU4gzZjkV1ggOzwVcrObiOgyLn7eNsGOFyv
PBMYN5yV1a+sMbp41kyRlBtUheFI9nzdoUvMdJ11UG5//ZRAosH23CjFoJHz
pRQKnoj2U3Unsx+rvLgiAkTB7ioJjM9013rhvtwDfwnBWK4kjiEqHElAW1IN
a3L9KUvJGR9d6FrFE82K3f6DKx2n0BbcZGJ5US2K+VDA3HzHm8gpX1hIwsrA
KoE4q8s+A/QOz6kYiV6eSJTnlORbkUOaw6j7c6Afnzn55k6VYVN+iMknHv7I
hScVovBlTLH2nDR9jeVDJtX4G3/+q/9GVE6pSRdKUa7d7QtraKKqLLCzB39h
hQkwmDX9R/3HgtwB2j56kEvH0TJHIjrWZL158t0McqtsCwjtP6wUm2qBPP+J
OEaCtfMTPLuWpB6yG/0IcpQO7lgckin7EvA9tvEqr/bXMWRaxdihjsnX4lIL
JgMmQxnWWwC1EOzmT198QFE5PCDupvmbuo9ZUgvWpezIG/P8+eG12lB35zcH
m/jZmL2ztqjxAG/t0Yp2haze6uB+JGGKLrME82G2/46p7Z2VeLIF67H8EzM0
6l2hxa2kVO6U5PU8YD7T8BS+oW18La/wDN1u2/ao5JnevJGvSoV0CkDztGuX
0qU9mAajeuvH0qUaFLmxE+Pqn8kF1APFMS/aoC8hkB2CIHzRB2iRGvjUP0iH
hKN5qms9OO3XhUyS3G6P4qQ7XZCv9Mm1qq/1NbNWweiDLxv0f4/tj5LLogB2
N8cXgF3nQU4XdfVdrt6eNMDqDy+AuUtmPek8i2Bg4y5K0TgWquHGzEKxLlQq
yzuhejeTGmt6+kjwMe3OFrPsmZXdZQT6PPd9jQFWIAcWWuE/T53U06lnDZ8L
lqYK1LY9z6m4doUdFgIhQV0b+ThSjWkyx1ZHJ/6gw8mcM8RY1I4pjLxit/nN
gky7X7/kyVQcURqhOmCsgYlzqWykqwXpfaQeo6zA+bSs5SiGD9HQteSFWUGi
t9tdEUsHqN/xmme2eJ0zUQMVxw1UL9p/gN6eSWfLR6vlvE40cKwo33HZNMMD
2AM3VUWNTsSRfXkVto0yv2njEv56aN3IkWE5JYVqiL1Q+ZH5glhx7jdTwUO+
bCQdJc1ZKLbZp+d7zuD9fXJg+Fq64cGwGZ2keKDm3a3J/bnEtNoFH8QoUIH4
HThYXu/LupuV2eMpHDrG+r9NgeWLaIKrLtcGrc7uhoM7gsd9WrIXVYCk3Pa6
6l4SG+C02drll+7IKucjaDQpUURPytPyf/zfI/ou9DPkDkdsx0aNp/IXOO9f
+adI9k8b5JzsF1tDW9V44iYT7ktaoCpLKhyEyt7DhcOGVSy8bJLJ87NtGsyk
IIrzxFYIbl7nnl1HQigIXbZ0iVGLrp/OdtjdEmxWZRRvr8O4x/d/tJv8bWtO
u/uyNHdufldZsDgkHLwwx/uQUFJzFQKayOIrIB7Sd3ORTy3bRyc9ZC2vClQA
tIu0fCKOp340Y3rxcnbQyUCX75jGBprbaqiWEwGA5b2b02TpJ4w2K/JSBwa+
xBOopAJ6KCB4mx8IRGJaElgiFULs3UMIfSg4acTsVJ3JKyn9jML7M8O0qLZV
lmQpsMquPllsOTRda3blawPOu6G40T4GBZ88mrH0y4OJmzEalotuEAQvPyLl
T5yjTnMuncU43ITgVbHMW6Sy0CW5s0mSa1OrrBUPRjUz75pR8iYB6Qv6YqSo
aIDCkilDAsfGL9xaa43ZOXolyHj0eKduzc+5gwVcQnioH1nAYnE3v8pz7VGn
/dmQNfD5PBj1w3pu/Nx1G07EbKx2yTnMpokRdU+YhfVop0UKgHfXAzMpKdAm
ToouOq3AqxL9bOTpa0fAbyANfeCX0clT1hZezEbA6Fn2igy2eygqp+v6LBtQ
Mv29qvCDwAKGkdMIMdPx2vARAeUlubOKQ3VHdVhaSS5fFkReVB3yKXvaJ54n
SpBv3xkJcjAHxh5fEm5q0ih7hLG5boyiJTvBSaGhnCLdvt5Lu8IK88xcDJem
BC8fh2vZNK1qTMUgasjgV2iV6G9qaLmAruIvF/INBcxKSAYS/6MApQc9sEGL
2hcYdQTQ/rQWshpBIv2qVinHKKhilZfNWe0FN7Us4ZZaF2QnarXpNDhTlBeA
m6mzPXhibmjTrgpCvpDqnzDvRTJ5sMXhtggL/z4DFN0hOmly13zxj9wPQNHx
AlbMpAV5kG6foBcO2RKH0yKYuVSxnGrZDF+NCHhmv9G4+7DGgo7wKAjas08i
Z0Tj175OyWMrjqSBS5T1/i+Doq6qlGrGGudJuX6wlmxz563WblK/dAfp0pVk
SXbVptM3VMpNgv43LJJMU/1WMnL7ZqXBviqnQyP9i3gom7o4QfLQPw/XGrkp
zgukhGAJjvxECktMCSAEbQDhFXJnGQ8y08+JgyVxU7IckEpskJhghNkKKjG0
SEm1nW8qs1Etp15Ghebuhwukq6Zb39R2yS8R01ZUu+vjplDc81A069wlr8Y4
GZN6bWG6BHzjhOPfuN3kvJpnzWSXYdpRkGf19KMPzwnpmPifhGMUg1aoY8nG
xz/L9OW4L9d3ek5zzxq2K2BhTEzXAGjIunKFyqU/noxHn+JXnFNHYXRpTHlq
VgzSe6qe1IZDj7odTxAdB5Zk+HJAzNp0knTVIdwvSx4zuAc2fbH9tz2S2KS5
3DxaBQPyvQYGOaB2IqC4KY9Gb0x6BPiLLAOhklyxsInPWpPb4OvXYWiPVfeS
v1CH/2Vf1IRBXaFLv+pdxIqL7b2ffVdhSXZ4r0UycbzTltc1oqokDZOn82sP
genbMxaVIc4gPpUYpIW9jR26Or/cc/YFUaOTuaPt05Urfnd157cFMA8AtlMU
iT7jDb/IBu8k+gccXM1m6LaU1bRpaj+2vYNyfvz1UxpUucKBbkTVSQL0vifM
sdhzIts+IbEyw1NrhPhLK6dCWSQMeDOLLdrjB/wxvsWdn/+yKOrd8h3stzJz
EjwiOJF2IwGQ2o4Ask7NZnv15AMF08S6Ygl/TshLv4w3hWON6Mvq2/+esoXD
tV43toygZqNLtmJo4abHK2QL/A33QsrGF5WQvWyjHq277snkBbTeYj8tFy4f
cIlhUSO9/NfnciLIYTxlehu5DaGolIttFKiSIxLapj6QmU3ruLXLZkM+yx08
q8/Zd2/SGS4tWGSCTtr2LNiQKIM6NWln3AoJnljCbi4pxOvRiazKDT0KWP7i
tLT7uiCO2MxrzbETCTh4p4Obvgb5uzFPYp7T6BB7y5GOwoixaBZUVD2hZsrs
eoaP8nSixeqJ2CLa/O4TIJTjLCpFMkBPFMoaOXSVZMZc8grU86QN/AjQXQ4I
JLom78FyHauoXT8H9IAfLllIM323msIG/dVoCuIt6DPT/S3ygNcGyD3++fDX
vwYgNU9b7iaeRPRa2Vo/18uABY+8cT4Rp+VE6PLhwwbLp4mGOpzDK4NRvUM5
qviJP13zV0BUGO02mezYTPGopJcjA8JiTTfIJ58Fm6Ka0NoAeq7BVSH0oQZU
sM+UQuWcx5EADS2gmCfBVXswWbk+sL6JYlf7EL2feS8VA37H3oX1BfaaPQjw
C2eNoTpfZflW+PxaibGaqJMfqdpv1sNhFyMHzA9zzCqMR1DnRz1P9op4I8dW
WtPa8M3pld/QrbaMdwzzb2XUn19VWPxos/bD7Co+Zh2KP/RfTYv9cvQaFn/s
Jx6phBUjjplLOWkEg4vJZQ5lzzJZv4Yw7KdJR9T7tx8TROE5uSD7RerVyB2j
qJNHjh+J7sPCOEq2YSr3UEpvAbHwhfK9ErH2kwrmW3vaug/7S6LQ7ywUzzc9
vVSIrbOi5NPygyYvl2GHIUy7qBzEKCHgCgCv+dYymFtI1YyM2xio6SakX6Pd
uxGxzeAakHEjMorZX75fHG7LcQnnT6uqHh9OM5NbuUdTySsZmUCUtOIWHrf6
XROXFusuZ/bFvOQhK+7doERlmDa51YU3LO8PmcD1uVst29AsKy7Ko32yFGNR
TGfFe/qNSI7q6Tn2rGSq8vGsUcLWvl76m8OVuf7epjXQIiErjQVwgO0HK79w
ssrNOtFyOMeT33a0zyEdBkWDeCMPP703+90Tl9q3RNELqhIctq8miRHCCOG8
K+XLWq0VnUMwOxZfI5KDgaNf5wgeeICCMZo90HeBho/qJicc/fENsl4tWt2/
nh+SY9v/etuFdXvm2RFMCqU4H3lWgML8iemSzeLYz3Ild+8amS/jB8qYuuhV
7F0cV+wSxEUWxncJdMdnPv6Qj1LnSgthmldJmoT/aWEVH3PPWBcmeux6yFSk
8BRMxVnXIOq9rGZsYtPs0ADMv6ojvZ03sw4ecO2e0lMN6BiXsPOjxJxSOItd
djI7p9fPUt/aAFRIkyugq6cYJkXofBhJfGoKGTRkGevBJVBx834ntf3T2Elt
q/d6k1Sy4EFwLVY9Papp9PunyOXFBhHvN+Cvx37kpef4++ar7NOpgg/kjUXv
OKnsGJUkxbw7qd1K9WtOiwCFdsdCA9R33EFSloO9L2GOB4KG3eiFWoKc6Bzo
DyuUitvTlBlQq4eeX6WthnVZdoUVw7bBEtDJxqgsNh/CEN9xZwsMS8irV1FR
0N9FVf8oFTIg4bCae0CZJE1A9dHd9OZVYHbu/Pmra7Ac8n2Oj30/52WulO7K
P+xkDf5G7fpCxGN9oH3Ar0VYFUAlKhrq967RPxedPZvf+OoAJ+RlQBt4cj6f
pdiEmoO/oAawHfPUfyB1FTnwsXZfavqDLTLpJURQRhjBLgVYYxqcprQ7n6wY
DGv0BQY4hq3ZffeYBNvtLqklasdaSW18FT9wIsfrtDVoIF6wm0KqTdlTB8yl
a1GjQxuF2Eq7tbqOAc3IYJzGNwNtq5yptSXdiJJFKBAYhIRmLNaDW7MWrEMU
Fgk/Gnt/FWZkbdwmmdWDRtFLRGPhJ8J18xJ24QJnME1gjtDejv+ptzNylx3e
xCAqCFKOMJK9htigfNsqlIZ74Yx1IEvgG3HZUo12sLINljlozFAqdxC5w3TY
YaQ28r6O6EsMHQby03+yhJlJbfdur9VqG1QOn0k5oPXeZIzbdF0OS6ZlDn2g
BBAxWyvcvDL8jEiTTn1u3urmOj9Rlal+wXOKXvxSAKZ+fdlbK7HG4RhcrUn2
4d8zrLEDqxk9jVA2B2dlruWvddw3k1HCAuqJ9btOil2OYeuaLEcXVNhL6S/4
kWSpOFpfhHdOFoBLFhOkzSzV/o0jm5e8SW+q9E08zN/ta3SXB6OKacYmOz0Y
kpenIPJkRxHJ2EF5M8a3Ok1UJTpiJHO0Xff2k7oSzhlyO0XSD6/7BG9HWdv4
3amVN0DfdoA/7boO+g95RcOfUGDNItTN/PKb2vMck4FyG9Tiquad6XYRS7dq
g3iaMgT9TIhavArOPCX3D18rkJh/imb5veq8OW6LVlf+hCLSy2fRxDBnBwI4
jm2EaneAJVp1uork9x8JaLdv1C2hGLKHRsWDq8CTff/OFlWZf81wapH/DQkB
pl9+kDwH4FyfQ5wqI8uUvJhkCAUuzP3TSLs1iiTGAZgEg9efmxZBLsWi/UPg
aZZRv4LhnxSOTWh8fVUkUXEVpHvzgwONZukVzFQSTtThZpCmY65LROWrOXP0
qniggvkIhdk/JE+p5HVG9SAWe2Aju6QMd32y0ukJLsSgEky8lyqBr83wBZVf
W8jBxlNbHAKSFcmQRCS3nBAnfjE/GYVOz6hkR2ERF44e5otv+2mvXIFsvg0F
rz+QsFg10L5ijvCcA+GWM0eEJP8YlEuJNz2Qtp2O6R0qGutE7GMrRedMD6Z9
7lqOPh0c8sVZCn39YXD1xD3zQm23ZK56sITd7KueEedyiu90K/SiRw+lr1BN
rG53e/HHJGKls+g6psUy+tAWsgzWUdj6rRkZobBS4jTBjOkbyFsNQVM5oa18
dKtZRprrl/90pUMThwG3OfDquwL1wvgW9IbYBR7lfTUkKosZFYKujLfGprcU
opeGPbstpIEGFE1wFc29qNrUsZb1cjwXhNZcLVL12/Y3g1WKTUhDZexQNb/w
plpwhaXHpwjRqkGY0g/OqnI9l/0jaQEMD0p9WXSsZMKolQNimkKWysj/gCSC
ggewE0YFiQy7tTy2uwWBAv+HRb1F0EYj9D8N2/rMW9JoT3Maiw1BXP6W5FXo
4mb2Vke0AIzdZ5ZVQ3t1CjGUuN58K3FzzlFfDak3/cORZv6IwensdneMb3xm
Bpw7IEzHkey1LRDz8GXraOlzguxzReeMS6h0YW9gDAWHUWlRzN7a8/Wj2vuG
GxUDRj4z0dPn4lDvT9qUPg+XunGS0LMqzpxLsVb9oxmhx7NAvCuMni/6kXRm
MYAWpyGqeVuBxR7KPwddDwgpuelzkcVqaH0gEy4lSNjpCAoe/EWW0nEbapWw
c9ThfHdNz6u8Z0Sfsp0YswM4FmEth4PvoO2wd7cz1FqrBzNHUtlMhD1iv29x
EKXeJPyLiyOgge9cRUZYt9xMUqjBymZY6GdBYlN4+kcKb3dim0lz0l8Y5ijl
cUi+jpA18UXipVJuhlS/T+h2PNGzJ3Z+jiY5SjkhYIWkEqmyBGQa0R+uHcvJ
BVV8bWKhPtmKDkGJJgUk0u/fjiqpCwnj4rG72zfWJ14wUz0yPpv+QWXGgRW5
zgtEJ6g+UVZifnrPLvEEr0UBeyqINb6Mm4ONZFduz2S/ZrKaJOnhAX4MaxUm
rBSCJNlyZ/gvqE+uS0elY28nTHMO3l5GcBmGCVK93CXJkr3KschuWN484kqJ
FZhKUz6FncTEP8NJSf77ExLxBvZ5ZwS4zflIN24hQ9ECHd8v4S9qJXxKY7MP
CbQdlIa2bx5QO04nPaVX73BYAbGAuvL4/+rslyo23afT/iIv4zi70S2kRn1s
uea3oYiA0/oOC6stY7BFV/AFSlXyc30OxVhEiNo+Xsr2j9Wc8WtfA7rysrB3
mJQJ+x5r9JjYhHBeRvAgjp0Ye+HgT9qMUB8bw8lPzzCxEeD0KZ1mJ/O1j9y7
5/sHCdqL0ha9+67LbKgUm6QpEsBAy2eLTi9UbXTEHKnUJ7IovH0fj06uaI/B
S/bcKyQ66KOltGO8kWU2l++Rll4p+yD0xQX7Jpbf07MhU6qG7Ub8FGHtPlhG
99Hf0ZDVzP6htpZGbLwSSHk1Ur+rXsJOweil7Y3Bo3vNNd03YJEF1+1F4l+E
jqGuqGoJtTWlG3XHU8LT2xxvl5V9zRLH0B5drvoDgrZtesaQ3N4NJXSlRbKJ
QFCg5q/1Mvm82yVMAIgdoiM6/vquLPjAMfJ5vGmx75GgGPyK5MKJGFSVnxYz
sBO3u29M1ZIlLYNUG2dWfhX8Ve+QcTHgrX5r9no0wTEZXZULQf9XWoAdJwNy
Be+sYSHsJEO/pURQ+ONbPuP23gZNY1ShqQWd5sZLEllE0iCST2cY7ZcJNas0
ydtliscH0QGG9tlhHYgp8pWm+D/AlGDWKpyw3HBr9GZir2lGiAcZTQTmarfY
RflKFfxGAaDl9ZPh+pSl8ivXBl3ifFnYSHe0PDHW6t2AG48AUYTd+cI7vcjW
JIHBi+65+eVPntPyjvT8antIBSxudMHDNrdoNernMCBa4avEaKwWx3Y9O30n
fYxOAn1wf5OmifCAZpCHHMOlF8TE2FzdLzRskuOehhWZDQQmKGXENkdm7pwI
Be0FBMEpyHpULXI4EXjCcz7Z7WgrOP9lFibZTxbw2b799vJVc3mtVe0AOiHq
eb57orQhEZBge7Q3xAhVdNECqZkCaGVKQ1PdNLR2VchbXkrsRqEQwQ7UeuwB
77ktcW3KbD82GIxh1gMNB6+QjQ0IZ/ec02KlWlUx6m6lL23UBIADOMH5cBMc
ruf/9XBie9hFN+vt969Fc89kkKdKXTTmOAbgcnhvnfXenJK78rjIgTm537B0
QdPiTlt8EiI5ppPaLcr79rdWZc0XO3acYtlmFtoXiq23qbYW5K2+dDHhgUf6
g0fJI0FuslEMBmVTFKa7T8WBMNo6DHF9w8Zgnjs3yCLCAyuF8cfushBNPRU9
T+Bf95QOps47NjmeVcIMhSlQffYxgHdzFbCk93WSi1RkDTaZmUg1chZ0aoYR
0ZynD4o4bhnsnrILYgJzxEto2xdzYT0vPphRd7dd6q3EytiuljKqpK3LwEGb
eAyVFT7Y6jFSKjkHnxKvPU3PEUTk7Auvb05NU+cilC6GJpgHImTsRceLWwWg
5FqYuG+iQdqLvku9n4EYqaz3uLw1TfAuMmNquJ2eLTCQ6wQMzPRdQd9s1T29
ZxdcOHpWyKsbQ1Sv48L+yCHXY3x2IW2G5LEWV8/rzO6G+et+mnKpT0NMQu+D
ZEzgiU6v0e427dJ3GuzVnR5mDfOkEE1nGZvJ/pbtaFEyG2pa3+fK5DDMdFl+
FtVYt3Ma1YfAwUhh4gioyuuKZqzdELoMgW2SyYdfUyRmaw5GqlPTRV7sTemE
MECyr6iPQ6g4sGQinap4GaYthcYSX+s8iC8ou1fkijkO5bU434sp67KU/M7S
jXHjgSwl5nm6ZW9B2bRuRTvgbhjhKGCLHatEwI0k/8fNvfvEkvcCWIu9kwgl
TYcQ9tJ9g4JuqcLRqIJtxpDq+wjsm1PX2eiC1VJaAtlBPV3NaPq5vmzAvGhQ
F0oajYQ4yLMEWvdHxtUT9X8tFpuc8+Le973ASyqvL1drJ0acXM6VjfwH3yG6
mw5RmJrN5Uw9OD/WBvfxeAy1VgzVy/8N8IcEUSA9Eei5k7bp6f4/bgqFkeHm
djvZtiY5N8lURuyGIFoxoV8iTBqN/lxABeUkARCBniOAgEmrfqyX/QNnpg2Y
cRddCctSBdyvhjnTQie1pl4F3T5hqGLOyO73wNlQ7MDYCTRHIhRqTmyPb6VC
dF06yuWgMyK41h7ka+zBzFFTIelseMLbV2H82nv23vrT2kt0AopQvfd53yNt
IIAQ8TfPNSdbu1k6j9OVpdR5JAUjZdAyU1VBF75qEZExoYnxQtrLkaLjD7Xu
Nqb588ox7U0JPOCqTs+J69jFcwvG0VVPdOo5qSi5UJpvJqwn+5jMuT6H8srr
fu6G0o3MnPjUQ2d/z7N9/sZk9WpjSDZndeKa99sLHUeO3n9lCWIlrFEOGZE6
kUTda2XJvgEBh9GkKFokJDIz+x9ZmxZGVsOUnyS2Ohlgg6x1PmfFjfEO8w6q
cCTV1Ji2JOnWVGiQg379Z/GD728HEuk4ivxsOywmwQPGFFKmmp9wtXh26v6F
tQLuE08x8vdXBpIRBeFwPgj4IhdjB04iO0JcX/I4qhIdIMxeKE7FiQQPAVCy
Wgbz4HbyHxay3rT1VprQ3ccBN/9LYRteG/4KO/WKG5Mbqc09qCPmJbwLysmC
vQ+NOz2ugSt1zgSQ+U9vmZv0hXwko6IqvQPKqBsEodhQZaCNqGEdCT5oGEIz
F23f3/PKYdohnE8kNm5QA14fnNf5GsuVu8EYClTpKj8l/0vdx5qxCaDHG414
eTCfHuHoY39TZ3HDDb3kIxbwJZGKBKBdfmaBPoir1YOvN7tpzSIbaS+i2fZ0
pce+5zhizFj9h25N3RnzAgKxejG/RHcEAwHPnlS6otqkFcQ2psfXqdfdWqFs
/3FBy9BkaBE1xOvbAzN8fv9fTmlgfD0OasFiXxlFK+E709sOQi9ZsWYSKzQf
uKFLK37tmoPGqRKg6hawwCSkI0C/NGCmUs18X4vUUxZSftqvnB3kilJ2lAkv
E7sWyzXx7BFiMAK3771mdTu42ZKdy0tQYKex9ymgKiBAiysyyh5PU5+HsHIR
CueXXHC8LdU6dCVqdFl7cAtW0loJn3S3+2CkD4fLRF4BWrgjpJF0rg6nwLqq
RTtc9tbTe+fCRYZCOEJq2MTeAY3/d0eZsQobL0SRlvZBELUBssekfpH5Vd3h
yd6AcIjdBsrWTr80hFHc/PxwguFKt3zb71FIMAPhbDp7nuw7/iTmF5t8wB6B
FPqen7tON7D8YydEcrqKiFjy0GPx1h6WBWGLY/wgL9vUnBYTwBWCzYMTRXjf
T4rH3hek0+f9UpHrdb0rwcOy8lDL9bxcsdfVR2iyMIDlAVg=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1K1PaVYXs1fZY+r3qGOph9VOpGGRhA1V/MiLJJgbG6sVwpctLwYcAGC2VAJa+GP2vQ5XF+TGKKUgvO1Iw4G1nRHqzMnxTpkbr2WHv/ct8GswrNYxiNueo6STFbxojJv+/C/zH9eBzrVfWlsoNdOMIuN4bDTNdACwLVhYuN9GyvWrvFa0AHNTk/ELfkRnqxgy/58477h8koDddJmcpr3uPkla0kdJGOZD6Dpcrtt+b5PScdIQ5o+80iyNJoKEZLykyEX4aE893TDqGVMQ5Ma9ck/5jrQX1zB2B2ZzhHAzHuOLtq3v+1V07nArzMyxPt0RZtpt5D4fP0lB9vv3tZCnU5DsnkP/8gd+688AIWP5qVehGjagpB+wwPrm9jtMyIDvCLvnRQkJZI94/0Kw7P9WLeh41qFBEdFYc7MQjA8Q26kwBctoCaFGvkJ2jrr616qp6Zu9isJINB7LmK257au8+kX4Wpd1OPAoEfoG0yAmvufhLhnAVhfkmuvTp8GDSfiBSNYNm2UPUhmUgzMuCGU7tgCkNHa4ISuq0E0ftJUcQE2ly6GGhSRyv/tqZevekxkpP5SkwdKyXmpYP3kisGuFEQNOBW/ocOnvjJk2vMFb8tEHqz+Tgvl9u/6EzqhXItkk0vxfUKlG1m8txLoEY0uQDu51FDbg5/nyJ+4d4en0rt4M5PZnhf4gao8oaNUP5nOg8sc9A3fRpNeJExGhzzpCKpZcI3QIviyKwXpSwEEVK0EY0YoFufsvUE4blNJujlBB+YgtlfZCtT5emlgEdITxp7Y"
`endif