// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nsNNC7v3H/xUXCT87eqptq876mVSxlwR4xqNK2sWGY+I3QnT3+jrz4+Dr5pz
RSYfpOMup1bdzr8xgJJ2IMIFHxfA2ZBioBl3/eRQgZTiTNP+iTyzHXnJsEHG
PAYVQ2WthnAJCITVOmchRIrJwOwUMXzOlPcNB1JFXnoAnmbQyChRHgKGM7Ft
TFXm15PGeUm1kEy21CPSjJ1bqtviBlHKUpLvFyWoGBCq8BbS3/5DRWDheU/9
l6VLP8rlleBlVduBc6K/lb2330lKBGzmRijgTkcx/JiwyTqvqMBJPSEBRl9Z
B8/zz/Yzq2m9ar5xR5n9hNu/mBpQo2STyv98nSHxww==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bHdX907LqfYQbrZ3tiw9d5n9ugr6++ufYqTU8iaDxLraiaUaohOklNz63kss
6RqkGflwDVmUOBnkeWFTShNaFg7FCLe1LH4/HUrvaigOxr4FabMHwRfmWVNL
U1lCxv817jLgJp3yy5wmsrivM7epoer0Abu+pdsQIWmLD6nrhsNCSvG59OoG
HpskKCgCtQoC26JnCiBfARnj9nEHpbKmFf6AQYzz3Ed2SxcRDqqwmRmW304z
qG0YzOlrXPGlKw1xZaWNdUDdEgPvCtf5AX79tmRQUsydgCvdqCXeSmCmXYrg
Ou7UaYsj10H1d0MaO66uaH91sYRZDgeDeUDTtipajw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jHDkKHvkNgtjKGfbI6pSPQRupKU9GDvDTrAPaghSzddhgsqNEVBzf5ATfeWs
5kJ3vRpXdtUocRFNczqVrqS9AjF9S35udy2cmvGkasNl5JtUFJ8YoYCLEA9y
NuVJELD8Wd5zPdVIOv1j2ydYtX5Ak10Hk3jMAFvNtnTbpnOXk7umSiCGFX3h
XOk/jHk5OlRp/JXb9AJr0s/N9bEtXhFMDYuyKc9xTQX7JppPbRuPw82DgyzC
+QNUd027neSRuSO40dFSbkR9hRGiNOCOq6xR5uAzNyysx3i0Cp2IJRC9eEXv
u+mIbwQCa1MDGQlGH3jsJdloXGEIN8U9Kh8qFTWV/g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Hi+YhKYQFe/jCEYqbqhBtcfx1LkZGHea7HDQe77FLU6pire2/kDMCZVHXr98
ejrEP5jADSDUWor2BlMdif8hN71ClZ/SbUTaL/xI7waExRBksYfCKZD3++xj
5H7SOLBSN5K/o8heTQqdzkXS6JGIxUUP31TX5w+i+70eByEn0nXt0AdSQLUi
eu73S6fU6iXwbm8cuqoPxBAmgXA4WGg0Zpyh0WxbANSNhz5K9c9/piQPtUXT
2qaqUxjFJ77wrPpvtY11R7tAanA2vrZ7Z3Y3TznUVpfxlNimdWo9lAbSbDoD
XbjJn4UqbrBctBNetw7/PpHr5VPeBXc8XjEnmgam7w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TmeAjJNjVwCCITY76c6H8epL+s+ArrNaAnVBD0/fQj5umm+kDVR6ua5laxKi
LSplzPKF4iYGgyyEJnu48h9MnHL0huPXIJ7Lxz8XpiNc4Vj1BuKCt5JRKYT0
x1Hv36hznWMtswzShyaV9c+Cj8RDYC3cAsHJB10d6Pv184cZGdo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
G3UgchAC1x3PKq6OivfRYoIQmKzZNYD1iweMCHUeK3ORKG6x4wizCWSm1OAE
e1tUzORcL8pWg6zk5be4FG5mJGKxR0CkLGKHXsv+nC4lydE4nIOu4pziXZMf
6y6G6jdLWJbYhcEd9wNbbV/ANdD/+iD+0ji6PCLxMQRUZXpW16JOu9JEByBl
hFtju5ieZKFbqvI/iCoGhmpev8OrXx3E23VlMk42KjZU5vVhX30U0EGRYU3k
pEIA5WtgvQnr10CR1acjenXnyqaw17x+RaT08+18qAo4x7aDTCTXPCutg19m
XZkZuHDAsi9cZo4jAjo/ZCSBspLaEkhchRBgsCyUDRhI2L8T1NDgGCsSyrrP
4v/W0J6cJQJEyYM/nK1IbmRT5LcLBvItJ7gPAtpdakFWeF59JxskaJaCY8z4
bkimcnV+Ix2VWocONMY8GbaFuQTep7pH1heLtuaWxI0IPM15TUp9RnFgSWXe
UYaMyOhv5LyclgHMu/5A+ELJPDJNDWwr


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DPZfIMWyPwFMwVwcEE5PYwLNWjE3uFNV2q/5XXcoSayq30ujhA0wFxqgNrUI
5w3jX55kd5tk9h21f5De6Sd2u0EY90pwyvWfWZTCouX0euOE96F8fIx8Z+Of
a4on6JW9kqLQlVm6KxXbyOuAEEzeuFEW6Z/vY9PGa1BdySCGo58=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dP05LQqjy4KnxduCx9ggDD3rtySeJttbr9eJdw1LeHC2+CjZrVwwWy97ktcb
gpKL8Rd1VjREq1WRZU79ottqZCoZwZs5NS/Rmef1vkNPuouHhERfrwsic0fv
LoqHndt76Rx1BmuxHawdM4frYWxwqIsTo5zChTOiT64s/TMNQr8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9024)
`pragma protect data_block
rq1B3Z+AH8B6+g1NSA+yXngNnWjQBee/d21B8BCc63VvcYHOS4XPYCaClmRj
JLXL42WrVeSC7TNtJCEqNizOxE844uXCO5UnZgIUtwUr4BORnCTU8rbcrLgi
CBCRB098lsbT/XG/0WMLi8G4WZJrRDg8yqxkgrWzY47NOyicFig/b/2el4Bp
45Nj37yXyOLDIa5k5PcfRtRfFC05d4IS7UFTvqwRNWDWZBMD+tdp+bdxaPOy
SyOicqnrpmQ/CybLO2eokKwDTO9tf4ZqegVAZDG8r4ZpHyp37UVXE4sv5Fvq
Mlwj9BhBJzectrK0345poxigM2cdHW+Aqt3n0YCQHvV88J9JP86B5IeUrAMz
KBfVoTy9o6/QFoa4W6ZzDKJBfknTGA0oVdnbwYB/7n7NMwX+aTH6SydGx+ty
j7QH5aEBWTcIpxiSNGlnRkQa8KfyyzmOtyj6u+8/SU3gRJlVWIaxrwmA3v65
HOeetI6fnNyv7a4oq2/cxEkcuo++HsnJNUeJmBN9bfalHiO6OcVKJ81pySm6
rGRoSJb1xtcHQghEjV8DLQRzmEheygwa4KxdTdZ3erptRk27QtVFCDHy2MaG
hDX735+YgRgzqWom1u+5RMwMu9PkQi3ksw4DJii2zHpq5bf2bogyLMJEJXeu
4t0TnaGcXRAT05yvxT7La6tPXFn/LmfW8xkX9m8UvaeBK5Fh3j1itfo26RVM
1Fu+GORb2+oKVKn0noQuGaE28n70ZELvNX+kjK0AR264w60AeDhijdpBf42u
ulyxczMDUJw9JZgltqmZ9opLaSIQGo8kzMcuOd+eczWnVMh8DYbxe1qUpFwt
dhbB7We7GxTaSor6JH1HKM4UgFw5ky36sHknb5ut1OxW1IdMDEwrsGcPOn1O
dG/3U+gICNjARBvdcXd0k+my4N6OWjVhNu29T/FCM6EqOhSEUdSolUR62JV2
DUUMaQgvRuLQDcTgsJraBLQZoAHwAqA1SayjxYE3qsxeHF73RU0M56E/m/4V
Qal7AU5pO+pY71rParEGOC7HHlJLYZkA/XOWWJOaAsjBxfY6q3Nhrn8EEkdK
8K3OQv2SSmXjrELe3WT0G6PE51O34sqOjTRggp+ePIuevkOkFxZnkkvysfct
I51NxBpo0QJxpg3E0yHsO1twKTY1tBMPW+qFBPMgBaaWtYklma7VciXQ2ky7
RJLX04oQyFO8wq2kc+X5RLHHMtrRIlemLdOuQmoT0UsJttI6EeQYXEk2yRSq
YcGL1sZhhrg6Zx7ghB+fkmzXjU9fP001Vt6tjmKnvIwjHXRRfO5JjEWIl8nS
l0Sf7aNe/NSJ+PZfUtffe7SYyIAuzWeeHa6y1s3jESFBL96EFu+NgZkpdd3M
kxcHjDxyxoDf9o9ucZGhpS8udeFvTC8NcbgXisdFufKLU6SqOe9WMVkktkOg
eEkFaf9UPq6J5e4QFJp0vSlgBxAfR2DJB0hx6QTYfor22AgPqf9g+X+7Qxhr
HKOO6meELtE4AuLRYPuKhq7J86mwsMZxhWvn/U9dXzLi4DZHORf1dFSRrKI4
Qq/VD+Ql0+qHMwbNArNvPaVs+Qbrn2rUvpSUAay7BTAX2pt6n6zHBUmbcq8/
suH8kVK0Ut5BRF2XSkTF0rVx/gycVuGL8BEas7+j+fWTCZKmm8m8zHZyFA8b
9q9iTckyPKAHtBk8jLu9gyV7VqTpHfCDiM/3F9HNCwRSARdeAav/4dyQ1V3a
udBUOjQdoFIOssJj63OTPk2qs4cUZHoKwI4LJQ/6ZywnltyMS645lxsbfTN4
rUjOdLqMjM4PLD5Ui2d81b5TiZCcUzIcWiRF8Z2OdXihRhLavqg+PquNfqCK
wTj7t7C9vNtVg6Ul6TJlEVXI8xFUSGvcNsUpw8W7oZMxSQCcDRrSux/JZtqY
VohOivmH1te63vdi5V5PHTTETkGuBc7CPgDkELZVi2BRmtkb2Fp+yrBzznpK
Kj0/fDY7aA3c+bw5Dv2cs3bRKtzu7r04hU46nXwE/UUMPW3PYdUBsxuTnU/0
xBjslDOa6x2HjMZkOMJJ1MD/c6o/9+xSkzsxwoeR2eSLovMZcMeIw1cvFZf3
0J5WMW+/icoJcIdiDeGqhCVe05VT7dQQz0P6u006Ga7/qOUSn/rSSkr52sD/
xKJW0KO4UsJYpDt7ine3M2LdntqPYXF095ebumI8sXBJ+SQrVrK8KarRuaHY
E4fH4S647zRA5+DqtAqIPWOf4MAtq09xZ7rk/C2np2LGNd4Mvh5PXHS4EouQ
y+9R8gHqhjJHiL8wbR8Q72AJCh+oEI06IQ8DwflX0cn0UgYOnjfD3i6CiKo2
ZYWI6jXOcXaUsJ/MyWCsxmHuQua4RUF5bc5hXnt7n9qFhrX9rdyB3juw/mSv
WzqecHSHL/m6jE85yBrHcI/SJdxQz6vIE8YBzu8Sc/EEKQ7hoS4MCf6xaMYC
aQ7g+1IsJDXZm1gXrHnkQcWy+z3zq7n9/ZIcqsESbGL10D62Uih4DXiSUJ2P
Iri244FSOeYtFMORv7Z9yTTrYAIqgIGWGAivehOJl1Y9XcO53X4TNFNMoC8K
jtT1xnvWI/3dpER7o3HnDA2kiEEaHz+F3y5wbTchGdH6Y/zpcdhpp6vReeex
HMavBy/Ya+Q2oDldSAn0hOq1rysgWzqnIZ+3LXJuPjj+Ibd0h8SbjdemGBdN
x0Dqzs3kuet5oJhv7ZzvK/xkBdMbCGBhbsXW39xrhLhG8fKtxW4WwyRZVelS
A7MtjbDPlNaukwOljJ524+jH1TDPshpJexugVD6o7cs6ZQiIhdbd0pdBM/Cv
xlZhXqQsgdgzLEp4uToXLwqkofE8PbXMDh3+1X/wOedI9oEG4A6LcnoPjCi1
0i6NnPI9KzbkAfy4u3jld6yq33xYfxaP5b4q2oQ81vqc6A3LzCcuR0U/3GQ1
zc4oqIqIKjc5kFKil6h+HSqSrlbiVq7AgPcrQP8sQPPjkh2iZGIDX1JLll2v
AnQzP5UaqpIVjkUDqpC0whh2mV/tq5w2P4hdBOwGWDDL5EQnYw+z2Z5hVzr9
IWRmz/SPHJtoaoJa+i1IUMDYuip1WSac0VqB8yCMOwr9PoMvkSQLqqeAslBC
3j1D3OTA1M/iKlUvyrvwQONv4sQHFE58LYXcUb+9/6Gu7k7gSpv8sy8n5BhJ
2LEdMLd1bfhya1+Pq2khdGhqyUOD8sHbF2hbQwcLgqAcHlIWeixaFUq0a1UT
OtHQJxv0oe7XxVgD1tmuZ8UN8zuz5kgZwwwtsKd0RoDQKMkI/UK7dqyLNub6
w2qK4t0jpfQxTNMgBFN6U7IGUAC1tmoSWs0vyIgZgUv23bjdqqvsUsF7+WiC
DKEU0NjRjKIKfp1BaarPkrZx5FAIsCD/aTDDq+JapGi5/8ZHX2pKhOoiN6WA
hMA+RhSynTrSTvfY+Dm3MsDbZsd/iQ/MnBR4Aq//B4Jpx/V7NAH5I6hLNfK7
WlhYCDavb9o5SVAEDpqFsRDEmHHnVoiC9x+CAt9eFVGKxj+oaG+tNIG+jI/6
t2kK6VTxISaslpuqoJCM9hZuLiZJbOjdRGHpyJ50+pvqcYYcGIktDlh1q3Ll
PfBsIYvRh3Nyn5wPtKHkZDc4zlaRlVMHmOSb5CAVlhIVABkknhjQNtjXRIRm
RITTArTO66cUku0u7n1wInc4KnThDESP6K1a0le0kPbFoGdqr2qsTqSwoVnl
P0c/0rWCU4hF+9raAwLpyPU42f47/Z0GIBS1oYBtEyHo8d0ssOxconoP3xtR
/jwsfPRxj6J6SvnrWznU56JreUuw+SHKd5peVVHWJDaU3wzLBlpTbu67iJpS
3RVmnO0349BpMKWpGBW9Ntv2tGZgo3qDIKZVQHkFb+agO4gEp74Z0MXifapK
CgEQF4Q7QOfBLghM098JQRAuN7dbi4lXhV/W+6G1VnhsnqgQ3ZQJy0zRLESK
Z3miRP1vPmIZUrXU70u37jB+EnidkrIIH/Xm1+Yek1Jw5AgSiHLnsBeMnlEa
ToEBO4xMthshJyQnobPRtqdg+3jsLHtY9tWLsZsHg+Zb+1SISKeC1bXB3+Lm
STqmQlnP9+StKkrjo1KotiiqvnEwygxvtYO+oqk2uLNpranA6CfQf+4QlCNA
YbrwQ9VxeffS9HGog2pi34YX03v+/YsOtfnVzxXboHI76if8JMYQLp1dUAj5
25SsYa9Z1tRPalpvngcQlFRlFO0ZOznH0JC5ZZ4u/EyppsQJcy4DW8CRoSHu
1GdqVbFMXwjUKOmX5RCHFspW5VCX3uKZ65aGTXu2nMLJdMAv1ENOWBjChD/9
/hLqkoblGJ6kXO9tzZiIhzaF6KqXHWA/gSX51aamsL24hokAnt4lkyORYKan
d9oBuVUP2iosccUGpMl31iONkmYSw8TYspCotedi9iDRY0+jqLe0NI/GxAKM
nZkASf24oVfa1JWri9vOivI5Fv/5nIMPARtiSQswRVv6JImonpwRoOXeZhdf
MwjIsk3tCHAu2+kB4JG4aIudW/hWZfsgJ1MMjwTAkmg5y4Nyf7T6tY3rt8F8
LUzsFdQbiktIRl6BIyR5mFoIR394pPx2aMMYuyEJERmcjhpTDV7lNJGSGFo8
blyDeLfuyTs9Hz/1u8JGlnjJ6o+yOL2lfy/0CKzVBUdy4TWBnQ+ph1sb/XYQ
9y1a/+Es1zkajloZr5N439neNBaYuAKUCzdZ1z6TYcxcFiEjW2LrgjN4BnV/
NLMK+qOzmI8DrGeqKo8A1EIPQf7pSrLb+dX1bs8Pt/pIHSBcmr50nBvaOzy0
0u6OWuhx51D1l4WrYhOS/6A6GEI5CNcd73I6tWhlKkMJoat+pEhsWkPT15Go
ca2PY/dm7f1yV51o2IlJCOgZktahWyKQ+Bwb7yV9VW7qKBrYuGhDKJngljY3
zqoMoDWyFk4gZUvOmn+KfX4fP4Vi/1moPe/EoRnnWUAL8FhIhXEj67M58tDW
KYPqDz96jsm/RD7Ijy9/UVzNS/5ishaU4KYI5L465dKirXDTOMYu8bDAy4Vd
3octEbhsdS9dH8h/boHnz4oIuk4jbK5R59iJNpkEq6ZLOT0iBgeBvxeTsfqc
2/x0czCqS4hUkffTlnhe7f3DmYrocjmJ69eGpWiUJWHpoQKgoNvRjbOw8/kI
AEDtuf5YpY+TfBsHJiKQVlkoCdDRpL4Dgnbawa7kIbjr8SelrdAwIai/Z6Va
Kpp5fIwA5l83/RcefWlsrevyfkA/bgS40k2teGYyO3JIUjDNKOEAzJn3VkGb
n4AW+67ompB/o7DxVoO3/pUAvreZPQ6ADEXXFm15g86H/lyo7rNJPEJjjCmp
NS8IsyDHRNiInV/I8YB+T9TIBKDmiYD4aIrhmLwY8PBAkMS/URJCX1dtNRu9
6D4XhqSTIVqjeJas3G0SDaslNSCyilpHDwTNAODr03+Eii5R5VrrG3c7MOpc
2aRHDoRuTF1nUpNAdELGCqd8n2rfafdqktI/Nm7apmPXCso9yIPaDSKWNNw3
WnuthOk5gYcAQhs119rGjvNlmE+RpXj5QKlN9NTteD8YU38mgx9Kr1wKQPmC
tJr9Qz9HUdnpVx12w0sX2DqIq2rdKmNj3doV+QJJfOtqgl6Y0KgNVPbRc0HH
9ppdfvx13ZPZjQ0Q8ekvARlCbAsGq/WN4a+rLbeSjmPXjOvrPT8q9a4hEBaz
sZim+ZvuYL0V9UFoP0YVM0pEu8I2fEft2XpI/sgmqksYRT5t66XqxEzX3e+U
zxW6bobjKDwMHLI77HQdnB6eOW4YjPUInTNgKKJISKGRt60rIYAb/lvdk69R
B9NecbqfBfyb9OYdRNHD92Xa6xxCyjck/A3y6Gx00yGN3p/jBbsIvheXrI9O
5wpOvBfX9vAgwJGx/mGpqbNom2OU2SuBZuC39J/ox/YL1KOK8NL6OkPfoBo+
scW/slo6Bb4DdOir4K7GQUiJ9HcOGk6IRHoFpnNVKpb1R3AtfXX/XY0U0DHw
96HvLjIZc3vr4mhdzT4+63Py6TUH4a+62DYKj9jMGhvs0wmyXQd57ois0/wt
J+kU44jCbnhL4EM7VWEwYgx/78f/pK0C/Geh3sUU6cv6s9syacr8KzpWTRBz
DKFH21lqfd42rli1ZXNJuvXqVoOb1ByKtNXXSSwOT9YMvuxeOU5E0RMe4Lu+
yWi9IPpQwJDeJvv9rN2nm/pZxv4rmw+XIDRxcsDfII2d7n1P5EkiT7TKyVCy
Sn5V9nfzawps7umzf3rKZ+bSdw5q53+PxPbyQcc0mjFt4gT5kLHaPEik+u7X
QVuMzWftXRWD1TMaUt6BBbGQRHBWhr65UNioSNxDKgNwV5N/RGv86f8TOjXl
01YeCDwryD09POZwwo1Wq1HIUk2FYHvBWJqK8tEbYTHNdXS15wDdDtYS3fhq
cfL4y/qoFBOtj2ZCDmElZN4j/0jUMQD0PDEMCAtX2TwtJX5JR9QSHQtj2faM
O5MlmMH238fRvMt9eTCZ5qUdfzPY70Z96Cpkx4/IxkWpvQg8d0f+k+LatB4t
NEoXUPRPU3KsBC0fsgPKkZwKjGJFItWiL5h2RVXXFu6+KUroKVw/0pMZ+3aA
IGqZGaTl3/0dZnmQJ7u0MoI9m250VQ7QEaQFPygiPa4KooXE9XiLsjDscdgj
j3PxWps8vF+gGesWbLEPIb9QNLHrJ5curdpl+XiHhxfErzzi/2qeBN1aRs3b
vKd1QHEwAtgmGF2Fln49iEuCBXTZCsb9XpoZYR3gKmb6TIiRpWZF0lh0c0sL
nUu1V0jeGeAisFmRf3QFc6K7N2Ahz5fIP4KwyisttdwVmUX2R02GMGXReUsk
oSAPInR5E6ed9+0D2BvYx/48gMgUZHqBNNR5G4uJIkU1DUmY2bnltliPzEd3
1P70dcRO5nr+7eckJspciE1XzDMH3Ug/ul1tQpo048q0nc0j48U6zhiMu5KV
TqnaWSWj5KPsynN9cu3ALJdfqvn0mffG3E70ROiQGs1TnJqEeHl6rFrtqKDw
nLDPq9Atb2ezWzzIduSZ/Bb//Zc620weUfB07enXH/5ItydIAc7ATVk4AvTq
OLqQSz4BWwAKTVgTdJMW/U0ZElTEa1Odbkz8O7AYHY8pHRcIuKe3ZFOvc2VZ
CdRD/U3VdgoB/cCezeCLrknVKe+50RaIHU6Bn3DX/J6LyE/Zo4ue+RzyX7jB
c2klSBXeu00rbWQbs1cbK/lHQz/o0xHkH42a5RV5NXwG2Ef3ayrBoQmgrboV
LDydC60FNJJnyj/uO8s4V7QZCTIXW7exZbRCFr20/R7v31sbaOvqudaBRStK
U4agHtnKcgVr3ADzC7IUiHCZFKxNs6S6SOCgAeOovv0zQcZJxL45qf6z2gl0
cUIo6HN1nz+2XZfjT5RzLt5WdoDLXel1Yb0zL9uWeyxgrYWmJ7f9bme8WM3L
E/4KTOb5xhpNyCmLm53TRqm1IOvdLLG0DI49xJL/ShTiASRYrFNCd/sjGtnW
4c4+6+Gw5Vy9PF0GuNl2EqDnjG3If6viUgUgz2n2F+mu36NA+odeiuZ1AKLC
99kS7ntl9qiVYJg/7u+ZxWpBbKO7DY0tOMqDYVwP5npBnTDFMmg7z0OkJq5r
xO9ZbZw2K47u98Xbzqt9tcaZxUpyLCjhygzffNG9oDgTRpxaUCnQyPOKvU2a
pgpU7oi3LolW/tvdA5k+3l73baKvkez+dni+2BabovQnGDAzESTd04qjaWKK
Gq5cumKd/N5G8reaAhm4dQ2RfEOIrGW9Fe/PxxQ6aLY7FVuXA4dtXr3gTzx0
NvqMRWn0CSpeoYk9J+jbhPbMWAtEu11lNYCnFJqzDohHFmRzqLdQjZZ6Ces4
ZsKOrjN8gnnw4f+n1MHmxds9OYZ9TDF89PNbiVOX4756Ua93DgzG9zZqUfv2
dtA/NNo26IL3M2mJpyNK6Cjrf1jp8f0Lh4QYA8g8dzXIu7Vr3BPqKxpUM0ee
ew6BuExorDy6I8q9UuAsMGTrxLeDczyJohMBQKJIi5wihVLfRlFbACe1/0RR
W+w6kxsPZTiaN1onQVTnU5lI4k0c5JJvq/Yz91CIWRRJ8SpIymksTJQG8QEh
iddLx6Hc9TeJbnLt4u+3Fyl0G/rAVFhE5RTnephU1q6WxI01vXmUQEq+sGtb
tuw5MhxjIELNIPegwMI+Zwj3i/2Y6cCgVPwR3mdvcXqOZYzg5eWguYgRqbBA
Iz65sVzxsM/YDbQhe1N/QQb31JmuwUEb70IbQH/O7f3SxvO95XrhU+kCCGgG
YPdE9k2NHgBmymhQJt8DPeJ9g55NkVXWuTuRc0Eua+JVmmTSjB6Yx3XJd73R
iVHv9fjIOEYfTSOELcC4ptwEFkNwXOBxS/1ucIa2zkEtLILknpyG0XoVIAL3
2mhqIMJZDAXa4Yj7YFCnhbBsy5RuseOEft46oenVRIbr9RYqHOE9YiG7sek1
2sM97Ryf49jNZfcikKXM8JQZzuX8w06DSCf0SWwwauxkh0j5tGoM2v0pct3e
eNdgW8I7AlffipfYNyXtS88grOMWXoHyf9KYuYzwqMPdjfhTKQi8QEkb19Xq
ZPWXpPtCdb76+0fnB3KtzbCXyfDMGJQLksg6cD0dH7FC5ubFB2OQenQbiJAY
PkE5cBvitYXy8/q0vxvPcLg299hnHw+IA6HOy9YvLU1da1YA1t03QOo8BYuo
6L6WtErUsUfTfTejTzLMp3k3U4kU61vzGRVhQfJj+LnVQGV/wxdtrY6agxEk
xrK2TA2ZBNu+WjyYa6+nQXxYWXsXPSvubrgO7KADdggTyeGUQ9HDcFaNh3+M
XQOYyBq0BCOEm8bQW/Iqz+lqBpk1sNiRQW5JqlyY2w6kMS8iNuVWX4sjKjDD
O4N+Wx6a05JzzmGhCoNFB9nKN+d1lBjicma3EJo/9R1eH7PnLIbPuk8ENXhy
MX3yXND++35Unt+XaIPjXXBhOkEex+7xdXSj8WPwdSHjYjZ6SlVPb7sszJBo
krbjmxB2hhcXjaJgx4uzK2wdlHFAZH00n1YRdsp9e/DGkULA+4eMrnkd9U3s
Bybt0G7MltaZPBVs5XPehQT+nzSg3Fre1myIpWzR4FhvqUMdxQCOF/E20nf0
+IawiMEvP7T4nChSKEmXaL+c+gWvkP6LJisAAp3+UfGNWxkJCzNxeV0mDuIc
dE88L1lsM6Ogo6BEzqv3RPpAq7zEbbPVQ3Oh/51y5BVYv7qRie6fEWFHEl1P
eb9+YVJSVJFkC4B2tOyu8cqLidJPvVdqaTarcH8ryOfWJ2G2rKpA8rhQD4KO
oIcjm6YNMSGqYNmMNGjXOJ36cE2kFvDqcQDbUu6AvwwQsa2VtfUYFCaCOqHX
z+hOx84/rgO44Od7uFy+bo6dWYCbEjMAYTx4N3emAtkp3fSIP1NZWFU3nsWz
mTjcLNQnh1VLVBMmADz41ARH8xJWvE1zHfz+pTbmmpGz3flGctkfXy6H8uph
Z1gNgQXUxf2x+c5PBb8IMc5QF3CQj49d9tUbCDyTTmH9bUnX/MvaWf/LNc8y
mMfOBp2T6XoK07p0LjQf6GAB25sJ2q6ISPKfcFGvtdFOgt+Wka9IM68Kpa4m
okljm+BeaQTV5hJEdzCuPyMKQ94+9TLx29VyZsOQaM7PqyvAOYjqA6x6rgTB
uXllhTZscGmtzeaRjkkzz2Ry1I7Vhyr0T1gAiZCkvHSibZgFrGVDRxuKpjf6
7MtjvIcvucrh9idDS48vfpRUCGvmt27/FPrgX0dGBjAA6N99Xjm1siiAdXBr
OXpKzorgxPvNUA0uV2ztvXiPnYVFwKU6YWT4F2LSDyAH6T05/1/+TUl3G/Oo
g4UPXzjAMlhJMCkSfQHT5d3XNUuzVRaLrh+YaKeMhjUlw+KeW3tg0JfprK+w
QRcn0/v6UD/PJuBgAo8OssmqJOmbsYF6VDYKgnq655nfUm8nfPNP8NXOau9K
BNPUNYnoUBu9iQ8hCXjP05S2dTcQ0BEsnzMhVejs4R/kOdK3OTdxY6sUKZ0g
4YZ8ab00cyEYxGioPsLw44jBx3U9kkna+4UxqCrfUwn0tYiIiZ8ETTgqd0jk
wQfo+gSg8PrOMOnm1yreWjejbGlOMF5YLyJF+DjyHXs8kLdIDbtd2pzS1Z2J
9+SmN0Coy23f+U0usoZ2e4yawlI+aR6VrOmIz2ZKl2XHk3BOGPc3o/qA2aa1
8B2lytu60+6/38X/oXQZn/jWM8kvjZjQXDa/D/wNAarvPwvxv4JVHY0z9oAA
5mvqiO3wHq1vXGY5t8qaN5jL8tt3t7RE16A6zcQVYHELaVxyGspR+ICHbeRL
bsDv6X3fQFQofG137A5wH5cMd+UCzznElFQWuB1c45weB3HzQW2uMXHv3zhV
0+UvDZtgmuddzDTj0Yx50s/mSSUfyLule2CLg8RCX6gJJjXsAZOod9/2HKa6
JbgNqEuFNMCOgSoBDrHNnPUMkQxq99Eal4cfCz+GHpxc4Hd3NA1YG6xj7Tdt
WjcnF9TsZqg/6+gTQe83y0mKn9SjKWgKkZunmr4EHndh+5dlXvJFi9PkNoCp
ZZ8zATDIiJ6xLxSfk1z41/y5PT3cPMhUG2WGmxzvYRI/1AdoCC4hNR3ejHG5
TFgcg3Gt0562NakbnhJA9x4+7HDVfRHqA3uTrZqWVySX9aCM7kpelarb3bCX
UZ9zhw+8zsO4MRgJ2Du0cRUfpEDTyog/X8DshPQcyUmqhdDdSDGoEwLPbGey
2kTo5HJIrwQ3IB5Ujr0Yip7lqNFpEMTBdKLj7XIOJBpiUURIjO89V5WRe46r
7WKdmB/k+NTkYH+JiR8XgGn8Ubtx2k6OJEhwcde8zTtynQFrhynyXoomGw6m
tLGfwGJa6KNVstJr7KSGelhTDdDZdd66fgoMIP9/dsd8nbt230bGAfcFjGm3
O/s9e7lfIcIYEY3zwwsE/D6csMZz3ogty74kiGo1T9gRWwc05Vmuo541q3NS
q9BaP4T03TrSsl1lq45rSClrVU1BY6Ip9TOHpwyng0QkmMtEFQLM57Bd2zwC
NuK34XDS3VyoG4VnHj57TUPEII/Oh3V4q6vDyjVdX7wBBB54ZsD4GEht+btC
YTpfcOOuxnjmbDyQV/HDhn/TKYe9L/KUXTr+MIqjLiB3AigvHGdz+2eEILED
D25wZyl7FA8+3+ySKK6Q6xWdDQAqQToMyOmfKtewuZv/fRMUf2aVoXy0ns4R
lYFirdw5cxkTXzVCMpVVrmRqqUo6c93O9Loa2L+KlZzILjZKKfZoxwwhBCNA
Lead6f39wFj3Zboie+cPLXseMg044+ehJ8jlWokdQ/+IVtP7vTbpCvL55IWa
yA7IjC524v91P+2LQjOPDkWwEmh4/5a64ulkIJiABDfTr+1cxIQhsnwDGgG2
NaBklcnuiQexDeDqR9tQc/AZMndhUxuJCBrs+Scjwlez38/SMv06B9/FzcXH
vgWbhB5sUCFHAMWLodmbi1/U0+yKVjVI3UkdTy75lC04rOr01WzJ70bhh8Ji
sCQ+5xaMZVWH83GbUtH+PdJK8XJsQZFRynQMTFMAZKzvAni1P3ZW6jo6i54E
Mrljlfw404m230upshyHPjpd0g5KpkVEeUzNbZ1WI4Bv4eZhih+Gqn+EQUus
BY/ygSpl8q6lK9MQGpqLnD0MreIqLPaUIbyrxfmDJpXKF7Gur9TkAjcaFkNq
NAtPAnZC6MH95rgsQ0QlyXWHav0r/OlX1KWxH7o8iIIaWMBVMe2+cquPQRmJ
8hTabC8AUGl8o8W/dVhNjRuqk9XSwKly3aLf3V4y5Iv6LXTTLZei1uN7p9LO
JJ90+ggGJmPdMCosv4cMGFnylK1HTX4paL2OZ8ThxApjbQKgmNxtUDN4nCom
YUqvngYdFgs/dAu3V+xU9yMaLh9qxzsnW2q/6Pp2PNdFltUg2IL7tNU0pJ4k
Pt9ye5O2j8mwPHjuqzqfAfiNIjnrBSFpXIRndSNjPL+4BD7vYC5U6SVqAcwM
anFlTyfnIoFFJOXSUxsX0Jbk9bLGx8Zm

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Kttctzi5aPKQ6vg9w+1g45z6Da0UaxXtt50QPmQzmLiVao+5Qg/yS2eSRK3c1uFoxS+G6ngDcAKHm0LGGibx4soakCOjaaRTqJmqblCXBo4qigRRJU5sOpNJWGKfxZC9LZLfFjqN04HCQ8ah5FN3P2yNU1iObRgi2dEkx758LbIsGmsSUmn36d6MTHQGWCnH/AC+2pgOY84Iul0q5eg7DNO6RSxNOih+2JmnF8szbMNn1n45Z4Lkkc721VRwIqdJ5W4gnHFZC4yl4NK++e8R1X85i0N5Ko/M785mHhQ6gN3sci2WLYxVq7aBFotNOPU/LDG4bhY3BmOvDsHBuK8pgilHfJDWd4VSjMaDJZL+fHNj5e34+SP9LtebpE4c91K1B5EZvMLyC9esmnsb6UxHLpMIhjDgI1op7+usB3EllJTaUhJvppq8aixRRSMRS/JwGPTNrffhCyX2ODH2XIjJZZwLajOuWEVegdkbKGOEL56XkKA+n4f35gqVED9/hQN960EGbUH6iiMiZ6Wud4kPF4FSwC1gvRJEGFAkSeTaM8DMwbfT424QAqSfV5mU78MYU6jtZFscWQ10bsbQlDlq6n+A6apVBVvWOd1pmGCTTmb+yDzUZoP0jWEeQKYwVrGSlu7QqpqkNCEVwPi8P41t1pvsPi/ea+MqLiBEMXwJM8s7i7OAHYIRdFgn6sF9VshpMGi2iZUst2e9dlxfSfu5MnU08YpzhyFBXC66yoSoscUf7zPoGUUc4ToeW019VTeMWq+jr6BwhxMhuTkpXZGdVTsY2dg38Xg+con1qjKjom5YKmIRDki5qyf7PjlxUsGoHhykTKBxu2unFz/l/MldePbxkM7DOLWbaH1EbAgKWj6II2/ur18E0NBDVEYy/QA9ys3mfFYCeCT3JHNSJOUI6kXhs8BisWwASRrfhsEQ8cgMXpjWO2Cvrz+5oKuHmIMD+ehdfSjM/Yf+G2RvXvC/YexHSKFnzXd3eRWQzi9LgOYgNltfVKlzZ+CrcH3PgF4V"
`endif