// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fy04N3ep+ddFyd+rHPl7lV9roxmbLxyZh2+gtx0T2z605sY7C8MndwZus25g
BJBhLjPkgQhwXIQjHTge50V6ZNKBzJnPtYtdIlqEiKXY7e1Y15pD0HKZs7kv
HJ9XhlB2E+j5s1IadtLpwY5mcPFrC+uznQ3UNua/9+jFpQFINOonD2/lpKRm
atIkZiofVIdRCWtkblD6qPTCeh+C4cswxQiqhGo5Cd3TJwok7bxDM83Zfy3J
J3x5cfiVwl23F538+ImHBKZcQNXAOe0pf/GTFC3MK0wlL/uXutaJxELUHZBD
x5XVHb53n4zRVtRUmXJ5TBcbxYTJa5A2G+sqU1c0ww==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Pzb5t6zcioweguR1E5M/td2q158cKdyNk/G4tzkDMSFZmyaaDux9MGoCFhUl
86kQIuNoszldfAqzoeWvGrE9GlJO9FImb+7aHFr4td/06fNQ2nSE4fld217R
2Y9pqWH+qnxzvuW6gHiOc+B3Z6riBTcQGI7nZDvx9i461N14MJ2b8sTe8wEb
cbRIFS4rxN+mQ/Ys+dn8DGg9cp8gxQoA8z+mhpJM38BmKQFRKcuFx5U4kPP5
hTnjwIRPns06/3llw68Wsh7IfX7KEai+APOxst6nFioeX8MhTeYWVaXs9YiF
dqyB2zSb7e+XTbj07jehv2AzwNcZcu2+cmRcA9ofmw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Jz6rr+GL39tsJnHMaaUuNSiQeoU7/B1U/E6Pqoo7E020dqGKmD8GECaZuIRm
Gu4Ed9XTrO89K2GNlxnh3JZhm2jodx9VF3WnoFFpqKOPYyVnVU9fh6wEZcKo
Mj1kv7ntFrZepmm1EmC0uBBQN6yIk1TfdYzzLAjhcD7FzFeb1tI8j/r1RxYk
UXwe8VRIeee9EUqWEqe56SDmiQF8F1hwNp2fwY3VmqIAoD5lktZbCYDatBXm
euCE/DqFlgafE6Hjry+EjtYa+0D+cAvBEqlf9rnRDVZIjRJTwG7VhdAzXC/y
Fa8nBHHPl5BJm9c9FiqJiur6oTF+V6D65xDd7KfnXA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HsN1EVhr76IXtGsdijF/AM0LY0tFt1yT6FMlBgebZdKxTuowgVnonLKB0kXV
ZSjvb6HlOIExlm0h+e0GE6MmnoMoHqPEC2r8+ppahyDhI3k544uoAtTI0Wcb
QbtTnzhZF600AXXAQMwKQfpLtiJroVmObhrc2vFJ8RH0L6XyufJDypYubB5b
/BCVbB5Y9edzm/+SFYHCdMqLyu+XRX5hAOE1zIuvp7WColQ064Hhe4PnQu2r
jgj85B7jqQJOdaQboHCZGm5bx0ExpLbT6K+bwdoYjB+sImnvwM11QgO/Fspx
JmNw5BL0vHmHlUcFPgj7oiVqzLx7gldoug78jzltcg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DsnILuBYj1j8Swae4ijNym5AsYBtnksD5uvBT/oEUe1xRLUwhBs/3OYAUYh9
CDKWRS18U9Ou12tYC+URIJmJTipB0qHpqJjo6y1tOSU19G5+SC6rlYsz/SXv
Jut9iRbO8W3ek9yNwCj+4xFYtN8i1qxpPoFjpYzadhO0r6SegSY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Np9D8AEFvIP1yc1lz30PnlPRNzcVkch+i+JHrjvXOYySG38c0C9rrMoI4Kz3
1Vvy9Wlq79eV22XRxR9fQtZEnv8hjskXW6Vbyi4YbwGw7bxfmjccTDQ1A80r
loJskfEn59zFrG8pAX7edbcKl9eGTAh0cagTSuw+rMXdUxF4NrhdssBXB/p4
mQ8r/8aZoDLLlHNaw+IzRUkpqer0U5ckfgnuTS9p0s9w3k4l7J+fttQlBVug
WSShe5r5kOii0t9Drwb94Gz9sTrwWsF9VSd3w2IctMyWdfDM7MdT8CRzD5CE
DzOjkfkMHUh7dpF8hyrUiBvT+OwSNqxLqG7R+3DiOZIU2SsxQhKdm1yup5RS
Na85nV3w9GdnJ5oLCztIP7oiC5iXjJYYcG3iPgos0dQm0GSFM5dbm1VYPqNz
8r8+2DwsMBSfGx0AEMfv96GUkB8gF4mr1Y7d9Wcsa69cUmPHh66WEZEMTzl1
BQrVj7cKYK8T99PpfHx8/za0iJ2triqF


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eJ/30zzVk/7rvU+fO8y9+lbZ3CqfhP+b2JrH1JLHvBdnQeyQ6qyESKvXfjd0
x0QRdX7V1K+6qm5iQpX3N0izVLd26rePP/crP6BDN3CE8VlgPLD8ZrigqDJr
dZY+lJhuuplC7KTC4bQAiyOB3rxyfGYHAFSgkZ6nvRjUrcodaC0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
f0HSKqgHfkWIdWVDe1/x2oSR2FympOmq8x3zGKyOIfGnLybaxUMd3ViDq5HA
6DHJsyndjBm4/G5fNU+N2/wL6ytPMwXcWOYNnQ/C1+r+4msEBIOzEvrV2IPn
IW7D+dgPRGtRv6YxM0O2D8LCvaUcDNSeOnXM9sTx5KKwdeVPzgs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10272)
`pragma protect data_block
ioaW1GnDCbFKgiXYL6KSZgbgs491w2fcARaoyfgx6KbyKnZu7sG9Jobg017F
YtZNRxegkdKGeRXb2vUQFLX2at2LOIZh4uqEQ13Sak2oYIkjgZFeEoVi61rU
MFCzlEZa+MsvOcbEhWDlghf+bVACUAi4rr0H9U47OhRD3BFQx6WkqYvHTquG
0UHYO0vACb/1560VuDkYJnyZvIQdhQT6wh1Sj8oe5efuNujphvQ64qkZg9pE
XdtIa0m7SucAWVtEcQGFa1R+CO2A2RMJaXfC4lUmxshidqyOZHGSKkZBo05y
tdjxe0ioO4RtV6/EdyNPRn4yfAcuGTtQkVvpON4UHD4beCWl3s0Wyw/A2QB9
UWXg+TLuNXTSSOgY+6Dc5wyQsUjy2CSzUr6G5LuJTCZF0fkO/y9n6ZTNdszs
8NkACUy7uQMoqzqB3O0Ysn7NJnrzDPXn7/9X0ZfeSlDr18vcUlJ0eqs9++d+
6Pv7T9WdbXFkbv6btMILTAvUQgxbN2jomBicGVzWxqjd4KFu7VuySeEFbpOH
CRgy3OCS7RiABzeHds/rdK//iDBx7KmEGRSOqHf+Cm09Si7YlbdJl4Vnt0WA
gspL22PJvfnqDnNWZZ5VnBP2ziIOMrQYE0pray4LdqQhs0SQNc0xOYHlaSR6
I67f+4FFlBGeCOam6ZoeW8FXBRjMrtciMqs1BjsjBA12JyCRr7RZVMNsm+4q
eiowAgHjAcC/tBMB6J70tsOXl42J0WeGb2XiIkU9O3EgEioSJCWSrKXE58Wh
hBgjvc1pEWBIKOggNBomHAVhTyyraDPo6Lp9TajwG9x55R2Q/iu3Y457iAGV
2xEHnJiVh0z2ia4Zja0pChoR9KCS+GckJWf8FQa1dy7U9WLZxylkXYmZ+WW7
T3w37BL+lBpCtfbALu83o6iFhiQkit27eKhcwJUXbwX86DxGqvDAxA1/rDgY
WWXWc5T7qUEBVm7OKX+gEW/QJ4i8XU5jdrS66G/DhmKfouswRf2FAA1y/rrB
EyQtoaKW8b3oH0lbJd9SlMrO823+GbOwJY/4wnukHYwG4TR/vIa574dXOtZv
QKobE96dfKyl5TogVZvEgOuunUKRThehQXR3sArJeJADmPzUz8xQaZ5T444G
p/bhvN3+RUAXU5Y/Dez6jkHq0yIPKAJbCD9myW+4ybkVLzY3gpNq5INo1t4b
p2Vg6zY0f0IE8t8RHWb1qneooCxd/hjgxgRpUe/FtxWCqKs29I8BWkeJjoAX
a5UrD5s1vVUg0JPGWas1UDcosUcH9VHaZfLdssUhlsXKsxF2d81YL5zPQHCr
U6PWUwT2UJSgGskKIQodZ79iaNzgbcBPFIMyK9wBZtMTR5efzNkpfZHKjakw
K37fUYDqDPPCZ4AkJ7Ds1+BjHJbRM0smpwaRZcEeN9JPffG8mPJHcWk+0cVJ
u3RCejQGjM5yrKPtqCgIJD3qelyOYi9vM0CH63upz41v+xLZ5bvJZpTqi4PJ
Ht1wr41YQ3sWq0AWgxKwB9jsFwHb0F8T0bbdTn3XiH7Mm3QXCCdDuaCJJF3J
PY6oAdCVP0bGkFVQhEJtmG0DiZmGuyJC+w5t+NEB1QImFJYAsMboLvE+kEDO
Xyp/48kaD3x1fDjJ/ULh/bt9sy/l17VEZLxiQz+nOW8I/eECKJ9eYyLVBogx
PDubK+ORiOe4FVDXLW2AhoCChuyqhn9MWW4UQUlfMURa3R9dLllJyN8TCnA2
BsjXpA9l0J5NJi8et/O+Oj+wBs1nTCdtPbBPoSTJaor7D79JJo3V+mAlkSaA
E7qCru0zcbuiu5aOMhhFgYqJHMiJKHLH1cmtW5XLcqHB75SDn5OYc331R9XS
gzJkx24ksTTFIWVlkUZ86moDZqMjpRfXdkrNNCld2gsuPR0McEIkD/EQjqSM
P/iEaLJ20z3DO4OpNn5Z2T74UmJ5+yjSXYTNKlWPqw/bHx9JpcYI2B/4JyrV
i1hH7Aflgls9MXluH8KGfwQrBQqgV2fUo/hdHOG26bKX6ZxCS0ObjxvyCwlx
YLyGWLJXMP+qBklMh2rA+tDv4EzlZ4pz7pTuLHJG9g3refkKFIHeFI9MTWul
h55CJ3gNuxtgbP+F8fXqJjHguqXwFhy4MV4wNSUM+CsDFoUu82XIACnmj9jt
Na/PR8IsGYj/aJUO9zlfDtYiXv0n+kCB26Gze7zhmWKUNM/zFWEzf3KYRykN
71HRVRs6JWxdF+j2vOgSgBlyX8GgN0Ua0vQGmRyNB/gUp87XxAfMu8TBInjS
DNxLU6IVFzOmjRZhAwMxMfIF8Au+bseYwkxZADDQbcmhi4KUkJYUtAZ/rZi3
tpRq2iLYg32pAey+OkbdfPg1JTM8FPSo+Pz443nGoT0GkFNvKkrGtI3S+qX9
OXPuATBhq8XXuCdYNU1qqtqsHzojqbqzq8UpMDdwUixG8d08ic102gqaiory
IVFnTPHj0zU8+cH9WpAZd+OOfK86PjAm60muSDvX+4CfZZRZ5TtYg5fiuUvQ
uRj3hDDR05mfar5sK6OxwWK1UOfyI6LUHM/F8dzx3HDiQclnUYyJTsL1S7hV
/2ly4DneWfCfHlzoQm8BcImqsb8zP74Ek7qSIG/YLqhFEq7lz3dBe4eXWNmy
ycZ6Q2yvp6NeAXFK5QAsPgsRyDBELmJFvp5gusZYa7uTRLko6hj6MXd2ofoM
5vzjOK456bY4fkLz0Q5/H/xF9mNGkpRMbsjeeGOGkzvNhrlgWClMnSYskWde
u0FHxKZhMv5PVHOqbPF4VuCaMuVbF4JPjS85lDppv141CKak6wsNW2IT5Tce
bIHXKPiL3qbrTjoHL9oxQCP/KLkHUZxwOD1vZuTixtTlsL9VgNvdaJiINhjm
C4zXIr+8D/e/9j81LMSUMResegHPaaqF+w8+zXpFcOl9Y3C7vaJneE36US+C
NlM2uxLHUKfxqniMad/xtZw3O3qslxGFY1rZ1/A0KX/o3SqfF2D3H1l7RcL+
Q5jPD6yZOil8Pl9/YUCAMI97b+ANPzFXV0XMM7mRghWhf7dWczxg4jGNkTTQ
OYG7uBpJlhZgU5IlXGNXjo98Tb5xpyToZHBJAdLTb1ohNJhq4a8hvnPGzcRA
0Z2aXNEp5Uq+YEaOjCCfqq0uvI/uwclqoeM74quaTlsEXupD8R1ShZ15FZGC
spPxn5ybEwrDrCJbomNfHGvpmSjSltjtYmFsHtrgpEVLYG7Hp7k2aApcav5Y
5Z9duktJ5rFc2HPEmfLjqrKXPYrS74g8WyIZbeLZ8EqpyOJfoshR2P+DhoMT
L6g+KMPZp8MZQxBUVUx+xkT9ilTNNIe/kQKppSW/4pFf2/0u/A9HQZk9+bF3
xdlQeB2ay7BF7MwU8rUCrlFiVD7kxPlj3KBiVuMMcI8ogxFlT8t+SJzd5XVS
ts9UyIYU1XiAjWH1VkiO2Wcq1PzrG7T/N+eSFPT+g1xzu4xXMOHC9ZCCJcs7
2Vl3r0qQKpV2F+8GYrxK6MJditzaZMCVF5mEA3kmidrSABN37l3sVlXLsW6L
E69IPZPtSLMnN8z/KZDkuLxL3iNO8BzvGh3Pz6vMFDHBflsTWh0kozeCfo7c
rPKasnsrbya+VSB0Z7+C2RXp+V+sErhnM9EySFBbSaJgZCjMKqatzpUVBTdx
1AWTayw+Z8suTLm6Ff+RqH85Ur5VHOZTyT10wPCunoz7bP6IKSbSNTy4SZ3F
/jXEtj7Tb4biDFHQnQKPBw+lfAgjYRchlhEQ1iDKDBtDcIC6dSwiaxMHPXNo
vj6F9lDoZdOBCsLKrg8pjkdVVLwXPFkpSS46G+DF6A1XQ9KxbhQYVmYjPYOi
OFHR5tY+LbDu2tiNcRsuacAIqdQn1Y2UpQpNKGUI2HWTqcP+AKBSImHmK23F
wQEK0XSh2WhAeubUUUqIiidcV3LSTPOLLwtpQ16VzRlQkT4oe+U6sRBwqDdp
H5Mv0sTp9jul0jMzr6JkKdP8Cx9EpW/Gml1n28+iZKFXYNpI3+eZF3jZNwoC
X75a48HHF380dOPMaCMmnUk0eWYlPbxrX0b7QdX9kBguBSTri+3ME//WiLXR
sp0JilvyqMb7y8BmA+hL4kAqtTALjopmzjVdS2pGMJh9Wtt8vcltQaEA6IA2
1TB/XQymtBQMoaG7WWNi9dfYnjaiAgECVVYCHdu05AvrM8ao6RggZmL1QSkf
Fhi0HTik51KuNUksjGVYiDQqnZFTylf9RGiUttQrtEdR2eqzw3u4gqG/fr/d
ElMRrUUZtRxjmzmS0TZywCQprOVlQpIHBMdhZdaujgAOBcpjx0PRgyCMpWpt
hExqYPpi0wa3p5MJcoHcnBPrrYt5F8DyR/Wi8pwdLbH+D3Cd7Z6nJv3dZlvV
29JjN13+owWi8WcSHrqsmftZAz3teHC92S3x4zykQi7bviEeDJjqNTUpp31I
dR2od04fE1nKmZz/o7nppVXGf8Oybq6J3wI8MVbPV6XPET7H2a3VvvWMcRSl
orH5A6ClQhxuLkCqL0W1rkFjxJBo7iRR/mP0ED2RVav3OhIX/ewrawBS4/BY
aT3N1c4WQB58ocpZHYedYcLyveqz8PseuyYl15zo2+b5o5PEjvtjgVnjLh/Z
D+9oVK1DdPSSXEAg9ipm2eqS1duQx18cBEMOkXO2pmjJIZevaQdSmEMYDP8d
vjxvgvM5jGGR/M/yQn/RVoH5iFk7a9TF/bFFBzd+WaMUGnBC4u2tI5ogJYSt
WG6MSGK6pBZLQ6/Umc1AqqjfgA2sD8vPq30EE7Al+877erXjdjOJ4n7yyd5w
aId8I/uxgLVk3V2+S+Jv4L42ouZ2v2/XfAWp4QMq9l1Rf4dvtxbxsQZCwa1G
wMqkRw6TlVrdffPfwhTjAYBwmNHg9aU1zWbmv5c+9sQyGfIf/lyXJM+3uO/c
cgnEwkXK4/9AA5FkEKb3C9H5yqXOtXLFM8jjw7Y8YmMcPsXRgNqJ6g37NQMB
TMRpByNF4cjDsj+RRS6Kw8Mx6g+iIkg56uvPqJ4vHVoq1AwzQ0b2nzbtaSoC
FhM5iJB+MTOnJ1WWeGp9oAgYEHzTqz2sf7iX6bvT8z1Cn32bNCCF0uQkgCaA
w1xyDNNNbM26s9VMdNvtKURw9cqh3PiHkddPllxJWDiWT2xl9yfPrB571o/k
LwXIuGgP9U1pKDuJnp4edycikImy3TvB0FI9SxIDYyoTBVy/FnMiDVoutI8N
+nx4zySLdTTlH0ru9aIDG0Ky6L/UDsyb4ibD1PDxsz1nHEEpuFdGfUTKTFWI
fgDRo5lVzGuUygjuIna4gdb9v62flGodKbxoj5TPjXxMErIAf+j7qAkFubyA
NBlILtFl8zxX+ozuzldeL9WHlBZjC8Pj2EH6bBNuZQJ3rChmQToxQwLFOyi2
NWgoU7KNrUnSPVFnEfhAusnTELzP3E176lh7F/7132MVTQ+TGaqfpbCwe4Ip
8Ocr8+HquaqXUw5Arf0tYMa9oNpCvAp8E7gdejcPTv/uxuhEW6KSRHY+PZRI
YHi+9xUSIsWOtuzHlu8Dzk+wba49HMUd+SCKkPqQU9HkaAOb2ahTYxSBo3hZ
EBCKGyJ2R2oI+nrDM4YHXlcxv5qUkoPWQgWkve/NNTZWq8oq4OHKVOhzHiK7
/s+N6F6576PbT2hKbRzbGF/9Arx0b22ejedOp4qyXbQ6rKkF7DlxlUD+6uLY
70NrKtBH5oaQ6JwudvTMRDNqoeRzS3HYNBFx47ZdT1Yv/5BIhBuWQV1zmKs1
ShIdhZ8NtT0/R/1/vXpoIV4AZbPnnULZMyJpHMNuDZwTFLYtEs4BSV07Wf/Y
XOJO/CChnbuwRVkuRlJtTuvNQUJprHyuh5u6jHlEb3VK7+jxk7MQlBfXp2Y9
MLblCtFXEH2UKvi7aEmg02lw9ezPZ/oJixP1l7izYironzZzfmgb51XpabIu
Mol6ilGax7rfydezjpD1a5Li1WRqTrbZkrqn+4ppqvFYYsy25b1cGVUYDCRC
s7qA37l1pxYmOTU1nyczaKLlYzarqbD3IPF3Cu71tU4I8hwfHM9DrbhONQ1W
T7npsHC3xsA/u/qrC7XGleiYOTIv4qVMHQn+GpjpSNAUdigG7FsmRKEImTTi
CO3hGWW5ph9c7VvbI60SXHxc7CYDJaja6i+ZQ7gBsluDiBEYInp3xzEIwiOJ
9SycIwKVE9oEYfJ/5rwfteKywkXQDTFtBhsD8WdzS02L21n3jqk2LA53a7cF
dvdYEI6btWF3ncA5K2vpMF6BxDeBQPiWkZ6Ddza6GQ/fF3YpuZdVYFJ56vzS
Vi6GcOVrTuphlPci9yhYbBI8iVP7bogmvNEyw8CGg439xK8WL96sfibl1FxK
D4vA/V+F+2dzDZDf5wMhZ6uXEkLUaTJsweG7U/NxXCkIiKVqq30UyD7ngjR8
zt2jxUv18BUXrBRp3GZeCACkoXqIhnditcT5PPwASVfmPFS3+N1RKYmKES51
sOsS5Aoee0U+UL0d2cQN6RpvxbFJQLODS5bPCmdrJjkiafp+93dJvv0rwHtF
bouNbcaxCV06zlic1m1O9iU82EVT9IQ6VVTS+V5R+xmdnbmJuBaexhOc3pG0
WdyTs20m9tc6cmzUZiADV2im4UOdgcwZBbhvFOwIUmCWqGOSV1kkKXPbtlVy
K6vi9+LbzacObh01KswA2sh02MWBzpGhgbYxEULeABT1Wgc9mfq/3c07s7uL
MrseSRRHtkwgUdd/b//VBIma/pv6cN1YNYc7mk7J5pxzsDrIW5W30pyR8Ffa
Fx3Y2h7yOayKuT485eqC3aC87euL5J6g83ZplVMQQ7JNJ6frmZEhekcoo6GV
Ie3omY45RVInILjUAj6K8YAmYgq0847mnRm+7/vAe8GTDkqMhrBMuss/JbFL
4i1PAcssD9ZYUV6UpNht8rOUOuQLPOt7zEs/6aNSGj3Lyhm7mkucNZeN1+Hv
kV8/J/yZxQkPMjULvQrSyoXBqnm6G0DtE/Z8QXpsxBFeg97V8fNDUciES9qK
MfqmlJa+/KTqkrETg8K0swweIesFoStumsmGxIAEsYT4RsElXLeRSKUl0eRX
ttssSHnayfLMk9ymq/fKs7KnZKyIAMd8amyDO8SQFe8QSR7CEkxI4WQlR/ik
RslJb9MXAQD+ci/SKu+Hk72Gt3L+1dS9lGqs+VAb+SPMXht0lA9qpWZ59MUh
M2lFWdL/fr7UsW29tEkkurD37Kar3mBZykyR/BRxI0N4dkijXyrXUsuBOx5Z
/j12mrLD7mW0e+Vntzax6Z9AVB9CLG72tWj0So9YH0mU2+ftqNYHxmCOdzKC
A6aenoa/O9EEesrRy4ci3MyU4RoONPlkzfF03kWAxhYl25Dh/Pp6SBZ+AxQh
TjWDYPiyP6L9BOAxvIyajoQKe0FY6JIQqAVpbbYydzG14ceXflrbT8CwGbMR
rHFjRJ1m7F8gdi6TBGYzc1ah5wXyddt+HWQ2bw6q5dBXS5YMVOT/Nn8glkYH
iL1sUX+NKbvFovHtYgFH5KiipWONn8QZOla37KKlEqmnAK9O49LEOVI12pSq
a0gBhensFBFsao//1cGSCjECPrZI2m9WhjjmWyugmCF+sphGBSuZiBwzer9H
eXSk4kkTLmIs+9CNS8RRI81ukrhP2xtgXGchryhYPgudFyQHrSFLaF9NJpsx
mzAr4dIwiPk6Hs/9up2S0+1idq8sOXQq02zMUvTXzlSkOtOqDB6CtD8wBbN9
smolUEdJUU6dQXrqJxaltqQSjgoYNRu1wGyFKn5Mr9YNXRWDawkdNvIKMkFe
Ix/ZzAEkH7Psx0AkvV6fhwretOrt/GU6Y2yI0G0bbjVqSEQfL7JjYT8yvKJZ
Cv1ECwoDYjmQaZaVFTOdb1Sd0GIVMvGXxIv6AFD0v77uLLZ+T5281fELSKa2
6qNEv9/13acTvWGJl60C8J2/8yNoMs1z4QfWdCQCNM1k0qNyYByDkigZZ1FS
Y1OdHIvMlLQmkARtNJ2CbKbKQyhJa/0zx5NJ6c/R1J5Xcf6bFGOqbfiWpSY7
gEjFhZrgoL1uZHCdtSv2S4Q+gyznnCnXlh+0hwpNU1XPLhcMewnXwAmI+g9p
xUKid6xD5wZeWpAvf7kB6rPfg1GJsyh4MNmox+q1rAlgsIadk7OHRuf9t1JO
6Fd24wVtTfAjpd7Ja+axPaPK3Cxi4jCElZ4/v3kUdi0m1fzr8eilb71+iD5r
DuY6MOnVMEw+XB3FOmDcMTcPeeRgiPXFbx6qbVXSnRTvGq3GaJD/IL/lHRDM
YvNaBXm7ifjVFnosmLCl3bYRTKdjkEVlK03WWvEaEvRsM7k0MqIQnT9waiqO
jRuHExJB0sEz71zHFV8J7MtVG5fgDApOZJ8DTWruqs6ZLjbFyXfVG81zr8fA
eq1X7UYxCD8irLOmP2AsNRofrg3Az62bEWNkRs5O1MFApEMMCp0kbUhURlje
jwpXh+iDlWh07Ls6HO7/fOMdO7dCpnC5oft1FrB80kcJuF/Fez0ABbbD8o9p
lzCEz2ZdubmJWicIUc3UAGs1uUAx/SkhCWgGH+6HJBeGPb5rk2S2hxc+j8g7
TDcUkY6/xTxn6E3QUWMbznz4W0x00hwGGVc8/tLT3Mkwa4Na1Et0OO8lOMrs
BGB8zdHHFdfAore5c74iUpASEBZi9txVlzTGc8v4KbpejPF98D29gcdTooR3
ojsNxLN4d4azNw+pME7vEuq/392jL3adzf8rVsyoLSjjBtiF+36+2m9WDb/r
a0G3iLQ6ewUfRAaL3d2KZ+mWqCvOtJS8UQ/zmQB9633rqNR/O01fG59bl6MJ
Zi3oFpTjT9fbBXSPEq+EpKU2W/ktxKvKkV+xM8eZsqJBscrUBxSj3NMjjzv4
XG/5QgJnnm3kuSG9hGtbHAeLWe8+fxwbgEWGZacgaRVS+cvYKYgG5PXxk+me
qn1HNX/Q9VX8lTKghYFfdPZFqFqJoqr2UEz/GD+14Bf9vYYBnR8TdWuM7zWO
WfJklGkxcFhQ/7JzHCX5pG5GC0CnLAFm5vvkemWOKh51PYC3oB6iez1mD9P0
D1xAccph/wHKJbb2pJsq+6SXoKiF3Jbb5K5qcMSt0bMH/GQKEo8vU6R6jubR
VHKXzl8V1FFhZEEHW4APYrPbKOXfUkMkGFTcGwS30Brcg7ZNtyX61PcnTLyt
5iNI4hpj4MDrnnXuBSHMPspP1XtkhBpdB9hxe2O4xehMtcfYew2q6pet0oLv
IjC0bGAR8aONGG6/Op/GHqcKFsEGIyXAyEKsMnV8PRWtXxZz6gMv0F4TkR3S
YrqG0NXGDsETbWhf7jfxgrHkftro6p1QQ+8mvwooiWjooQ5PEKzUYojAqt45
LmhhH+3d8jJ349HSCSZsMf5UN1j4pIMpFVHvM4V/o+jT8mG6vsy7GxGOQULQ
ugkmPH6PnFUw6cV7Zq2gfRK9Cr+Zj65JMT7hx+tX3NTXAITqyvnCt698OrQ/
NLNrVK2vFGWHzunIfUT8xK2n8SLcEOVzohhFPkuIxlTvS9S1J0z67wlLA8PZ
m8d6NH234I8Ur+lTMzeRwv4x9k42WfBN+1kZ/pHCdpZtQ1R6eLNVZ0d45yo9
GpAgzZo+a2xHBjDZ1kt9crg7u9k4JcZc/EQfSJHY+KW3FdUeCnW1AVrVkkE3
FcMcwzkrqGTMizAXFGwxOZ1jE3/iSZhVA4IX/fW8yjcOuE0pV0H62RfI4uqr
YtwAUEmoK8rY7a+wqP7bXpn2Ux0XK2ij0PJT1HR7qNHUQk3BHCzsP1Z/nErE
+b55Q0YekxOrFNUq0UOtZN9lDPytldaYROfdWXk6RkeTKNxLqEVfnvg8b8Gy
sPYCbpKQahEA/fr7EPnOpRc2U9vJV+Zg6zbRSzii0k1w54Yzbev+M8re80LJ
y8ma8idR22ey3GQYbjZ2CmCNaq1caJiB1ls051FxspilhinIAwZQnfGYCTCQ
FdzOizBNzPzwiFgkp3Hm7DRflZm99U7In0BJRd1MWZq3PWdmRVa/RZG3JGMI
O3ToM0wva0Jws2DmAyjPBbWsSWP2cQEydvTRMpBY2eNFDKJ2eamHWBbcYlDr
7OKZb3UlNy9MMFCllSQprkTiRMTYWCSXcvd/sV9qt39Ydl3mIw7VR7Ikld12
KhvGgwdAygm8HPSrin3QV5s3eD50GZQpIN0qKshiPn3Uta0uYnsN5FE1gs7l
fhmk8iLdEzerpmIj6MhvUmugVRxfV/X48BdPMyiAWizJMGxKD+mZSZhGFKZp
VGhcZUTLnkn2adPvvFDFVb24HkyHG3r9xCBlPevXue8pRFMbQqlUoH3PikQ4
0tWt32cUG/GIkHPnlW/AS66pmnX16I76aw7ny8XHjhcAlgUhfyFHBfRH8zSY
YszkvqAnBNOD0IqsJo2qI0MKVdFN8/OQtsu6SCVYw6lsy0SJacRqW8u7Y08K
xZ2GYfMD5cdjKToFEV9w0HDxoerAlVasspv6eMu4VSGfMxlS5yyuXdww/odx
ArfP7/i4oRHxT6rpNx1QhPqIuPO16E0MBS6kyq22xTywbNFZkvOAQ5fbu8QT
mgORYJ4c6k4M2eKwTvt4KtokwfpqgE/5EB02xQzd/APMtEnH0G7+Q+BZievw
dGgAysJOHsWKBtdeJ4bIbenbCsYM4GWsT6pH/6JGfxskjcD5aoxn4b5TM/xR
vxLWTpJ9EFDnAVHbzo8PNzB1Xq0zNO0XaQF91d3r/Djky/n5AXQxtNc8ij/4
QxOA/RGekIqIPWQTfd9SQC2+9Sap0bmRsQ6Pr5S+9ps+8YEkx3vra5V3ZzI/
gfzmEevbKD84TOs+gcbIs2RDWOjw6VA6pKhqQoAon3cUNDQH83rmRh+nmmbV
dsUlH4+MYaPCFut31bL0bwzxhzB2E+6jHzR36iDjJsuIHQJpLDBS5ta6K1+Q
CSWjnoqC/PlfrJB78yNZOrLx9lWVcklev+Om1rW9Pj58QoP6gNw7uHaZE5JE
EL/gFgEqhPfsfX/b+l7Vp1oeKTWNePR9E7lrH3fzcwcHHalh/E1A+tg6GgoD
RIxs+OTNdsECDLTqPAFN+tZpv4I3KjR3FvqbeYlfkYGsZSa+QTLgU/bK6PHt
HkJb9f6yMWA+rP83zooi/4OWaKNzA9yR5kslGPMjgq769jsmvWMH2JcgiqLm
YbCxZfpjaBRZtNniwYeTsn09j+xYR+QBI8dNNHYxzOBNlYvCn3QvAaZToGUj
/7jaQC5SNSvkKcJ2QNXPevtug/SVVc0CVA8KYWYkrWAQbExV/MbeEnI4u6AH
Cog7K8CXWJqrca6Sqn5neX1yzrSpgorYIzo7gbtrtVOP9Q7oPShPCwMlTo9J
1v+Bpvxox1nkInVRuAX6fsLDc91/7rDShBXi9murLeXmAoCqGP/XVkIC7Z5V
QTF9Q4r3GdV2ljn5G8EVClwDnThTOxw3D+sECbBXtwEOhJdWydpa4E4m7gcc
lQZgaz+hfo88qQeAEnUv5XPvN9DM12yb7mQ+cJPo2alD+PxrAcKGKdXXOH7M
zmpBbSZfy2oqh66x51d0ZDRb9OODuA7r/bqD3zDof7fUkhV+CVhaSWiM3Drg
K8ZizsUzfoXADAzY4w/FF+dGAgohn1olAoJKtHnNozFBhodYqkFsnqtC8Phv
1PA0H9xkoHw1C8zUSKheu5SK2dphPDEzbrWZII/t73bZ7RPWqW8ixEFgqp1O
Op1E0/ZZOZiOfVONUzRYm3kQfZImLGBaFL6Dz6i6vETgtin/b0hpl2QqaHBB
/PCVg0wY2EyqMHSXlYUsU3qe26nxzrabggny9cuM0zBR5CVjC6BdWE9hIoTj
FD4QFHT9ubxr5YcfSINc4pvTjlcjwIUrS5+jhiAL6CEeJXo2qHUNxjzKTDaG
NqxEaAKDtznc9kL+g0pMcLjnxZHFl/U0JRviSugpuSN1S1CCliDc+1iqk+BI
uB9FqwAe9XVHqqcSu9Uso7Yo2yWZWsxzxTJ7nsct1a6kDbI1MaDrmc12w6c+
sxnmAGlJiU9fnP3D0o29EBU6IPrEzGFlwtCwokMY6y1zFW5m+v4SajElQTO3
3bPiuX0qB4ArDDhHQlQkzsZAUhM9plYQGmhby6deshhLY17wh2RKreqpiMky
++CWX7RqmvmvrIUymJOHSio31o5eNsCz7UcF+S1fTVCTTcoGIIV1e1W7VROM
7xa0zlUUDV4ttMaI9CuGqhb77pZj58OhS2QSR+EFUP3A7zRG6ykPE3IUEmVH
6WIbcQs9hAoyCSCdLujsr4fxD7rpEniXSnfk/gifrZHVe+A0qiCE7Dp6nlWg
vEyp3Pm/MdWzzrXWhrBtwsJ/sZjIExY6FcySyXO+eR3P01PGHJUkJ4zU/DSq
68needVYK18mSjwSRVCtvYZNagmnvbxnRgef7Ynx1M9cXX//iRM+ME14mSNQ
24Uk5DHo40pOtErMX9MseSFmQSarBOEJ5WjF51zYLp/3eC9GAVB4Mu+WCc37
KWp+gz+ieFi55t1EZtK3KqW13yeeWmpRDcPEzKneq1AItqgO7aLwHwgfho0M
24yEDBwcYChF41PUNWx+TirpXhT4WOcfu7gQa4/oKaZbO7ziXtkGp3GPGaPj
T+MKbySbF2ApKHiGwgc6s2y8qn3Y7nBCbdAkjOthfBiEVOBcpa2I5HtE47WG
8A3W5naU4R3bT5XKeqZr0SQpizRtv9T8dhsazNPK33Pg/sKt9vY4ueyOzmNS
OnPRtjniYI8suA5fHqxOpggKKRRo86cRm/p1kn4KMF6Whfyc7WkaiQx7kG4t
h3JpLOqFD2U7vsF1uEwj2yf8ZVGVFdURtjhEdqo7Ld9v+6MU5eZIDWopOlUh
XP1rKPa9lo4Dspii22zpmZKuzlWFxyUV+qiEP6OAyuLX0D0YXD7Lhu3rgKT+
wvz+4gk3ysm0pYtGDNAAl4lizxvQu/bHzt0Zm06erXukHJjJbWYa4vbZd5DF
pmMtUracj5XLXn6KeaNMf2Sw7OrHa3+l93OeHTHUdq1LWkEK2VP8E/QD/+I8
hjzKjPtIpjHHX8Ut+YvC7tu/zIDaZJNxZ8OjwLto8STAtA7Kd3QXrmdPFtwb
CByXz7uywbtiI9h4BlzOVvQ6jZoWWNQjD08wQ9G0IH5p6jShpv71ZsuEL30n
zf31Y+KVSak4oZ4ZtlnCszyZlGBnDv3HDxjjjnfv97G1fcGacYSA1o3dhKU0
3SrL+U1mDLMtScITQEb43bIq4UaGek1ipKybWdXYItt9b2LPMcEg7Da4DLnY
Q7+g+iVd475p99dANe4QqNQXzHwSZO+tBJPQgKpDY9rZthyvOJ/WQh3o+RF0
eyDf4xt80f5uBFhhF6KzxNcTwce25m3AIaki5NDb/d1hxX8X2AHb63hjM4De
7Wn1oDvempndN4PsyOayFOT68CkrgTnfdCuVrjJiSGAQ5c5s4eO67h10LsxK
eGJ717COP33/sxbL9GzWwLmUsS98xJWlCJ5zWGqkfbSbUJ5BWXiRv3tXU9U1
xIO+yaFY6BTXwcZM8Ro72lb29aC/6NRL9+eBrf9YrcXmAZ9gRPAuGkq4WtuO
x8og0lc0xHx9u7OWOiM9RNTCGzUQ7MDOpGf1KgfN3ro7UZrTvT5WleNfkvAz
PLxj1ld71rXhpJvRj7JrO0B5Tg4AxAjs4I0QUIp+cuKb0+TCvsXS91wZAQ1S
I7wNCYSDh1qoBdAV

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qTw544HWFlZ/lcbv9tSjBueTBQw7msKFsUeP9dfr/xG+AExY+CaWtceLqvr4zgUhHi+fPSULGr8eAi3joxaW3yh2NWYGVBM0TnZPnVwCrpSepXdgLAF11mvFUuwNLL5+6CyANq/A1fRj67+ZJtWv965MZ+rNlTZM7rZSZXijVj1qOrGwB8DMJo5r5HSaFHcz3hvdHtu728Njm9OfOwpqbrT3e3oFemMqUN17/CDFP3LAVnT0VsKcRVvWOfM6hN7WsAXm8CLyl3UHmSz70/cDFqov+H9vljIoeq2quWQwM4Y3xKHQwn9y76ayU/ggC7XY8kxE2FsAHIpVvnvyGDmq+NxyAXpIPIIGUttilk9BuMy2RJIfKJqMAzM7JfTguli4lKQaeUdi6WAYNaoWSmR21V7S8+lQTaqb5Nt1tsnJCna+0JgnnmG4jSqYyd4BYqaeQb6H1+/atgYjCetHMcmWakCVqqHHyowqjN32YoH0QbiBuH44eWW05yfbilJO+LQx87PunzmMz4Rvpm5diJwqFZVCTVl2gZ+Et1bdDE2Gl0ypERp1G9yWXSDe61QG+FsTiNepTjlszkxoV+y1uNiHeY3ESV0d/SFjXDsc3/6vNF2debCUV7qXwCqxPCNx67/gx8BFwnNLToE+UBMGMsQuMoKRK62n1IiyPV2x25xC8uSpChHtOkVDEhXTLUS4mNrQ3nJi9L4eiG4OxNFSZ4+x3incuyixdrZ+tVuLaHBRmesieplkNlJQtmNlO/1vO3zaIOKm4xNW1J1q9T2T6zCAc8d"
`endif