// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nWkv0sLodcE6GJURrsjGVOgVUE+Ql+Wd1McWtUS1Oi96IHQJxeJQxy351UYQ
lVuYtycLKShloqED6cPh8026rqLObMF3Vh3OSk3/OuvmINbTVlAP552E8YUS
K+0jqlnqBVFNI4frJ8Nxdd+9D5/cCHpf+Mrq2UwwZWkvymH5ZMaqYV8ZXwMQ
OtWk9bWGH/RwDBeUvEzdRalhJQwMkcm8GXMJXe3ba6MRAhJqQtH8sG/BzesM
YOttggY6nP2oV7frYSLDD63PjF7hREp27/9Ey49GWffSPwd6WYrc5Ft7Gzop
ijDVlSI1jApk6g92CTEwS8FXezcracmafc2DP/dNRA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qyrQ5VF38fGmCxrVtnFvb+tOYuBJnqjwtPFfSNtFk+ubghoWjv5751skJ7TB
NbDHNOnt7tZy4iwXpeAWjH5HzIx1FWAfepWPtdpkZbij7+jMqp4E1PUYfdLQ
K/rWGdmUAptVv96rw/h+iFzPiSk6Bwl9B3Zr9si/YD8jqGQ4x+GVjgGIjyjv
wubvCUTqc5xAgBUnzJtfhFrNxOwpL9g7HEif8u1IyLZa35jLPSarzobIekR0
VE4SsD9YCwvW8L4S4Fs+ddglBw5+n5bw3IVolFXPTRoRsB2Y6qbOujVb1nUa
GrwEnga4KM5XZZX+/EvCGEq8chv9b5dz+kK5iyfPhw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iE4Ewxyv8mu3Tb4ngjngM+zLT2QmXMQs7R63qV0CEXOx+Qk73LhYkuOrgyDK
d5hAfCtFasroPbNdjKUxdY7UhqQbcT7zJ/RknGqFa2mk+Trk433uTOtk6AbC
Z9awFbdrtbO7xkpBpPjuC18h0s57tAnTAof9iGh0vcx8gn0mVPax1GmlkBJI
ioL8gnsm/0VjmPn8jp5MPOPOFh5t4oZ0UMo8cdObeb/0m5hT5EF5JDvkqiKe
b/VtUz6FnrhMI76m5A212H0b2CIvM0ZPLu9YZPYncfwQklBiJmyKEVwIPZWK
vp6Ziungpz7b7eixecUJChr8Et301HLruAiD7Be30w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rYKL7TOcPVMk8E6QjujNiVpDX2Oig91xIj0Oj2rROow59EHGzV3g58XtSr/4
UPGYRp7ilxW2Z6vhSgKOBB/Vr9hZnFvDk9wx7a7F2CNLJBYtwYqnkSKM1HJK
HB3dfFlZdeutFNl7s8HzaLS6REliEjwGu+Ani+WXSqqy2MaWQ672rARf1vUG
vO8m331uU3tRO97M6aLNxu7ZhoN/tjtCqW5rgZYLYUN60Dj9ybz+ndrsgCUc
fq5fZcT+S77+nCyAfvMpYrSKHJj3JjUPg0lTqJjuVdFti04+AQEdYU2O66aH
VPWSXroRNxIwfpH6WXA6nAMyYDa73l1LrtW6gUM0WQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iQbvATR4Y8UxFRu/F2yCJWEv4ydNSODfVmlo/cGbWWpmOeYloxivITP2DzFO
XIO+4PLfXzw+xiIW5s5l3oj5fOGCjoS82uQSkW/S4RPQIkS2AqtVF0Z+E0va
EelZ5U7u1u/yz4WeLM8Ub7VspEdWZKO8cgfzB+MeH7AfOy+3dhE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
euPoBjbUpXU8Ar5yVg3Qu4Y4iZ2unOY0tDzn4wq1H+HjEQM3C5q6NkG6VvXr
MtLh106K1Avr8XThODnFPFX+rApQAMJv8o435+ok6vGGqev7bGFdqKOCYh41
/NfoMbZfs1XdVaj97VtoqeIQPFGgxyh6kHPajSPdL3xxrMFrgCYjYz5RU9MO
yZYcMvrLUaiKi2Bjd8w+3gx30thY7r6nqHndd7/l3BsutTn+6freMP1tlEg3
lzurS2iX6thAMg8+S62T1zr7RixntC8AYi9jefjOBTgy4kTWS6tgbiwfn2pd
saL0qcWMWH+XWEYNhw+anwMGmm0v3VAxQ/yBJMcIgl8ArqqD6W5a+Xoo843A
rKlyMsFUXAUa9wnPu0UpYjukj6jRurnumw7XE4IYp5Ad5FadFiaw9IN9Qtwx
KypripGnlN6e9+j8CF2aIQtpstAGYuFtO01XmAtyxBF4zuOEssR1Qjs/gTSf
76Au7c4DDSi1LWwf+XZIQMChf4X8M206


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kS0YWSVF6+X4MJnhIT3Jg6yYyrhnwYbPuPY1pz4T6fXqpqCKKaG8/bioIOZ+
AMt6OVKObgzmjjhvRDJuE7eBp+FfuNxYBkrIUth6NZfLKyvOv/DMjxqq6zzw
LYmiiukwOXnwsaOm0a4pC9tL9xwQsBIKfyA21GBF01pjSbulhoE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gSY2jKAzUcmS1FFJY9rofS8UP3rthaui3DrG5KCR26iqVdIC9uOX+CvMt2nc
6fnJTnkHEBxk2yfhZKTnlP/Lf8R0kwZTT81OxAyHO7b1lYPeIARJD3PKECZs
3uck9PExVeOgo6xkfudXkvKazs3l9bRwIDwVuYuA2L4aicWihnI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 21472)
`pragma protect data_block
PbiIH6k+Cx04N2EnxDp/kn5WSkrJ93uiwPKCmdhvyi7iMrAj34or626GRJQt
9LSw4UaLgORBLQ7L9ENhMp9Xwq3yCa4wwjk3XIDUI08qIkSAAuk44kvYQZfC
PInF1JOGD54xRAV18gUdhwjqn6YAjvOp8ycFbjzWP4frbE/sX2LiI4MqaoJb
RCbVjIk0okB3y/6sk50ZUyl7JmEA/Y33w6Mr2jjsSEYjYptXYdKiTSq3DFy+
94R3poBLMf342An25JgT3cg8Ua/IEXGW0akNwdPfbos2npntLknpDJsUDiam
J5UIp9KAByIQW0Cf5CDZE16A1EVISYpMaFcOJICwlMBi/z0+DiDymvhqrckM
O/zWx5U9Ywy2BIZZck5xsBbsGtanV8L6jk/kh2TAX7nO1mOX2ksi3KGnIxvp
/1dI6uj+EHysqYWywpVzUdzqmOi9wye5DplyAwYEWd0pPBPBownMGK8IikhT
9wnlbdRHN9N9d1eC1xHK5kijlRMq/1tIUznynpkwMCp4GMmafQbogJXEvkgA
QwzUZU45tBdNDjSoKXl35pj+sU4aYwRhYvK3qWmbsHEVP4/3LagY1MBADGFG
D3pUys97MRyyJWQUaFVVkqaWRKB5eqVM7j7u+0wN69sc/1/14r3Q7yEiAuH0
0RRjJy8jBPvKkkBGZ0GASc5i9LEzi7i8DEHNq+TUR4TpUES+LzNSDkK1zGga
G9QVPONFD0dnCk+4ntODhv1OxjSB87np7lyWkuCfkstYv0ZGTi4F4WnmHC4O
IoS7QNULJ9DMsFjL8/kM0dQ/7fJQTfK50nuGAckA+7sMQkQzXj3Qfyaj/U30
LPqNgpRptYH4MOHfxJVpWB+JXWWhuHpMH5RBcXZuKrmhUVqdox8bOzPWE39X
GcHSkjKV5b58dQtTSNkoU1sW76mlHBXzP2hxHv2paGHO/H0MznpXzMYHrN13
cAcsMY7chwwLhcWRi0D/DLZMc+T5kTUA4DzXWoWhe7fo19wXlyZJz5I+f7d/
pCnKJsKLWBzmXAmpMDX3Uicv7sZTfVCbqjB74DXmJO3vNUbgCbhE4slkpSKE
MqvCy2rjFixCVoOjmZe+XXZi5GWO4n7gqkBWOT8WQcbHOZzrjiSfa//fL+7p
+dN5D1rjvnGq9LSkwXBP/iyEta4oWyFudA3OMRGqTrW6pTuPQNRtyuGh3NUT
16sLCWrge26jl0lxeJOHQ0uwONEkP+EjUV/KgD5OPE09W9SyI8Umq8k0EIz0
tdt3bZ0Z/34tN9L9fLKAjU73TMMw9IXJjhcDQDk+tdw09kxCQ07IoGHbSekj
YBu8HP/jQIx6ljM7Dnmu1GUqUrNBgMWkC/I14XlWPJIRBfiEbk7UH0hwMprR
AH+8O5G2P6lIDKYnk778We/hg/8NEN9rmQpKwim8PtWaJ7Xl/hGlHnqoi4bJ
teXxHDDjagh8s4g8CiyAwN37y7cYhR2Zz/IDhAgoArDKlh5GFLidR+VqYyuI
4HJ4xbp7rkZ31uyCrGa/8sIHwRRlfw4Bv3e7/Uv4SxCuk23gyQHSTLq/rjbR
unfMb1M2xHh0FTMiq7ivY/4/ZKJjj0WhscMQN+IPLtBLOs6DupTtHEdPgzBw
Xq7AblVBRea7fN3gIKF7NwUEpSJTz91MpgJS/LpEyciwzIBsNiIs4iOXkhkH
gYcpUm74fVA4EMnO02RJEFDyw8GytW4XBGhl/q09hnlbt7tvjDSB8ArQJNpt
lpxNXK3/9DB35Pbv/FOL+3+S1HSOIBjFesGu9lN1uhZGFT4qpwVgcWbvZAdq
5RYKKkVnMTE8QpwwfOFblXTl+itQIr8Kj3UUzo/3RixfSDO60ycS4thOu2BG
sgSifLpEonTWCUdZ01Ed2vUz7zmXulE37dASUX6yYSE/rgBvNMSyNo0Q7BPl
7SsMx7vtJL7TUkPDZreHJP8BYnzeLJjQo5upbGNz4bZagVKwr24h2zEl7dif
48At7Bmk1YLoh9RAFyAYM+IVIPT4ru54q6ol3sk+sZRSIPzlbT1BfKNeoFJ8
yxvKwivHZ/SQNOtJivGpq/WHBgQ3xjGHwkixCkSyaGIAOeq/nvnLTB1Nq1mf
o9P7Yy0F3gal319fqqtmZjxzjsw2EAEqjEn0JcLu2uTc/UXnh+CW1rowxuOl
Ua0SfkAmqcmwXpBXm7EQVsZXq2EyU/VZSmACK7T4PvZEEe0C3gHmWFZvtmxs
I1gVIwK74tn5vWTlCE2mSGx5X1UayFENYNwOk/j5qx7N7YzdDK4Ke0QDj/0s
iHJnv9EjqNp5JmMxsc/pfpUbiPiFBeGJYjMUJhcUTqKrdPaYs0x0jG0ZnN1Q
VCZvnpN9IDZoGohwxqFZOzKaa1A330kGqsx9FghXi0xMAJjhAS/nitpYwzWJ
w0qzQxg4UHa/avhv0jzF6QX9MOgGmDVyfVzFhMp68MLQGVfvBmkOZC5ksA39
wnGIEojl0apkH1sMf/f99scqXSnIoCYmKqIj5vwHCwMJtThcT9xpdEJ0tRWs
OOW31XcQf5DDzEn1WlJ8nq4yFF+8uIti8lHDJIrXfVZZcOqO54Xg+yyq0zri
A8ambFncK4x4sofj8LbDzWn9kNrFQ1842up7qa7kV/4nlasW58vEbkExg8+2
CtEzyCJdDpvhar8r1dxFIu3npq02Jc/NHoD41jrkA7dIG0QRM6JDE/uHH3ap
G1b5EkOy5ErIaCaLcJSp8uCatcYnWXh4Orc+ETz+ll4mB/eB1tize9yWJKN5
wG2MxAnqLC40tChIXXZA/Pjjb+C38Ek+c7ECRfDR4eTvzM5t7uA6prh4jQU8
HA/WxU1NLusDmFoUcMfh91uPgJLm6swM7RA9iZel2UhPybg9soV9sS/QTc1M
+uKjgvFJA3j1++S6FHdk33yEPsoY4QnqKAC3dtCSEAU+U9aTR+DWlV7ailF5
ymEoEIBXb9z12iLBRIMTlCgL7Vz/lqIJdTCWpVAoZ6P+thSI9wh1kkzFcUq4
QuD9enWOzIHSDgx3flG5wOkfP5MFjETsyS+bQmPSUrlBbbTujRY64NPVP4sZ
Wm7khXl2i3iNC4rWbxCdzeNXMJgTsHDNbaKyQbqkKHRx5VDBVrb9zKijDGNl
kRkB81wQeEvU9XQiuKak80AfGVL2Re26YQ/4yaJAGerW1OwJFJwSBxid4YLk
VvX5RwaceMJIT0kckHz6vxomrgsPkv+wTrTqgCN8a9Biy+OAei61ZRqP0J4G
CsFHhOiVxu2qORG5gxTl+rqVZd90OQr0JMwgDvoWSv+YOwnsQzZnLPEJkgJd
1HvuEvY9peELEAmm+Q8U1nMU8b36ai4bfXiBs56A1ZIFMYPD0lHiNGTiKwAB
OYsKoGLPKHtjuzMBWkLR5pwezVUXP0cACJJcT+g9jTsApv6EmM0byJElhYax
3iJm6iMlxAnQYDJ/jV2o0ciVqgqo4LYjv71P/lHNGWtTrE3f7NGTQzFv0b4K
/y2TSv9MOsU6c6RwOGrzauoD9N/S1qy0YflPjh7EsxvNL6DbJh8l3DLSu9Ks
8SbpnB7A7KgT2stSVAPOJj1wjiLjKX56mGG9U5yo5qd/RTvVqA5EOzNFF4E5
4E0Ne1xBfBGSYaiiXCmmLZJoNkrSS9d/tO8vB2rVceWFx8xxTFkGPcL1ofVM
6IuzsxinUejK9g8y/Z85Bnkyh+gLRlYgXA6+w/dveawOuJwBn4JPk+r33hII
I6VipXkR4FQeT3Y4vfptYVsrzY5byx5qtTzqQ+RfplFv+KdfDGREeifTQKtE
48hrvjAL/QaZH7CcXToZIhMsvxHWQVe+zjhMpdg//U1J3nue+IRodWa2AdqS
1g8x27D/XwTLri8ypxjZpIPWG+eGu6SubQdwzd0f4rWOnvawx1uULB9zhYz7
SoYXCNbgaoJiIKcWz0wObyJiLNtRHUAg/TJU41IQZm+v1vId/TxFyE1sYyeO
6CAlfsrn6gY7L/TbmGGQv5Cy57lCf7wTYIjTaulUOtP8fDyQ/FW+nwyuWxxv
BRoIGMlvI8nk6p+F5cupCyTGiKwxA6yF1O4+w7Z8dkIK/6Fgx+7A3jldbM3m
QDQoBJtvnf+gJxSc6OAis6DcJv4tcX/OVFz5RI+yg13em3ju8Lfc/vjuhOPy
SIyxpTwj6jfRXui7+Gdc7DG+hct9EUaappBcA4L+A0lcg23QUiy2Ln4XjPej
5P5W52vO/Vo4z9gB2DgZJrMHhqK0kzftzs+H0sV/kg8DciDTnMZDkU8rWyq9
hbhzvQd1C6ykRClWhSajMm+Bgi1r1ctqK+9hPaa9Cr7Joj0Jt2wkfoqyK1h1
Busx8/dAqGNHeAaBPVkGdFyjAW/Gpb5hGdQXPNgSCS1EUZirWlkxNCMjhG6k
3SUpgh6tXCyMEpUA/lx+vUFwg9I7p0M0N7LQcPdh8No9xfUjNXbLe5iLBEOS
hVyvcdymSoMoVSvv0n5nt2JyM4aPNJKvfHcsW0bwXezijfWrZNyqOmLLReL9
YS4UZf0+z3pfjwbHnAe1Ui+yZIpcpbRJnulWp9FvlE9I3GORD1ud897fhplQ
eezbKwuLZk8Sq5NwY5hXUtyrRhfFg8xzUKB/0mGINNhPiHH5qD7vSpM6nYJl
e8LbUE6v846+Quuqn3hOZztb21WKMuKLzMhv9YpLV5n1INS+9Lxuzj7AbdfA
KPV8g2NlnqqYDuD76UvFtTyGWZfBpgH6yIbmx5Xy+Lk49TS4lNBjYZwlHovy
74hfgfqt+ae2vNd0C3gQiiTnxWd8f7CWgW3ipr1dqB4eq+AfueeKe39NvU95
UXAPnzoYKENGpmMwfb5kqWWwy4Tuja0XOefgWDR+7sBOEzRPDI69tO2HJ6u7
wxF/2WHcQ6ioVSDODAtkfpbQD+aaSK3pPTfrakVPZF2JD3fGbM6kLU++eqdN
SLxmePvg62+VKJRyT3PfQ7H8S4T2ALk//Q/zAb1rZqS8JGIC7FedO0lGMqhm
Fg7zbZnmMiW/a10deP7EnAAFwX7CPuHbqdjt3HphfTp9fRW2FyQRnVzbE/F7
A7YKOt5ipTnOJcZuTOd+ar+k8n2eQ3xDz8qjEmI0KG/MZ/GJRLLXxrhMeizj
lKaBaAEwP+TP34uGztrqriCug8uylggfREmRFx4P0DSGMl7iXKpfSYZFBDWJ
AOOjNy9zpwoSoBFlqmUZmtdWSoVSXe9X3D5KDPO7E44x4L6AwUOZAlu09R7h
2hQ5BksQbtwRDvLQUeS7+wn58tF272YE6WOj52yyN0qnSggtH1JPCeutNKa8
KX6h1UVuYszjQEVlUsPWj/ghkec5naacYd0ItHRNHi1BpJRut9QTCDZOB/t8
90MhmK4HH07XIMtIS94Emq7imfi+xKQOZtPqZFLoJfNavZe1QI5ot+5RKnGZ
YrLjiSXr7CJi3fA0zxq+4yZL8Bbbs8IUdf2m0UM3wQcHPIQFl3ePt8iDaBrK
EUfJGzuVTP3YHGR1eSgl5XyFwFp2AJpf8a7nNFZUPdjI2fAwMlNJWkLWKhSk
9mUcFRteXwemNn4CbHBFV8cBs9ynah0qYeZsqxVkrCKSlZJWoHwWb1VZpgih
z2rwRlkcpKuFYL2vAjcz+DN+o32GUIKJ/feoiKO1jN43PoUs6Mh9SgQaF3+S
rOF4V7jdfGF75mU5L03a05M6/ucU2JgfyJ3fm2a33TjPE3AuJSzD8qfl4hfp
bOGjqgzkgKEB9csixElFRytP0XG+x7qiFU49+HpNjdNlcnNUASeeVMKAN6tL
ztSAbh/1iq8UQc0W36p855+JcdzUv2mTGAftJ8HVUHLYPK8nodya/UCa9CFt
KReYFkTLbZDYp9r87HhHkjrqVLSifGaxQVzsU7lAip7a9K8h+Pxu4998HhX7
XSiG2hbqem/3yscKfSt+NmVXmArphJBdqfoHkh4ydQqjlgc9B0ucUCAb0nG1
ohIIBQJKL8UOgA0WTHK9nfcqGYfaDvy+zOceDhlHi9WJPcz32mX3rCtHUK35
2IXrM9mPE8LQ9AgedttAtTYTMdr97uBxVdRXM2Ag2shP38lvNaxrFF3ocCWR
fR+Msr9EcHsSrLedng7WEoLEUfQvWWdtya4REFoqduo9cFeIHGUEieifaLwo
n703Ocp3dPpxNg1sPnhn+uWTLgn0YTQKJNP3SgTwy4HW/K6BsV3xrwJZuLG3
LD+9SZavIDpfUi9pZ2pLNya1oaqhJTVj7UuF+hJO33JIfPJ8nRWjyHDrhPRy
4yoj8yWuv3nyq/XbOJWc+Wk5AON3rkpMM/nJ0lqIdELAcZY+PaBTrHGg2DCC
Ii4HXtnjLkGtKvf+XZbC1F+as7f1OXvBRx5TCj/W1/LLNssHtTfOAzdUSZcp
lJJWRcL/9gQpsskxhopWxGuJHG/Kr9TsWeimQD01Choi1+KNXwbPg7x/JTnA
ghGz8k7Fa2SRG++FuGUrL09n2kIt9pszvyv9ag3U52Vr8ON6y3P8hwNGHpK9
JEgyFyalxzLVx743/aJO9VrZ24JrHuBlV9aF++QF1FegC73Gc46Grkf40Hq8
tXt4yXMNyv0CsJtn7aizOgwfCXuRGuMXJiCa9b0GHX3RaNG2fgtvd7czg/Mr
8Iemx+h+bgpCG0GMbS3g6SJi65P3oYsUyHrj9MYsWg+uDNk9uI2+OMuvpsOC
7wno0ZC+Og9m+6kjKdu1udknEl/Im5krLYBSaZ/bhaewMLbn9rDkC4wlJjrk
fP8JbwiHfZ130SDZ8TcrHgOd9hKQOsQ8gg+8HwHa2eZwMp8a3IqWJRkNSTc2
/xBwor5us6NpXFvKG8arAnH4j6SCiifJH6lx4yhsdJDbwgwQZh8wNxaZCjvo
avkUeceGGZVD8V7JTb3tlkj2knrO+aM1gKj84R88ZICZYqtk5arzlYTpDm81
1qqciiiSoAk3bf39FOS+BsPcdk3DyKl5LV2fCQi36YBPfhk7r2g2cXHC4jfL
SsPPnja5r8J4akt2bpdgUbAxBZMSiH/W3xKUM9HhyoqRjN67jd9B8zYsFWW5
qOJ9E+7HzArJtvsJloh6fZ4w30V2JYtyDMc7Qia7+mSJLBBUDlC4TEdq32OA
4X+WjOwR9WDWR3d8gL2MYAlZ+S6ZNOgiYoz86VWpRyScqZhJZfoucWn4hYpV
kzCF5x3E3cTAIogKLbXdJUbJhN8FrypIu04CsC6AUjIyGM3DcRNZq+BSx9IB
D/FzJh6+/oN9xNovcbbfQ047/jV4o+IRGASWJokn/cD/E4CaHJ3xjbTTSqYp
c+q8jyUFbIQhQAp7hyPX+eU6ZsnXPGQrRD+aQ3f9SIxWOYArHBiA6YTJY1vX
hvnsU/AxePlTjvGWRI0z7Oi48GLitznX+Zgbcnj6CRc2qKy/Ktc7/sXsxD2j
FH2C0Lfr54lB3vdJUIVhOwe61mkcHa9l6/QBxEtxSF7MjSnNJmrXhjvRzlce
pO2uU5vPafrBBRRur00mrg5frWCfex9CcS3gqmKdvlK4pqNLKkhF7XQkw3x4
AojKLQ2JYi4NRAM9iimTzvAElgDfJATof4VtJUR+J4+kID+ypWFzhyvrhp0X
PlfkafZ6Fyy+2JiJduEUCzduoZO4pnx7Cn9m7UU/dV5sE0mwUcBxZ6k0z9/7
0eoVnXIS+Pol3ky/nXk1ySWMoocpHRe6sSsqKz+W6GKBE0H6fnT7khzIN/0t
nRfaKEUrqORK6+OiGkyaQbDqMxqqsv96YG+voTB3Nch441Gk2jnsTc/NjF9e
yFBscBOoEmdovBkvZrk96iqOkzhF3gJf1k4M7VbpEaAQAkgGLEMwphMs4yYP
1R2TzFHFI3su0JPngNUI/1SZnJWrhyWbFOhtqanvYLzehm1aAN0eNDDZS2oO
6JFH2ZIoCVcP8PZ8f+xQZ/OQ1SS6spMjk2bj/1LRYXWerdKuGO3GR8Ks6kHC
pNQor5Lpc8n7rs70VK/4QH96rMWucncwmFvaEBKkP9C+5TO75C1E6XD389zg
b55xfYmM+BnU1qTlHqWMR9DpOXWWaXVgsN510g9gCEIssp35KlYuxFQ4/5mf
87UAX1X2A9csr7KJw/uMLIBwiqjkz38+x2OLebJ9z1gp+H3GqKNA45Ue6xTv
aHTCMOGDxRmJmoGcDnhLMSucOEhBOciU1B3PcxnNlOCtn/VYkYJuOZqt5Ilp
bdjk3GJxlwOJTa0mEjwkLF5aq/+aQTArLGyneWIPXnUo15VgkwrdUg4+r7i1
7CA30XVtwDHMquYWdgaH0bzwp5vb5pvkIDjSx/B2B/ShXttVY4fBxmTPysRp
WnXlRhpoq9hchrEbz4ttPAKcvDy04RFhC9cJZbFgdW1YH9oUzKrvtacDLIZY
h9DAXBZHyLsRHwOMjwKsmsy40rBLXxBRYg0+kVz3oaQ4Xn1AhMSGEN7oBFGL
okXyyIMCGQdoLu8bBZptS78dDrsCAW6rLBEroRsE0y/fAv4Y9ouHp9x5NUQL
aG1UPJkbQ4dKVVbLmcvxqjCACQJ9oKn+AXRi1nFxA8ItqBBXREMPv4vpVzCw
44R3INiLUCdZ/HJmGmOKqjBT3dA9Xvd5fdq72QMBvWIxBHjCUnXYNJUpTRHt
PeJN9w9hhm3VcTihk34E43iMJMB7nt24kKgPE0F/RpHWtEL+k7tHQhc4dMr3
+NqbAmNXmWIXERw60jb0ihcG4MjptyZWPy4qfojWK/D5uVdj2tF4oR7EEMq2
MVomYMwSDll/aDW3FXPoqm5GZu+RrNQN7TK0xTCG4Eo4TeqdqWtChXZMZxER
oNjPk5ctm3ENYauaRGfPMjiZ9ZcV0yAEaWHgh67gwJWEdNydrXV9WmRdLS3I
JhM1akVM+3g/RzT6nKBVol0JfS+ZNg3zogrAjBxGXNtqIJ6lZSBp8wTbqTJ3
RiIFN+hvty97PYVUDnLhcYgzveLxBvUuYG9JK4tsrezIkpCp11HPNF+kZyPL
vYYbMhGD0D/tJfeMNZ8Y8M8+5GnNbVcwerfEMLV5Kbd8HoPVZ1UUQ0hzUnfZ
wXfXYBM0qfE7PkV7yDzHkMpVCEe9DEBlE8aSR492id/yXFkBgDodChXJfnPF
bUF5y3YF+BYoN1LBmKMm18HGNKjHg3SJQXv/3a0gq344X7m3R48wCLY2t8nN
IXE8uqRXVWEwWF4XWznfYF4hSUTtBHPKInnNtHym+kv/zzgXokmUhIZGFvtL
nZnlim62LSMjmLLm9i8u4FX27LBCIVHShznS/NnYRdW3qyyOCJYRlnPPwhHr
+UlUdERuv9OBQwxlgbq9C/jstsf0nSF0unBtvgTLvjKraVh8ZW/hGsOT6SwL
Uw2ASfRBq6hoZATi6aAOxjr75e0Oia2npcS8Pt70BsWvg3b4oESwY+aZTZlx
dqWssQo2Mp21z0C2k/AxRaJCRLE7u+Q0zixDhYvOXO1SQLJhg63br6c57bsy
ZTU0tZn1xkDvSdq0adBLDkjG1/1ZppxOb/d5DeJwbMQITCRAkgIYZP4uYHSt
IpTSJDOKDAxt7WGDI1F/4iQdfnMV2T4L1zz0kYHTamGz4d6mVzGC+YBt+hLi
eYaYkIJ0s3aiWTnZv/uvTjFu4N0iyRFaUFuU9vrisAefQlFbGdhQE3jSKRQJ
fY+Vde0Skq+jIdaIn8eQLx7f+n0YHvHeV+5Z4chRyeezf2Bg3flTVp0GjIkO
EIgPYi8FKxIuFQ7vasJnGqaVQuoC8LUNI/a3AlPARzzw+fhx5cEL1k7vHj7d
Vk/bxkn6zypPS7Hqu42f1Z+DkZJv4bx7VyLp9XBhVKKYZKT7JurgYtqMsq6p
kB2UWNL3CrZxX0w3A4Qa0ANZpPyj7lZHXAegwD87skooh3mJduv5tCOz+HA3
E/Bvlay8rm85PTJotc2OzhoXT/s4Ijoeq/HKsyhnJ8qMbiyoMtLXS1zo57uQ
5JV49K/FNM/wvuyaOu/M7za3XZH7PUrZXSL9wQLuMFxCuzq6dBzC+ht1INb1
vPrHWlDdp6gYnIG6QDU3bThKSVInZ2u0VOBQLygxFmbWQNrGSk/Nc1ijK6Ae
mwb92PGhzvw5TdEhVZeCB2sHehJkwPWZth/dQdN6C+l48lDWYs2WhIvWHxc+
LkomqIxcdeZKR5yYbxaswYwLx4jwOHfPY5kgTJ70jzpAFBqPTUPASvUBBhek
eCIJcat3PDojKqrY1rhcYu3wixLM6dKaMdlCIbyG/lmm+YnsOnakkSrBQstZ
1C2En131m/Hm/3r/riBr7MB67ptrTMepeOUg8R/7LqcFGHvUuGc+FlJvSQHj
P4jPqmE6uxBBk9+RThIh4G42EIuoSy4vJugRFkV2OHsEOS1Aha09MejagVLL
xb9w2z24Iyuy+qt1sFQVnrm7A0EBAp8ije7hgORyqbvH4qb4VkpIo+rWlMpV
STXDPwqd84u+Nxt0bC1HhRE3a9EqRb/CSEQ0m+wGXK/6djXJKDBz1T03TIpZ
RRobcUI8DHxV+++NsRNenDqgzxNlMSfGvRwwDus2y1zSUe7WbkaCiQfabqjT
obB4tHV0C6l+QUn2lxHkauXKVGxR6lNHGVGifZrNq/lY0Rgav7vCD0J97FpA
iK1JeTsSEF97AeuPv6w1O0g14MxlhN2y2xFEiGOgfEb+Gq0IM5ebTrqNwhA1
Ml3wQzz0Yu64ggElyR5/AF50V2iQfGIbXLZYyFY97e+2Kg/H8gugDUNaqDh4
RWfM3bQVqzRZpuDAb3LQZl0Sm0iORaNMp3ozh/tdbBgb7/8dAPgbPsGFHB2y
sDlhtTEvKNNZtHxg94JDOBuEMjdoF4ajeGyebhbNf3PV2qCE6UbCrH335pTI
9EAjI2Hj8iw/P5BzDNwS8CkPOK1AfYik3xrsrX+xadDuVNtEiHe4wdkdW0l3
mlh341k1RHAXMz4JE2Ahxyz/2nIlMsr+HWvhqw59NkbSmo04uVNGDur4KmoB
RMeIBsKNxjNd1bpV90shzEPI0e9f9aGGftXFNVXhGlOtAJvH+eFVhDnwAEc9
PCpAnkX/BGslVc4lqSYQ9Ldiz82e/Tvd1grItZGOhoD33ez9Jqa3AI47ctjn
+8IRgsBKg5airDybU4OS7+TSE8QiQxU4HLTqqJyp11nSR6Znss5XxiyDa9vU
SimFeIuXeFjde0IDPRgHe0QFzPW+PIiJn+3wjOIpbwMoSOUPThTarr5P35IO
cAH8Yp8mrzknSGdvNs1pN5ZuCbDzHtSHQsWRny9daRTwJFTiHosiA295gPwM
7BbGJB/0CaxNfRxNcLvs4trG/2ncIWapmkwROmhRF8kIlSeTKpMM3paWoMXq
AFVoHdJX0fqJ7c8ZRQ7OEvVo/nnovLm4oM/y7A8N52/AUU/uqxhXK40F7Fc5
z9awWLW3hJkbyUC+rg9keKbDF6t+/R90OySn2N6NRToPWrus2x8oDuzPBMHv
Chf2WxIujzGBb/a2QDpUt8NgCBgzwc+Ri9wTq432sRndZjKYcHf6dvRtQIxx
KmqQ/zo/zjzWzuBqjqGL27XS9/P0gS1QT4jlfSSMtCaAY3BmdSdNtEAO78/g
rijD8+61myUwg2SUrdVnjtaqeTzc5aL4hznKQ//KED52Yl7ktR3SSEhyTcJy
Emo4OlC7q7VJsgLUV+O9pIiXsnroPdxOUhewm2aZzISDgi9MeV/8AfcigwEO
ERk8H+GiY3BEkF7t7WFprdZI08hYy8bE4WE09O83tWMgw2yz2bkXSbXhxHxr
5Mqnup7m17cu+4TWRekJIktHJR5At4rB2DJn+nLnm4Y1EySEaChiyIoREgo9
LOhNim18PmE4zcQ+NsxRirp+UAY+05fzIBC+f4rcyp4hAIuAQW5B6ZShb6F3
pYcmTF+f//Gkcr+lU9xMwMYfehn9AtJAbUFCsWEYi/TA7ehWB2GVMwuY0MG2
B0511lEDFmoI+MBiBp36yTY9UHVBx5cBFwxFPmf8axa12PhdMAJbSlIlLzdJ
R8Yoj8wTzC8f+/20hJVH4kmqbTLe4Yhh4NcHEwFyQ1KrIP93nEsadlhPEhkC
NblTA4+uUtsf63xPqnPRdsoTzL35DQXc9QK3ybgdbfuOI4LD6Ao+tQh5Zw48
FvZc6/p9Bqn7qlklkOfKNVXKFkN/jjOABLSp+gfoN6YP2lYtGa6FbKiLJTRo
TaZcoUsO9sfjYddTubHwzIutdG1mCEO0OlmUXXZzzxzamnkmKT5jdDtXJ4Ph
VVKor/c68iscfxq/ScZGeFqfuNMezQu51sPdCa0xX6DMzY8XRZgyW2lrPWEI
MCZC8wcgzproghsHnrOXl52ygb9NX0vvsM7cxLMOVxFafwPWkQb7gK+jxyIa
M3BjtiDmxUJElNn5RemdTTkKsdYRbMUyGVhXQ4iUOeRpzEQg0Mw1lieJwU0d
vF4qOD3+zgPyLhSPnHqpuApzru8BobF0VekdtHDyUMKh6K7PD305r99ynF3I
nSyQoCcUmmzX8dKaASrcBmDvj+fktIFffKPvD3Us41TILWRQUYVqDyP447pF
oCWY5ULQ05JphdvVpqsrPNJP02+gwSF2jjtoGMTPpWHzNHmYDYRFCJFcMacs
4vl1g8t2eEn4WIflBwfOruN/A6u2mZylRCPr18qa73yIjGRhZ+/E4UQ4KrEs
Z/8JdS/XQbSF6YO3+AcRNAc+uOI5uO0y/t/9LGxVZhcAOGNosQxrsJUT1f8d
HI9PFaNlbvIVe70Bs6e0XlKyb0fPLcvLL8lt+gBvxiOJwNOx4wo6mwaPx8pK
g95I6cywk97Xvk3ObPnHf6EIIkiC0JjuRh2DHYQFaG7vayn+oC36jKNYCaCG
biTpFrNqniUMV4Bb/5Vjq5t9xHMaGKnplU1nTxiIrYn6ndfAVTR+o8weTSHC
sf7P5u6Lx2BRh840AiTvPQH+RaJ9wRbC2n6cRw//SWThgpvs6NwVTnjA6kXo
7x4KI8jTcgwcf3ZJ+k3izZ3plKC4zVHKX4lxsICH/OW9xQ8tKS0Aw/1sRdVN
ThIc4dI9a/2vfSKIPrTvy9EixsmhqkQEn5qReahcK/0BXcJ4PN90TnMNd4JM
LpCt7K6Kxph/FhT8Ssfr5Cz8WlCDgXOoz0dc3y2UDhMKXZgQsBNQ8FMwXUVK
8RnFtb8nT+baQehHdzV9c9bvcMMwK5tQs1SgCOoZ0SBCysMvqI/0l/oITa2m
BVO3JKkULz8bD+OVfjO8bDUsdD83KlhrO/lJueLB4UJoyRXUL5i/6KLN6ApQ
C5NmUEFwhLVbhp2em3uO/bURONSrnD6Ei3KFE4Eviw9LsvxF0jfJclF8g8eR
uVOcUaA0nGk4R7H0Hr/rzkC/8SATB/3kNxeFr2bbp8wJ24wi2l+q/hnzU2T0
Z+6aYq/QWYQCc9egfdseILrCPtCI1KxwZn3IgWVDYJopYGlNsZIQlHkSXZLr
t/gZsYBcqgsaDgKBRgHGGMKaZ+zyRkM0/ltXrL7CUkFyPSQR+QIrpYDOKpwy
41Z75xtlIdKQTcrJYwzUUAQLI2qJzucrNqovuZrdl1Fcd0BvFR5CQBtG68oG
hIS3m7xCQQoI/sMaUCb3t3EG3yEOtDxlEEYiDERvuRb096IWx/Cb46diXbNz
WUYzJJvqSNTsNBKoQSCa5N7gDkaCjhxNP/LEaoss0TONQi3aktUU2u0e6sve
N2cC5DNqwed/jMC0l1V9OP5k00fJ3MOpbRW5eCY0NSSWwDqmCKEoTAV2Y73e
RZ1YG/qcc5+IN7he/Y7UQo6lDYCedPg2kXaiwrsQO/6j9r38/BYmRq1bwGu9
IxnkIpwpCsHvyagyR5WgFBpHLL+iGS21vPORX0alkdHD5avaX8eQyl/yMzCr
C5VpQgA6KAVRTwY1etmOfnLQSf7EyVqogItZJLvhkV/vGeHSkRrB2PUAg8uP
p5t0Za5yynkNhDZGgjcG3uN5sdlz7MAHvFTUjGFjljo/I8ZTFMcj/RFPlLK7
sGEAmrYMB7uy9DcOn5dedrdVUNNcO8/1eYcE8YCIcXDJ2yVHBG6Akk683RDf
Gzp/LYmEluHPkSokwo6uJk9GGtlhPbT08QzASzCTUKO7rXjlVYyilNMugSh+
nJiXULAf13Tfv1xxFs6hTKtkJYZBwqyc8YNHfojZh7wjRic2gh44YkxnngJI
btjqz+HfnLqaq3DcG8xfRrUd7GVLiZhZaO1qKABj2z4En9jswGlmf/sBhCUp
1ukHWgQZJ40uXyIbu/lsq6zw3F0KTl1hKt06+ucrLOZaCqYQ8AQAybbA7emR
WlC7TBMQbjeksF6IiHM34+HOutR3s6P9IVU7YAnsclatKY/cZISw1EbKVGyS
aNnVZ1FAOfkO0p6bplbAtmDtYJKKvm24hAQKWEmieiEAmyE5XJM/MCFfUQeF
LK1VjZUf4iRI5oaARmHpcwv4pjaWH/vAGneS37A7DM0J/WAgI7nD6hH6FhIx
CH9D6XAGnj4a5KpSRRy3N/Xn4mjMuE5w2txBmDobLWGIqNrL/lQQD5QWLUwp
oRnyW0tvYgr8MIP1a2NTmP6kPp/ELE3xhiOEeRwEbghFit1KE4yCCKeKq6Vg
BKwQSIlqz0SFW+pn+C8Jy3qfIDlI0WONWXOyElqvK1kNlK8NsW+jRQBaejJ6
OfFpwXm2xfoyIIvWshfy6XuDKfWvU0/y15k+1Vh559hAUuTRDPNffU28L8K5
tNp1SyY63bQ05zCC1i/7xfrBM2/CA65KEO6hlxoZJwu6qiAf+9Irg8f3u6n1
Mbx5nhjwqtMlmhSoMROC/3f2UXQRNkPAjrqH/35hLlMa3Q+ZUVTdr9vgevB6
g2wZOxddn8MKa8hNW9J3IAX4sZuUNLuEGd8+WgRvNHlQBkvmoOO3WXmlmeFj
Ets8rFOYGVhzLphpox68DuFbIo5Es1Ue/fD5k+PpD0p/Arw+2cvTZb6G2rAI
ZHo4Mfvoanotvo5JZENv/bVYpUjg7Og/yjAwdS4nWn6KWbt9kzId3wbXfH+S
iU4VM+z16wGPCc4czx77neeh5mOCGyILqmEBQj/moM7vymfV9Kl/X6PjLV+T
cLxl4DTp9c6Q5OI6Tc5CZqIoeU0Rlp0M5I4QFcJRzkPth+s6rMmnYZL/0fZ0
T/9KlHv68lnl07wMU/I/25kfyuKy+Gil21z8yFR4p+Bo3+vWzSB1iVu1JFJ7
s2Wn2I6cICmooV/nRL/O5hD3EmdhnuRUGH0ZHKkQDVy9Cf8oNGDdEDNbXo5p
69RaDVa6HZ7/9Vq8ivUOpNPgLO0o9ll744gLpYmuPbpVyNesx5kgqtDOrsTh
0/RcwAFNLVcO+nNLYeLrXrRyARpyQoRBxTK8zHeN1ZHtHSM7N8CNYKYdCzqI
OpuMzPQnKGWmRwBmG/H+uxxdXmFtOoSH2jxL0SHJHagnUmBbR/GdbcDSQvSA
b/LdTA0Fdlj2ys9G9EWVMPXESvSl48F7q6f44jUBobay9Z2LdVukiVCREZvr
pDh3sunkd+GHzMwsdTAK+67QvDNDRu0nr1SkcyA9LvLp2yOwav8dABd8Pi+F
IZzp0R4ksMXytT+AuFVhG3qswujnu8FteR/F6fCEUNAiAIhHME4jJFhqHnfy
Yp2g2b4cWLuHG0pQ0rZASjJxqpU324LCJfp2VCEKscvZbNRrr/qn7+qKv4IC
jCAsAzLI/EZNTLyDN+FFZHNDIJdVbek4yM6tvRCzUBtQkU20q/X60hjwTrCJ
s4cPVzVeQLWKyc43XsXLFc0TcgwbvsAqF7Dxrib+vBd0hsbHonMzi2QgowMR
uB1UJjaQNjVnyIax7eZn5Vy9VSDPIvSOTgnwn6KNguPi0RhKZuVeB+JWvOTD
qRpOZHOk7BTRGqRN2sMP00d2tHkf54Si3sJtwBf6RyjOQuq8f0rcJpjSopsn
GUS7rv137esFF673ONi47E7Erb3Iv5kgAF++0NycKwDb6heSHUlAcnV1fqyu
FWRQs2Lr1mFLMSLDkKJ/95t/HaPYKXOwqQ18SBSwOXU0HqEn8Vh68/N7/LBE
QTEIcVLrQjfCyJwKRr9wgYkymPa1qS4f2gdggXLVw+3AF51J0s48YUFkQWZn
sSjdBd7/EEtp60PrMMUz5q6Dd04ZcolvUPII+xVCO5OXZ9r6/4h6U6TWdzow
MAyDA8ezjcb0Sq5u539lPUB+EEMFpG6r8dC8+vuloRQ3AJt6dzkFJMfsQPPr
Ovoz9wvFOVnUeoDYnD/gfEK2mva1DSJp810W+ihzs4PKOvHInf6/ivba5S1e
i1rkavOXi3ilcAKhPwgs/47figPju7ZtUv9AnT4qYzmGIf32v2hx4odngcqQ
KVu/lHl+XH7g1Q/by3qxNpQyiu9rDnspBhbfxuW56Jcn/x08jXbSHOlO9mfm
Dt0Mg+ZGs4xi5r7tn0dSnJ6Mhp+gzMk5gx9/RPJoY0tOhKLgJbrhm0J8/crG
mP9EJnMdrJ4tdl9lPZ47L1gRweYKr06T2tX1WX9hUspn5zxyFhViFHNmvPju
FAMr+g9G/5EbcGbGc/STOUlTT4hIFu+CXmnvQKp1t6SxusGiecD5x85w61Z6
2ceO306Ge8hs780su9pmW8p/jSJBkMtoIpT5dQFEf3Q4T7MPpTouqJP4w5k9
WVa6Ly5kcSQA3JC5J5gbansN7/EtSEPo0adFe5+PgL6DDeNu/j1lngFa/PQ1
ZC9sILNalTHrJvaX2MiwJ7/BNjp4Dhj0vy4bM+XQV7hY066erxXrMOIy0kmQ
dtn1HUgWrR/JvqPuiBtpakXSmXzt3rjbms6Fqj6liIVCaWUlX7qP8TN+9bwY
d0ueqOO3mzmfCygVsPUd5xWP31PfdRKq+lQuc2qjzTs09fy5WJlMyoup95Db
fjnXcDK4tslwKKCzp0GeA7jGVqdTjhn7hURNu9pz52hm1KSA2NLv7+ZvhuLd
THgVZbCSJ740/G1dthJF1VEAIoUOnaUIC5UTkkOXjBH2YFQ5IBGkyb8A/uY4
SZ6xOMQDXwCX/8ZzlvD1T1WE8UAkBPEjA1+zdlUi+SLq+v1yrApK5bjAEovl
a1xsWm2MlR/pHvFGgcAJK5UjSH96OhQkJXuFfD4M5FS/5GVqWIMvoJPTxQ4+
qnnVVjxkkRHGeDoCm1A4aJvFozujwXS9mvVcPzdACXte2fKHjfSNDV+oDCIs
4XLReC/xSwQVBMXwxstUmYIx/906z+Vae6uZVQBm3Tqp9IdVnhGw67e99tSG
zxWlhmWSDQpxjBmRNv7B/K2GtogsBc+S+aFKXGtGUCx4gDbZPdVMK3QSSbeN
Bf/wLZ/BTgrLxp/UwwB1cfqmaBU96IZDQ61SnapU2EsK+oIJS3Hj5anaTrKR
4Jlwh4pourvgqaVD4nuYJ5Z0kDRUk6yjW8hjEjN131f+Nw0jxpplyKKrWWFv
56rU8dapfwbCsoTCIiBHxmVDbSW7I/1YfCVKvZp/ExTOzPdUt3NuSX/TR36Y
u2IGwfjkdzUTGosM3odw62ekgKpZ8PAxAfYFLlGje/F/2Ch2Hx5c9Kt3vrxQ
SDv/0iSqqZVSZAy9kB8IYPut2tWDivQD2WypI7jiYvhlh8SUAC2gqhqcO+VJ
OVUUTsnXl4B955wCg1Tpc0gzLqzR5gMkMv56ZBeEFjVajdCn9R9zGMpHAudb
nxGIIrH41PI8aCNdU2nEPGQ4wWTra5Deb45+GISutg0mcB84eKYGMNomUfCD
52EjH3YJ2546cRWnakjsY+lruBJ9A0UccoCqTC4qrhSlaDG+jkabkX0Lxfoe
0szY92Nk4sLXEirlih9Y+1b8O4IZom7zDpiwT2JLrUzbaKNz1v9R6eWtu5Mb
KBWO3BWEiPm3hq+koJxzDvajJrmRLlsXip/Eag+w54Mo0UiSYdhsHhr7pnvY
n7xH2FHS0EMWDiosVaTB94OUIuTakNWGIp6UMOf79AIgYauuoWl3CObKr5uJ
piiyEE4Ii3p+k/GmLDuSMZ3H4WGGLNH63YHfxv3jKHiADojKkZI+Y7bctkrq
rT3JYCB+FH3WWUOQrZeF2N3BgtvHTqBqi+dRZDLHVP3HwPAwbuFH5P+KYRf2
Hp75iUz4hEsWE0eoQMrMv9bCKAJCv7SY5fEpucrCJODh/Diby5gGr4OqmRij
JqWvR8m5860uCCNPAId6d1+/A0fJY6cSJBV7xaSNPBP4uKspiEUM6hPDV7Y1
rLtF6mqDXzm6Mo1QIYqRybRm7ygTE22cVNBzKXGjMbJgU9woB291x+A1Kf/X
C8ttgrmIEBD4Y0biGmlCUexhhEbjSHgD8Jp39EwmpfDxLMXfJTg+u2ug39qK
JqYppduBMtJaWoD6jNBP6RhlFe1IRMbsAVJ2T7eAh+3Wf8GEd97IBbMLWTfP
fIyqgjpJeCNVTF8H9QairjKLEAHSNmlCVIJ2nYBReG/sXaxIapliFqOFWhG/
pjQ7jw4NjGL3QW2lpqVTSffOsPDItlxiMRxoqeU8uoq68RDF4eCM9G6f8he/
NXcn5GgnmETO5uw7xpTyqauRKAfC9/7e+tdpAqi65CzC1gNsd4Uy10TAlpm8
bpzGS1yvDI45aR+68HekpDfsS76XjJoqq5tqJ64QsMi4+vY5OLS8957stMfy
y0xLaPETZYB3lvVwuYCNXVfBzYbDWjxwETGF5ntuLC1znA8UVi3lbS1AZSeZ
HCwHrT9zYOqc/zF7bS9hZth8jMVbactwNjWFPikEKTRr4iz+Fz+GNGKrpWRd
X+JGCpa6K14mCI3h/TcrjRoKlkoUgt7rQNCjcUGQfGd/uR3QEqueM2IWvJUF
QGPVKt/kyURI8XqjJ+ptHcwCOtWBGrBFfGnAegCL93nP1C3ps32FAFjYgd3K
7jamAVMMkdop3a1wiQkXXXTMbOymizN7zbvU7yMBwIwErOW1LtVFndbvRi16
x7KKdrsj0L41mwMogW230X2ZzStNQGS3N3SSXGEJDREhCaFBYhWneLD1jUGV
Uvzfi1/pofuKrwHTwKXfiMOSH7wEMBMM6Lfh4j+fur+1fSQsbRVnPSKoP13t
RpnlqG8TzMgWzjK87KR/YzT+J73xEILeHNx607ImsG52Z08A3gpJCHgeJvYX
aDeTvRgTtFkzDwlyzylMNRRcre2ftJmD46wMRJzWyrhuk6i5x2xvBn7OQMBz
T/MEjfcXDISrk6epBKt1LMGBaMUR80fO4SSVPeKfgxmYvXDRSpHb8SB0OmFg
+BPYj3R4wmKXvc2Fm5jybakv0En/zuVyGoY8f4pt+mJuBUsZOEPURJCAnH0Y
hTT8KhtHwUb5HPLek0CrN2Q2aWRJicFGG0F10FPayJHtoozmKrwQGR0JCqih
Umy4YgstZ0hH7/EsPv7mpngqsMC+5VnzYC/OemAf/xC4wu7JTdBiC+8OWx7R
LhCGC3G7TV56vGxW1i3797FhxAegwZX6stjiWNJcK+LhBu6nklK5zkTsPJfm
OXEu/Sfk/0lrjCHPtV4DewjyP2wnK2sQyGqKYpXyviDx1cKuwQKTjkG+3Zxe
x6zfZvuLW/61SWVpgKSnlSeK8YHW20x9RkqVaj/A8Ng3/WW716i8+2Z7xd6n
Uk/Hy2/2CqG6HjFih2PvcmgvgcDuaHfR0kgs596o12Js/3z2hek4HcJYjxtK
e61My8PqlhKVDFDWys2J45aFzVq/DYEH7pOCG59SfNRq6SYsxwisWXmyu9yZ
OCCB53nZPYZbJaApiSL2paowtW/JiQZI0YKNwCTDLv5XMowEVejJL8OKVog3
xeVQmdycCCS4hTaYB2SjHoCEJDM3lh7iz/gNYtQ6+zzrhBoGTcOPK2fIVJoR
Ad2teoUwYvciHoMXGXtDRIWrUttNW2ac7QtuFnpXJhQIisJQ6KBgd7o1b88C
zHWjYdufvIfwPVCT25Yp3I+lLqJBo8MAxz6rjws6m/l93ZoGJWXCEGzN5Npr
DVPsEdn6voaegyD6NRi7Qwj9E3QBtzouXMsryNgkIjmoePSAbMThQIN7jeYr
eDJuvyPqvsL+3c/WVa6AoEv3l1QlAf19VdzeQEngDOnMttvTCvESJtwXprMw
NK44XMzyDEgv0B1sl4XKos1LKpM6YBYN3rEVssomT08B/CZy2to8ZMXRJxEq
uTRpz2IK1+11UcIgcPrwF+Y8M/IsK74hrFMaYPmwttYy84uz74CwIQjgN+3X
Fnrdo4cCvJNLg8f/WXCWb1GuF1vNU20ojhCeLGDMWIonbjRd2V3ZmcE+oiEn
R0KxrytwSofiM8+WIWM6CKBu1bXOV55/fURmQcT8Q2TSv2apLDxtr5IM0Ke9
lyjjjP5yoYoeJS6AzXLN29FoFLY9QCbuYVshEAwwxwnAqTHwr2Hsu4mllB0F
5v2yyGZNJPnnFdFOKRrlg891hE65vSlV47uGAHtfrejUkM9Uto34FCSb9N+l
2HhnZFnlC8acQoy79aDtpcrWuKmODeFWBDUTjmNUG2bdHSNtZmojJ0hW8bbm
CxIoIcKnxPUtdx+u27HzS5jfnFCp7/EmxtmAJTDTvUYr2Oryd+xJYfoFLWSc
Y4+5bJeEeH5vXDjIIXBgFoXwohYOCYtj0Kc1JdH1S8fIx6pVsNyLcl6edcV5
DC/zDJxznuVTZTOm013bBWXp4qh8vj0wRUpqJH0LtivDq0/Axw8n9VPnlujA
T0XemYB3pvulbLnQ3cEwq9NmF1S8DYDSY4u3ekq+LZvkBNnBXx9P3ZSC3Wqj
EXK9JFFppWNzt7X/IPwmHeNW+liByA1AECHSVLnr6TPuCtgXO+YwMH854bl6
Sm6Pl20ygbvwBcR9zvGuF6yrj4KwEaxkxLo56W+sMzncD5VusnVmxzZG3XcL
SSszWmCV5LhuPbrleasRI1b71n3u9NJFZTSue4AoeYBdN1GNot9qg7cqMPDW
HHryyv19SQvJ5eS72l/L1dwRZGf9bvHZnmzKYdKsiMJSH6Tk2zi6N2T7W2PM
pmSvggWlaCBejlH73Gm5hF4AX5C4CWA66LbjlfJesgLr0j6NjuzZghs+iUTd
5qeZfMxCNve33NhpXcdFgqSBqTX+qug1loAt+V9MAIBiwZN5EQVr5zUm+pSI
osv4PV3izgdLauhwYN8tDmMhLDRC/Wg7hd86jarz2KrYPyml7IpIFmNWoUQg
nFX1c9732OINBONfidHLesOtoYKjfT+Cfe7uQrsheOyM40L3RneQA8k4Xw1n
sYQc4mIm7w/veo9OZ67Zviwgkk1qXbD4PpzAbl6lNgN3g5TsvPQ3NcEriGQ+
CfPBEuleuEr06m8iqtbBjSzNkfShNWY6kfFJ/Ty5IuPRxFZOh3OxFLit1hkp
OAdG+RwicaxCUbYQTW21r/60cRR9O9hooxamP+xYuXyIqnIgMe0sbovoAFWt
PyiiI62ptxHcCffqNMUBWPl4mIoie/iBFVr9vQZqQzCUHS0ysJNNJANkZ9g+
Vjzv/Ze5vIM9RAoskasa3PPbFAtpJNo++35TQy0AV10ap4NNDXMrMjhm4UHo
vqEDm8ch6YLDRgnstDBrF0v5YeQXk/I3b50nOMqrsIhhgSx/CBLsb9rZgrwB
5540QE+aaCb7JcLfW1xZTheVzjlME76uaCD7XoYlC1e5VomWOIQwI5iCrVEB
hvr+axeN27K7X6H4A8X0piPqDxGjwfNfv6bZ1fgAioUMh1nQH4A4w8N8Plzx
IszqyVpomhk9HqXaRmjduBfs01TjSmR2usM4AZbJ61ykWzjtWEws5tYUL+36
4wyzhHHN4jbd44ZYNCpJOoyPpwd437OpS6kVI52yfbEnIl+20jcvURzALJE5
twSuHq3LA5sx1BB1ppykK/nFKPiZve2ojfY6UPGzFE/8/jV8xPv+dgWrKb1D
chMNqdNM9DjmIAsvCuKLUzNzz/iwhpnTN9Mdx1auM1n67e1pAtrfkjv2FMbw
+bh1RuMkzhHr8CEMkEUeMmX68S2GEPuGj0LD/RExMDMQg66lsThHzXODt+BB
wdEwOciEKbDKTen2GgyDHs48P/cgoiBPCzGIo8TH1L8DNSjKMeWf/vMikEn6
dUvr3o2k8/enRRFJPGvQL7RNy/4mIlr8t0RJco/Sb1zgX8xHYgsMBzjMqNsk
MvhHt5sHDQqi/mkVZFh8q/6OjGUoG0n+UO5iFGwyI6G4/zLYgOk8BbOZ1kw3
1jhNq+ZDTTI5SF2cYjwzb83hiduZP9nUTpGAKcJe3c7f47/9qfDJGoCZ9PUB
7k7HoXOTL5YnRCFPDOdKa/5wXaBkR8mcFyLjAVBSvLqdsd7awniuGIm4m9Sj
8v4D9spfjxLQQZO/TQFablu1OndtSO+3ZfUCjNOCLa5bNNYDujgNwyyUr2eQ
BgD/3OWRF0oTbTu9SHzUk7IorM7jJjxTU7yT0fc+X4Ybp+1XPf2hZnS+vCkN
5RCE2psN1Glthae9qZoo6cKYJs61e6BaCHn9Xh0lwqSUGDh+i2PMlZycfzuW
tTurbHbjzr/bMZsrrlSKTizYY9S03bJ8D7ub5spWI7iH6fSFz3y/CgJBHcAn
D7ppL4S6rLjpvl955Fc2SDJG5A8YVaSN+/5KqNkB9eQaySqLPsTr0I+dLkZI
Ngo/TCvWg3DNdckHyJkrCtRUTuLyRygvKI3eQVAKVIdAIHNmsIhzPUyhI1L9
1zQtxGp/d9oVlucjsIrd8wIhzcOvsKZCx+/mTgqUK8KX4VLGgX9PMZoSio2B
fXVG53TzFUg/SKUtsjeENrD5OkoueUvgCGkncfTLATmGRTDOnaiFooSW18X+
wV45s3CKigZzXI6Zwm2CviJgSyN+mMK3zgpXTFwvcFBjHack+Fs0Rk/SIunp
LSO3wpU5l7GGfvOtsZ4GPK0EtuuWGyqrPVECuKebhdI2TMyk9ONk7XZ4XA7X
X0XqGqbn8WsNPWFTlqBtmXz4jTFS4U/uEfoZv3nVfRAwZ8OJfmEJMuwCSrRs
VFxfTFFciHJizcDNB3gUtWDNVf7EQNrn+geXpN68PgWmCgXrfu+9P3ufjRng
/JSTnYPFuN/k0CCHDNr0vtyIwKlTvY2//CS+MoWDWNjFz23YZtdB2paZoDnJ
Jlvz0ihx2/5enW4Zexex/BhZ3r/qDBPQaIx2vD92J+8P05mDCcMXDJAhihks
Kqm+cyUELZTMlvr6behhCcp+TZuG2P9DREIdZRMtSZFNKfakVi/KjhWVVOLi
E2s5rvImJAnQOhtmej3aS0SSPg8xmrjyU9DysLMYka7wwJDS6d1dWXEaPMJb
cIiKhTajsch0SUnHWC+aYGNWFT0/+F3kJ1EXrlDwercZjnF14YwObyVqbMzF
UFsJK1FNLsvuIREE1o7ELyT8A2LBGWWVC7o6y7LbU4opxIeypFihmbuqR66n
K4J7CBwEICnZ9JkDdY+bGxIDc7zOhAWZwLBepOh4is7vhu7kgcZlZdy+XbqI
F9IAJrFYK7jHfhtVisEnq4qXxoQAiDaxPyTYOVTFWSx5ymo0X0lr9fljD5Sh
ffeLyBm5IrzHqjYObNLM0TCRdEChEsSQoJLZK6BcBRCmwtVLbw1czLz/vB1c
qW6Q1crOIZvTC8jYEZkLCstSmGoaNjdxasfY1lrNhfjkg60j+qw/u5Zvgcak
1k/KTYvPc5dv9mHDZJW2G2tQ7k4ctwiDWfmiNn3cN1NsK2lcMcYiZ8JTx/Fr
DGgl39xsu8NX6x4T1mJbfFqYMDLrgKy3Yf5uMKAi+n4JypOzn5eJvyWohwXJ
BIJkDzRwQNq5nQ1KZW8UtejLZZfHgLzNlAFyfIjnRo6Zu1ff7uqiAjW4cFeG
+JhZTim4EQ0Tjvp6MKRK7WeWBlFXXc64aP+0/pucJv41mlPluRKKFYyYGydz
TZ9PVZhH8/OADU6/l1ZBLm2QBSYN8RYJ+xa48iS7K5FGZQvfHZdOz3IQ2E0P
2ZoIeRXuhAQM3+WeJpSKemph8Xc0EOTAPX7UyQrx8K/WB3of31zU7Gv/7w+P
FVIT2Yz5l9qKhimCuuKvndu/OdGR+dYbbno84pf0cMoOSPBwEwiTSGAVTskF
680SUwjvfgt1eYURSLUxRBeTCK2A6N3CqB3V021EKXT87qXHK1PLIo6I+U8z
wo5JDhKNBhkTwG97VJfZ5WRu+jV2N3DG5OXteZ0aSSUb7t2qo0E1G2Ng1+VE
batmOq9k4DN3q/fIDP2RFObguQm48MAT9N8uZvHv/BPUir9KPHdZs43CGGcq
E7xPBvEKi6Y5kHORqGDs5ysgwwxwwt7kImKC7r+wcUFYAkVa8pBFdF3BHsIE
KjQEe0PIWlH1OA71dQICUwbCB1DEA6CkkEAxj2WI4ByjAVYC8/g8Y8y0aTel
ESy31sk4+j2cVtxZXSpBlrrYUcKO07RwM7YlAn7ZH1835jJer/KmM5aX72yo
Qs2RIdkaGpIHMNVbctQ0rN1NC02XiYq8I7GzZg+8jwae8fgM0LR7D7k2zlfH
21/sCSv8K9CPeevb4MWIcowUKCDUdjiCWbRJwjy5xIiLX7bznbS+Jiy+Jp0O
WbOkkOVfoLHBNEqZO2DWREAxF6vSqj3kOfjQ4jhJLNx2Qff9F8VZB+nYlhmz
cS7MgaHugFmD5HEgM1ltU/UENCq8BadebToT/BVM1aHRGUp20Nzeq0Sk/fG6
ZKiUpFSDpmtvpj0i5kQPfagvCkeKsI/4ITtQt5loMDhkXyW1nB09ZnMR1jjl
TDOf/dsCOaQG8a41qUa4jJow+NGTYL0izwHCmJjoV5da0oq8o3/n0dwq7Dis
hjzZrO7gQsjavRNA23FdpImcvS4xJFPWy091apywGeqTshIu5eJX3a9PgEKE
ztkxBKjaD6TMDS63cyr873JEZ8RTueT/KE+bJ+0Y4ziJnQGG3Al18zw1TUEG
en7w2VLNa9dfX2rGlA38jTtFXzDX6HipBxU0UJbKhfumtu7KYPIPTMTtMrEm
J/H2ugvhRWfIlvbIcy+1AMrF3L3ptKqqXhjO/TFzB0TZa9mGwhOKqKmcxTYF
HZxwdLocKp0jyhRPfy7LcXAQtDuL9R9/L/Sca/uZQ7/9Wf7jeBSJRYrRGjDs
oDcN1G19pzZt/tBmY4nstwmjNcc4lPE3Ud2z5S/hGMyMSf4JSKSni1ZG+hnj
5MmuggtpsLUFjp5fPXOVuqzjY8mX0eJfFm0u3NNQ4yg65ofoDEwg22yxORyF
1MsoPv9c4ZbUQocn55S+Cfs5De7TWlRkw194py58HzCtT0GGPiQ/2R4LoWqg
VCsPDKFKhUncfRmLQNQAHcmAiRUlriUDeNPMjxUWcE8ShnzD3qCPWkIMCU+R
BWDZiPBE/mATFC/bX3dzeI+S9fsSwePA4JeDwsFWuYZPoy6Kg5Bl+IGxTv9n
JQ5i/c8hdMMhnUnFFW8z1bxj4oQN51Zr2zNo691gC4QMfg5KnzNsW0NEJxc6
oL5dx6t8uJSdByUNMTls0PZ4fykpuj5k6w58if6SNyG01fVu3SdG4aJYvQmQ
xRaCcyrzw876eKzCJAaLDbzjDeqJIDAKlsSooqOcCyhkkAA1b1Bbg+PjCVYN
V3MF786XCkJSO1I3OlGkt3JCqwb0q9MvrIFCdqrJuGaOoZtk9i9sYbJ0Zu4k
RT17mmhCSUCXw93RZX0l8H7AM0xvGxExYni5+e1YLS5OW90Fp4+rjuo9a7G7
vCMBczxcRME9010GhlnLlTRYVQ9a24imlqOgjNej3SvibdVFNN/hfUQTRZ5g
saeMzBuSsT9REg5cbkQAvsVPW9TLklCqXjSrBLQD0zlsLmZ6qufUqjJixFny
pBIQxVBH7qTiEkpMuCgTrH/09Hzw4ycBMo7VTXpOzgdIxZlfd0N9eMm8qirZ
vEnpiJ9WGUvj1KoRHJilTS731mrHBwt6onP8Gm28BlvS+7fcnBbyFVZnn0dY
3sCjKKTeilEm0qIRYEiQDtOg78kNC5RDNy+JSLpGr7Ye4KBI93E6BrS+uSah
ujlQXNYI0LHaZjuzJxN7+YQksODlD5aVbDqB+9KZPDAwnG/PmUyhUijwzjM5
omVoXMqDm3tDGv7r3m0X1UlqnoxymjZAiVmwPx32ZNwwE9wIeW3MDv2C9cTq
ARcQopAWbN0IBIY+z4vKIofTrRKlSkqAr7FLV5bSG2DkRfvn+B6olcho7zX7
MT7UczBklOFWYTZoXE63LORr4JgvgaHeZa12kdGjeTBTzp34DAhc4RqwDI7x
+NHBYsr2Pcz0PjCU3nVdLqKN2sCsOxrMCleyMYEQ1UKF5Wj54zr4NQ2+F628
ExL1D/Jd0mcs0/b/OuEmkmiyexo3Wc1D8BKcl4BSo43qd0PrTfkNYUuJUjjQ
iHVbl56mT5FXLmaQNiEM7giJ/QrlZcHr8hylqODIDI48eyABs7aXd8+54jrp
DX3+3fpCdvaa2ZL5HUPocpfMOyZaYMkvIw5gPu1CGHvC2eYoObEHVb1fwDnb
2DZQOMTpUaY9ARdyBq2pSDk3gE+yu3i94WFGg9vecHN/9QNa5CsuVQp1ZcB+
3xRItytbdRpAHYmdc0e6ynKc+jJ8QeFstYBMkfhmB+O1kDbAwG+19HqyRLKt
0JIP4IEJcpLR3cnCO10oLTtwfTUvcA+Cq+RxM8+nKFlz0rr6XQSCTDZ3nZlT
w1hBx0ukVq3S9i5jTtHXQUUcklKO0+zQXwEACv+fFDFwPZ6/vf3ru4MkHfPH
RPYyJBwdgIld8w7YWEUxoXfA9qDoGAcXuY8YWLhDQ71nPGxaC8Dfz/Zwz2UB
ERKDmrFS8RZGXVsMWlxAIuiQ/JBerqu+RAaDcleOe6a5x+JjA2fT980xMzOV
SeNG64VdikyZPIkzEYAN2ZjBu1azpemnk8jGmOa7OcRM6HMBWwTyb86Zhlef
+ICxUw0A1i7RuuHIAjydjMYcGCxhyiqyRXb+TpRk2BG+uLjQoLDPh/4z6v9X
FEeZxMfjrMWT5jNAQDO9vm1TpqDCtwn0NBvlOayMiTuA5FVehHhD/MYr5WAf
Vd2QwMewqRx2Ju3Yuqu9bI6AyNW1sJrKJxfNAGfVMlcoGBRSAFAm0Z1vtk3L
vzSTVWCTm2ML5CEK91OvyRDF2qRSY7arwm77zg7iu+WlRwkDYldLty7ThCwX
fjguASbSxP/TjSjxnALzB6lSwlRXOtmQ7DaIQvp0OXdjEkNmGSXM+4NdX/wG
q1XL4SM1eY3jFWjnQWxYF9ag9c4T24QJZxw1I5a16oEl0vw0k6EaueXT6Bal
rW0kDR9gbTUJMhFrGMCDE1A1E7kNQn060iVFnwAYJIC9ZzulCBSmhnKCrTw/
YLHdCzzWoc6LKoHUFw+7GIrRgQCeNAmJn6PGBqEEEnMz/nPykiXYW7JXpCYt
acNVGfmjA2JVtZ0noxMesSnfNrSbFtNjeDiUvEJFHRGEdSYhsv/e1uMg6ubU
Gqio8pAe4+AecHewCHYxLnELDU64/wEiZLd0nYGT6w6N5fFmRIsRABhdy059
9DuSZWnNfIJsfS7RPTsLW/TrT+440X75SrLjF0zqnCUQ4tlmdEVJsA6fVuKE
pRk0HwVOutxDbqm3FDuOONarsYFAXpdYPdZ7R9rO+CdpL7rJ4i3huLdxx8A2
QxhtClEcvoZUX3B59wxegyHiI+3nqUIOD3+PW4j4a+SrQJOdeYx6mu6O77nC
1lO9gVyxUpbM3FzugVTofFhO2NO4jOaWVHgnFd6ow2CtywJqrAcA/XM21bPT
HA5fMT85+NSmCja58zDgLjj5sROKR1phjH3xnTM/CPWdkE8u6x7m4JrP2WiO
9WQIZmjpP+GY4OQ9U5MB7UQkyyU3keiroc8wVACV4TBbT/NOs9iiKYdfKFWX
9wBO/4vnr88OzRxEB1KiehzF+DDn6ESVHdstUFgxyCfA3z83VaEDdvn2X/sl
ZXj13/+oeeKTI9PwhSmAdZ2bLlnSAwyOLtkfaBBMJXW50GOWEdmN9OCtm3HK
xZjPGDNb/h+5r5l8um9X0GK2uUeUbRxSuENry/CIHEeFJ4TKFXGFxOvmQhlv
JA4A22HeUT6sAPjVUu0eJapVcHupc0clcfomVzc70GidvV52fJO2bG9sT/yy
4Evubz/vxDoPJPSPTI3JEShI9Bytsssjtzzua21QAetFOc6WmzipRS8DHK/R
jNb0o+QLDeRhsTfwCI/ICn/qDU3jxukSbzv1xq90gRz5tBpFXOSiPJIIfgGc
wqMeg21kwN26fiAltb0wugNhrYeZ+QPctukQ+4uQn/Xuw32jsvH+a8IxJusL
ohdo+rnmJkNimBveLtZatqfwQWoQgxdWtJA7WWDBr+m10Lb8pVFqLPWxcRKJ
L8waPF38qXqFJsxeTXgTfNAk7iBatvDqQdMoNPo8VkWCxeB2qpr99N4+n8e3
FwpK/nkCKsG/6oaEN0O+5Y5jO57J21g/jn0Tc0UgvquJiXMHkdNm8cD9mpzq
mVjzFX4Wo+n890d/peV8/+iOVjcZ5CR4g++OXAzTKXs07zW9CxJt8r9ZVzQt
D50rg+bDLsVRJFvuigetK+1bUXkuC5VBOsqSE0i9YUGvXxlVtZ0Xzf4hYk77
d9S0bY1j1olJ9rjgDxM52Sdnt+FFtoMxnkLSxRgf3KEcsjhm2LIPszm1oqDR
3nz8C7LG2brjMlfG8eP0QfuqPwikXELC8vEmhudSPhoirzSXTyd1UQW14uBR
mFXINtkaWoMORuW/lz5CzoRW6Qufp+OybQ/tItxZlyj7pYzEl+xiMqsUArev
2IbHkUx/fg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1JseNXRo3+FDvmKdcKVviSynYhJMOn2xGMtltX7rSCxqx8jsQNkTKdx7HgRGYPkGNC2Qxk0bVVfO4pDq6hzjKifmubXlvEL/boR2V/XHyuVqEIT+Pxi93FLqrGInnwrMYjKD2O2+zRNrGeltuQJOcpTw4VZF1qA9F3ODXqHaL/WC95EaID+snAb2z6b1E0QfsXFKvSHOb+PsUQXUwnc0Dy98Z0IQn7kbPE/+HLJcmop6q5ajOBSz42b1z7fKzxQuJZMUYAzV0pF//AlYtudGEcsEL8eN6338jLCSDWNJRK7jxpSBNx0b9/IjkGJ8/Ge6LbCT7ri2HsRmfJIZJII1IMZG+Bot9k0/OMaWlEzKYBXG+y3zsYUon92XfmTP/+duB7Hi9vHjl9hGvpOjCiHhD425/rtjZDdJfWpP8mhS+Uqs10ygJ2cknOYLpSRVDB4deLoE2VhgsytWzHziBJC3JPAHdhca+qhpYhfMWBwDQvY6mAJO4Z6IN+gwzqXzrxFyE0VC232kdMOAdng82dpmFGhm+BqDV9yttyr4h1MoShf6UDARqKDY/y8fKD0VFulM+Wf/8IhWUs0NXeDtCB1ivdcDfXujeh3L9Cg3Y6MW7sJ3dNj4+pgki0MXw9GNvm6gJIovWxfVjKSg4wGhsPk3H9DKT08YhFZmN20waqEz0rqx7u5pdVH6TwPebVwi2O58XtfpdgOqcOjzrdXEj9t6RmjA9KxzAWiergz4yLfSwkWLqjUqi99F2yYegVS1C/ymngjZgMXTf09LtC2V1lGl9AP"
`endif