// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ctcDnyy+9WL7G0ywNl0EFo0TlIfPaG/41MebRwkxvViMNuKs2HrzQCabr2dx
icc43f/pCjUuyp+AmZOpV4mTE/p8hgEAzcepGp7EIXx66RzJ1dSUd5uXZuiF
O9W16EWBE/eTpBb5Z7tljU1yI3QDZHeIr6zak0obBjLXghIV/kiQCfu4FV2O
2ppmg9ieJHR1ol1pGu+Cvdt2Da5SW89P7/+WJGViwPSiSwGwqPVQji4yw4mv
BJOomxM5rBNnmTLdhXlAEYC/DDtwmlLxlzEodvFriGykRUfo3ebLzMzhRwVA
kLHXySSlfhANMg6nB/pTCSyWri0Va66lyS6IiJcCJA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FTT7kicRyLFNdtTXHjNj3lTZRE+0MbA1qRYoF4u3bZQp5tINva4ayFP63i9m
E6y6LbE1Agi/yFNevSGTPXZZkjREOhs/2TFbBNddfQH/3xmhYqcv1sRnKzvI
s0bsQpPz1YzpGK29GYeRaIwaVMZ5qOU+ceYCq0UONCmQ3sUf0VP90SzWtpb7
itxT9TIaUzPB7B7cfvTGLMZePqlstDcgQFtwLuDMDEUeNYnNjs9yy30vR4+Q
YGEf0D+IZNneOut2QBlk3r8tluoQwYNI/9gRDttXc+PP3LNOBh4fPnweVA4E
rG6ScUB2hs62VbzwIgQDU4xLpzuk5XePaoVgNEUybA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
V+7t/c9r3acitIHmN3zNdKQXtHlghv9ELrnc/Hki2ltYta2feyfc77y9Ge/c
vyX/Q7RZx7kjmOV5yuqYfEMt0gGXBx+2+AHiMh3bv65ulgtm/0TwQKM87AgJ
fMRx772vBRRpB+UDysy8BNcLD4cZWWrrIH/nEg9/piVQbSd3TvsC5pymHP4Q
qsQhG/3bzD8JjcoADAvz6WBmxl8pOVh7WQfga3XgmZVDLURGInVxlESOFYuv
Bk/y2rlkCZc1F2czrJh4pl7S5+qdq6ehKvT05T+R2x2mOodW4AaJszECTRDR
dEo0tP8pcUk1q8J5oTQu8VabuQ+lzwhGZuDibF5wcQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GyB5KfUXwcJ118WT8YIv/rfu0PuQzHrk1LOWxHCrHqxiMFYpQwRO5KbSHbgR
erVUlNEWWhuqudk3QF1bLurEvC8qfXy8BbMZwDmVgWIaVUrnikEZefPwXgyk
O+86x5i0A2dV7I++chPla+P8Y4mRVhxB6QyhFlbMUlefw2k7XgQXOK2+MTwJ
cOuj8ZPWLlWK9amx7D/EWXLJc/hbQD39+oMeZIpMLGBrFd42jfIRRQnidrN1
CBnuRpYaNlWg8jcPNB/MXD3bblVgpz4ai97TikYsHmI0M4NnKJ5qST4iFxaO
l7NBhYagzPALh9Sx/Q9HgCYDT8evDli6i1BFS7qf1w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PVZtZnfceHcKfi+EBe8MLugmlsbzTtLYdzKUM9MqY3JfTX1D7Y0PoS56IKVf
42WdVvB3+7OeGoTgvxW+UmasCOFl7Sk3FhW2T27n8BGRYkFeSETcoE2ICcrG
A1otF/znyqL9eWI011fIcpnWhmDP7HUuD122EKPHmIUYWirzw08=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
E8Z+bFoMqygyQxpn1Ey6fRAyKa6IbGaY9lD2T1MxcHtZreUaTomdDB3PH6kW
+ri0+vQv3xOMxi6HHJOMxO/IoGZSpZbMczac9l0kFlxkDFIOKBvOI/nVuUEo
+VUecPgrd7Xl3w3NKFdd2w2PgPY7TZRVn7MvFVXYc+OqR64OTjZQUQqWgmVa
vyGihUNFb/3CbzO3LgnnyicM4Pq4yXZfK6QpJkOita0k6xJf1PZ6vNwkxsXN
eIOYlF0AdWhfOQjLzJFiVS2OVyvCOxHcaIXKcdvQlCQ1AYvoKIq6HkzrZWQT
1muBrk6IeQOkPAywr3/0m7fFdezB6yVc1gnUKbv/6GmgAJarCuOtbkzYhyw9
CU5dWBvIKkPyOjGxTiqG5jQ9NlSZCa2Yc9VCEFwxPQqAbxzAffAgZ8UZJv5a
UDTRkDnwg1Cf9VnGHmtVuzeDfAOVyVl1Zq/KVSH9Fp9jl8k62m57BJICkI35
VPQHw/kpAKg22Uo6SEM5jYrdY1c6uyZl


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AnbmTpqx2np076prcudEDDJbUi77NsIhGha4546TxLqmmPLeAtIKOjRORDv6
fWCnliOf66ICkj+qIjuzQ25YGH7SIqmBVSHqF+qhPTWLRo3iqiR4VET+SkFb
mSQ5A38G5YXJlbw4jYhqitBNRh9lqCNso//EIHX3NRFjjvVk3Cs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eLIqTsDWR9LVeSVF2JWgqBp/NWYg5E9Lp66o5DWshAQrEtOBKGwyE8zZcTm9
PDt6FCzMDUg1BUWqd21klL9o4pMPWsdqP57w2XjLI/uc77kHXb5rj2Zei9oX
WFhYr3bP3v6miiGhF8jEbf23+vfxwR2DNNyQfDLX+aKVvcQ1xXw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2304)
`pragma protect data_block
GctKK+8jPCjXQD/XpVrs55jbNZDC2Sq1ZHLNV0ZG8aze8BXdQOCQ+7Ny4mGZ
RoiwMnSExvgjQ/+HRSjuScc3yvW+kaskrsUYKv3WC4jz3F6w8MF1Tpy4dsgd
kNszQfFfPY1p2IHSx9YasKIrBKP22t4offdzvtyQ9MlVi+kmlbFbRs9CHnwe
sRzNqA3VBLuItBUTO4KmMyKM7m0KQtTiudIb58ImONU/LHEzeh4om14qGf11
RrQVnKeMYMVOhDZgnVsTrt2RMJcRs4lvYjh0gRz8Fx4T7Tb04sOdff/Shp72
4xrmaWq1EWWsutHFpqjMwVdBaeSNAQ03166HJTazJMyhB+nQWINDY7wbPI5t
rbbiXxDfxnrxZmXH42upek98XLnj94d6GJCWMb/Ep5N3wK5RTIP2N/i3RbCz
Ko7AOAHfNg3SfAsdRNPpTS+GcXafJ+u28qJ13KZKwX5fXm89sJFPjg9o6Z7C
rcB5Wd0tVbvDsYE7/rJx3EpVbEW/ZaUgWwLyahr73Kl/3KcNt9UXQctLFihx
C+AsLW/relY/438yuyK6OeGgwdah4GIxAX/zN/EIOuXx3hGfPq4wAQduE1a7
efLAN+6q1DTN4s5XAci1MQ6tkOQYUu8AELNHE5j/XGmvS/QUDd/RJd87wIZB
EQUPhwKlfKAl9yhhUY521dGDQaY+SVgFo4O5jbb+VtVsTxTwWiGYPZZe0M+u
8iNA5Jt0HudiZQL2xvved/exJGdTcpdebH/VCoSjzNwZqahoqz2yTZmRhqlp
FneLslUEgRMRUwSva4gYtXJwzlAuWUo8oC5mrAU5sO1yWnhbgsZR9BgAbNZy
VGQySVvoRQXI0l4ZSctvU/n5R7Ht/lVBWFlRCIWxSFYvjEO2ddVf3IoUrvHd
Cbse3Pk+DYwJ9ZNE/3elTHYyaYpWIfrKmOoMWk0l7sZw4l5cLMIdd8s4R/Hc
wTyBXA8exzDn9GCzoKQ209Bn3cWktaTXEWJ8MbT+cDrDuWkIv8hbMalvaGzA
PMV4+1f76H4HtaPbYxK7hPqbPfAxvyFz72yDy/y4Vv8xhvznkl0LtP+i+fbC
cd1D3kf4RMvgBrjZmR3to/7Aln4904ctHiwjtLa6UOib50ZJrfoJKzR3juHV
DPW0lJpoRAmINAkYb+cYB10+2cLWCos0x96spp5C2rsqlcN5y54mAgVQ6lGo
UYUzpoucoXu9/dJaKIct5a3KT5AyyGlhDZ+sjMeHvHMttfWuuEM2wldkYrzK
/y6cYlKAMmfdX+3WKmuUwGdHo4zHTrvF3L1iJSHFUfnGmZCq1FTERS0VJnap
qYvwh1FLrz9aItLTTN4wQMw4lFn3wMFxt/EFYdMtmC8f5rzoCxoKmihLQvA8
8VEiJOGPqUn1TZan0GB2ndowBHNIBZgo8fDeI3IDDlXlh/pBA++yOFfWVN+H
8XwY6cWsC/q/9lebVXfSG1NSSTBxbr0yNqhnbPT06v6Tb1IvZOsUbQWVGhSq
/+7u4gweIzdh421760WVQKLIvgtIYOIjQGlUGkIPD2t/oo3bQNbu+TW+wsW/
F2K7p+dLa5fBPfpcOfhnWa9qkhbDlGBxwfTZgQAE+0x/kPegSOWgigYXM1eB
R6NxvUzZ0p6biG/569Xm8tA/Uc6moz7icbkPmTPbDCNswOMhGfdpJqi7m0l1
pxrnbU5leq/YmPTGQ0JWukHXC9A5+MEU9mgRv2Do59zh0qOvdT6QavnY+86e
cNj/qyJpxI/71k6gaC3vvoK0/WsxBkY5jDSfi23Al4t3C9oO88TLkPip5VYh
T/rChTy4bg0AUQGJxX/lpYGNIFc+LrHWaL2SNkR+6ZtUHIZILledSvgf+uXM
9iir4CYQL5QIwM3Vs2sGEReOKS+p4/0YXQAp12eej/bIjRVvnpzpflzE0g6g
MBpiCev6h7XGtr8w9AK9cM1cZxxJEJyH7qW5l4sA/QzinmCxFkcoSH4iJXw4
4FvzRD6aJWD/zbTYwwARGYVmAaaFphT+Xy3FNukBRC6W5KyyjtzF7qMGcz1g
Utgaxm2rqL3zt4Im7b0FDHO28Nio9Sc8vKJI5VDNksoSfM/boHlF8XKz/ay3
Xc1Q2Q5MZ1kK7h5tlMYPcKRQHDaD46+uQ9gXcqPypVpmQEzAsWuagM9SqnEO
EcZrLCgug4zWtQvWxhH1iFeEzQAEH6iFbZTTJ/jtqGXxOEeV/8eza9musJ3v
u+MNgOlyfnaa2yEIzQV7e9p7UWKQvPQBBl/5H0y7lViITQK5EVD6FPJJy5Y2
0vw7tQoHIdGhlbso0PA07G2YR8aIRqw/EX0+Hd/Sor4h8LhAlTX7gKMLXaSN
rvtFq2BW+R9cfNkGxjejAHaa1LbZgmcJ9Ei+NNo8MAuTOBNw4qLMO7LoUJAR
9dnIQPCtFDi6JPtxV9dR1BQYxVMpCLn+IIp76LHD/e7803wom0TklZZfyxFs
t3rtQaSKrBAludLRW8xv93t4dD4OOJE671m/ITQmisIwVfRFWd+vptRqRVuM
+aOwVJozfpsLT8uxulB+B+sejO/eXKSCVqMxkAu7nqjQx+50653CQDo98Q+o
+gV8zlHk1f8OjSVLPCQAc2BaMRHJDPJrwsYjVnPX+x4tDth7JpvU6nd6Kaur
LXtPqH/aW+C1CswZHy/TgBWQAzoiV90mMbDz7MfBtOZNF3CN/U1ntBmgjTK3
OtAxXA6pSAzRlhc9NbnCe4EskVgNy6zLLG22RKpMmu1cd42f4Y57tJnCKF8m
lZkdlvVqPGJFMLQpwFxYIaD4/iCsO2GV5WQ6IZ/5xALmVzdkTylynS6eIAkj
uSFJM1q0MWMLzPN9FhF5CABC+1RPz7HX/X8bt4mxAWhNhJBNlbqpWIB8aK9S
06ry2rtFNpMOYhoYPekBIXg+u+Qi02LcIjayHXEn23t901aFkgzsPHkUZY55
hhrNnNr+6wziogYtAh3nBebwil8nhyn5wcYqIydt+VUV2W+3XH6kbVS/y4iA
ShZROclqQjVj6htiUlmXy6GWGrqMxW7gwxtMO8rNqOmz0Q6Q6zhJ9qz0O6UT
0y+o/UETDgWQ

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyI5h++oL9KGW1ZMN7ibhnsR/kMsWeRmqbte7eT4ymkaTOfKkVL2w99Cpt1nwo0LKM6GYGKYZYwphDJCjCT1BzJFGPcgTUCaBNw7Ih7vo/g9DNDSwDnb02q9VieYhxdOoJPT96O4Td5j8yM0e/q5CuhnQFzHRZSaNlG+o7ahaiusZr/BGz7cRTPtT+V0eOZnu7bexady5685lAGDRCS7lGaFcNxll9COGWCu/HKwiEHsTBSEiQiqfWzG5Ff+LqKd3SLqbE0MxYhH4u4awGNki4M7ghGs6n93B0eYIXSE8reRMI5tVpDCtmJcBCYfdZFJOLVMYKCwS82KyC8wvBtWbypxwDMtofChhMGY/5N7po5oXKjGm3ydY0PYe/2Ol6ushl4sSyZ1bmoO5oeAEvY7No/s/BdF2I2ypb7lLNE9OgvFG8SURjkLkgz+NQuVCGduPfxZnOiRJwLss9hqROQchylFTAab64H/K+nlE6qHZ1Om5IRy4PkVmR3FhEuX24g4yRBoVXiQv8U60SmJAksrzuJgTVYh1XMR903bP8vf1kq9MtvJL6BFJpkuuhkgJEhZKC2leU27cACMttiBqcfBLWA8o1dgKg0W9psYL/IPyThz23dKAVtEYsg/mY/Z0XTIzyB+Ci1CvWSotbcx5rD7t4xAPuDmpmWdHhOvhPZdex2KxYQaMNFGVFaa6Ajr0oguilwvg/JLnYSLlzrCHUk4+IPv50FhaOFpT3XBwDixvJ6nzdCotq0gzwBCQtyjhJbWhlZ7+Ye8b6dbKoBk+baATuL5"
`endif