// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SqbaK1HJbuj/vHB5fJtVoB0JXySYVYcXMb5pECELuea5G7VVQApjYD5ge6Wj
YvyrP9cuedjVMvFTAOGoUdg0SpkwXzy+1got6FNQgAnEHl1nQvYrbiuWOL2d
mCt2HVaquByrBXf/p93aSGYbGiqFzewuiFsFD6vVy2f44Tq0JT9EiNO8VPPv
mJhkPeQGlVAZgFQLm1sViVLbB4HVh7pQZtbTJV3n7/omYF9xERo1rsaAsMIo
Y/5iV1qghfeZmAgNa69rNs02UsX7MauYfNnKG8UAzeakLTZ2O69A3GHl/Sxu
vSu+XntlffC1wrHhKHO5tA0hgFfmbZHlFhBe0e5paA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AAyiQBzdwFJfrTbNpGIysVfxHhKx+3J6/OOFC7lhaV6peMx79t9kRKTpfRmN
N7qid7HIbSrC5APXlJJbs76Z/uToMwNKq4000xcuO3NswUxAkO6jLMIYtjSj
vqa/r2GD7XNIBMjYFP4oREuXbdTI4RQpHugRa5I1fsibRbQO0GXPHurfCWN4
mCo0gzJJC1eIgwVAwpWA4MNSaQOB3y1//DlZ5NAXTFJsXUVx/8PXL5mYjGE4
w41JAwEByvMQdNUKhLuRONXDrBKBR5taWpb8odidcvM8+C3jxFMJFxut1CVT
Ki1ebTRaFw4YxRD8dXRUDnB9au+GLgcNeYEKHfU2rA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mgobJjx7EgmMUxuuU0jjxhOvE/jQ7UAQwHPOpjSeWKMoIaqzp3+4MOkTZt8p
vMqySUYG/bAU6mlCNWwc1TpskVsrCRehk4TcyfydGmtOGtpkBpLFY21lOLod
h+dNB/rxQi2pU6hxnHo/TTak16EWNOlLkcy+Tqb8aBKt3M2TXmE8HhDTp6zQ
9oEd5RaljGXKEBI3pw+tmUwytMgt7ty4pMLkroKbN77R5upGeRT67D9ahiRy
Q+M+4Da5rvf87rwKRQ8YVY2ftKvfZaeZf/O5xZyYF6kBV3Ut2ZHwc86H4X5A
tz2Qyvle9tAemMy2M6Lso8M+9Pmu02ISrog9yW5OeA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZrbF6RGOIhRTuo8GmUUB7KSS8MSFvEkehOVRyTpj+MHCYjlvmUFtAB9nVNnj
7tX/8BDHl+wk7BFYsyKIJ+knZ0SlaYarBsW1C28yHtmjISaBdWDfqs1PhHk1
BKr50p7Ql6I/9Y7YgyGRL1NJ9vtplyb8sdv2H9xzMt2LteNascbXfb8orANA
5FP2m0JMMTddkkV4R2VFf1v0ChAYpJDvRyvlNf7S3NIMuhPLdxvQ/S9AMFN8
pE1e+sVu4mVPkYt7WymAM0j6UCXqFy1i/jUpXa7NYH4GK92b9LVK0NQ83oJX
WyU8bpBdI47q7WUXNYGFg1fqubXUftquMjKBK1BMfA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DFuMhwquThP3W1cQPvbG+eG15eQJRnOvxywkk/sR0z7e1lIGnpT9F5O6Y9m1
f07dykrOAg43AdGH5CBvsxXUXXmrmVAVQfTYNW7B+vFFS2aVkrNlj0fxSjN6
QuFtH3PHqOgv13NlNBsepaAdwCZXo9lZMQBIldgG/nVv/PPkNzQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
MMWRD3BxAvXHjh7HrvTontRUpeRLyYWBq2ILYEAfFunBcKIh5LejItCFnIgC
5DyYKM8KW8iH3dw0yAuPXlvyJlWmE5ylXiURnstzBsj0kRALpvJMafRAbued
rndQAi0b3eCvR25tTBxc0MiTaKLlTUZPNKrOhuYoQLVrg7ut79PqgvZ2oStn
BV9bEjkZgnicAnuSNOkFWlwJSLRChU35TQN51PXb2xKZQTnQ09e3jIS1HiQs
lCuge639oFsT+HaK7yAlG9MX70XK/r8/GKtFsbQIu1pqaL0RBir3daXNU1MW
QIYMuXiQdTlvGso5NHjqWzn4o1ROT265Ok2S+Lfjb+YIn86rMWs815G40niP
ZtZmDHpjViG8j/NQbwEIP/1DkUJS7DKekrHzuaAnJyVYKRiTaVbLLj4FwdxK
KoaO0nHMCzSzuYsLJi7UJUrbV2lNcacFw2QqrwgqawWMgkyQ3x04MTRb8LrN
wrTvcK5hpI7UYGxw8s6eRdl4T7e0gbXF


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pNx86mepCJPwlInWP3OTepCzvMjdueFyfz6Q05dfjD9TDxPBkAHpXWL75ad3
1vCDR10fNhvQWRqhPjBGzlBUgBA/6nqasOvhbL5XVWYhSjaqUgqhFve/PtX4
SqRFm2vSQ4PSbr/99Os8m8HVH8rYHy2hQOtId8PJF64VlpcS8hs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cEXJmIk56qPcfQjo3ddVXXXmDVar4rR9AO2qdmTDniY/h2B0T09DFQZBTPDu
IJQ3waTTI3ewqVkIlEb00CUTlgrFrfW1PserYVmD0y7x5Nq/hRfyiY19k+wF
veKI68r1/soZXxV7tw0ByFxENA+Qn4bPoWni81KQWJmfg5VvKJQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 66672)
`pragma protect data_block
zKJyp9pTRxPkqe/Wwj15ex0MGycdz/ZOyhneajxUj+bjYgeT1X1wLp/z8LAx
CezFIsn52LxIK7GtS1uIrhpHC7UUSQGbrCc3E4kOw82CAtAti+Q3f/zWUCVG
8+36g8wHo3T7efZqDJMC6TsYV3YNCmMm2+nPLfTm8h0PRPMSpt73arBLFZ2w
dnsX4GZqAVPqgHmjHsH9UOzMSWopVKMhRi8WM5piAJ5DJiM3GJsb7s/lM0c4
d8/WCpGgeCXHINDhkNjxtvyQlMwd/enbCMVOB8OrWIbnW2U4C6ahPTSsqawB
Rd6vdt8PF8ALR3aNhx249JHUTVqXD/+WqaOE9aD0plWmyJZKZ9XGWlDl/b0V
IMORyBkjf/Iv1F5uwbcvso2aD0TA9Dhu6cTut/MJhvyvRzbwcmogEMhear4F
NFchQIHcnN0SHY1s6Z7Ia7H86ues8m8i/vvfD07gwOybNqBpnBdeQxJlYt+O
l8x3qP6mYJbD+pIvXghjYZAqP2mOZXuiwPPXf6f8aEbQvx+4+9KeE5g9e1uX
1G1Zd04P8tNzpR6aRBK5Krw4a4YWxHGWqMdf+OjoPP+epTaZyuBnoOAfTznu
FjdSmCXBIcPmBRXVU0z6P3nazCygGDpl+X/j5klB+iH1F3uClefDnQ3F/Fi/
MPVgi1emp+/Itv/JpVd0DDVu/6oyuU+/4EhssS/1iEbzxPUwPA7ZleUB3IgZ
5WQmJVPtqgJfPR47n3xsyBkrlIP0WvQjqKi6NQ1+y1mEvMGSCRFqVyKaGLgI
VXpsr37TtdtNdL+6HYVUGwfkg1d5GifD0ZPhvVfA4rkCDhaXIq7dMvmJaRbV
cIHeTBtW5Y4che/n3VAZTg6ETPDz04J14rzVN3+y49EACNxn3v8Ao5wLchAL
zZl4RjjBi+V/ZJFkPBP0o+h1u/BR39dWXINHDBasD/LK5AKR/qOOrVGkQUvV
AQN2XDH3TdKxZ5KbjZ0In3eMoSrlMoylNPEOGgHdAlxk44BtpJu4KtETURz8
WzkIMfykXeCpJNdsYytYO44HR2RiQBgR53D4gOCY+rLFJLW8oxITLS97qmic
IIiSMNrAG/RQtIxAuVKtL5DYJZIbgnvmKleIOOtGLlUfxtGDLNLm4F/c6Q9J
yaHwwLGTiCsStYyzCOnRnXlOc75euNRwXrqFuao/ewYNBPR1VaX4MK/7TdCX
hPguGIQyX998Ljd1UWc1j1JODynKYt06/0mJDQVHLoDuaHHHFr0pyXEhUMvC
rE/52zsCTfVHMC/7b4mvt31/Hrq7irJhrFr6D0vyvzc+11MJ1VdDfW3j8nuT
bxt9anCewK97A7ZnnWJx/5dBAh2iv+jGGbKrPQ7g9T0rlgPcJOahHLqb1XeD
SYsoSTGLTzlDxc5RMZyX1uOT+RIZDx0BLx8k42+A9NLRXD7GGnPPQGSI8sqn
pEh+bSbldzEZB7oB3dV+lqPriIeXniCwp7gvmtU9cE9bmYRE+Q0CEg93kmgH
+/hUln3CyHl/8MkHsRy41VSMfPmLgw+B/n/cZTdsMn+VexdjSVat3k3kRwza
sS5cp44ZfEKRcsAMsTcqyO4bEvSNtj9JcfSoYoPJXWdRNlhaQpLu7b0vFFqi
93Pousl9gfscgMblicqPezmNKnifswznKW0Z4lPNdiLEd+Fkmmw+WYT5jJOy
ZpbRISdWzwMQ7tcUtM8b8sqEgcZ1EWqEU2bndEdicIoBL3HEdFy/cwZgLE7g
LKbsmyiHPcuulYwldj6wORYGeD2J5Zx2Rs5942+256bkT4HPfLTA3OF2gAUQ
9cC6mQ/VUQQtvaPT/MDIbtHXwsB99fOEz2aUmSB0aZXXFZ06xfaHd7Qo/21Y
SNraKquKEsj+BXAAZkZvYUG+E7jreZiGGAygNIvYG5CN4gI0ybYxtliQpCC6
dl1mnFZ+ytLM33Q/z3HCQBGT2o8Cwsw3XTtxgEWKfKdQFt7taat5rG0M8WMj
MLGbrKmNVFK01Efx9016yU8ZQyA5gkccARcLM3bevXsb2BF40iK3itj2Q6pS
JKu8PipwRf2k6ec5h+OoXP/sGY07DfeaEAUHW0/61WxH9o15IpGHwjS/H0qO
1vyDqsUukZmbOztxhWAoAjG4BGHOtMh2iJgWRAZirxJLCo6ewLriVb1u7cuC
W7mN0aOnk+WE5X70aXIlStzebd92qsArDGasE/iQPIykE5p/cfcbeLUVIUQy
g/BPL3bPGaxpbXBVW3Qp0CnNFzCxeqYBU+/ls6YgJfpVM1dxSIFDdA0zQEG+
qC5Z76HgubP/e2Ki+7sLn6yoVLroguzwxbhhCQVPvcCyzUHK3fWZgYjDqMvD
g7WKENqmyEkQr9zmchQ6O5EsyQ/O4hdpQ6PMHWAZ45IbSNmxHFY2Fy+hbbQp
qI3S9tZHVHbpHOkhbUdc5wcxAboGdmxdax3UBwSKUoouKxf6HUJFSc5+hWqC
qLU5xHTshFwQ5Ld2wfcBlxsQTdY4oKqdH0XjjDStDHMMSCw/RI9pLAJ3eXUN
v2taErl425QPLhuivQjdwr19Ah7DztTvWB3ocWTh2kfG46IzU+opB8HgsNMt
Ns635AfEMBj2f9pXsPkyZxmxnzbPgkXO2VC54AW0TGs/9/ajuE1Rq92ywNxX
fv3+OyobEjbYetusJ46sz7v4HDewoEPfCE3bR65prdCNTUco8Yr8oW44L+kG
cSP5w5tJCM1I3jUf/m2Z8rnaJs1edPn/4kNwjusZhju0pZa1hEn/ILgx2Jh1
6MiVaGkUoOfpocZ6DFQQsfLINKmx1EN+GvYV2B/X5HgzPVYqj0MzXigMKiWZ
SCYR/aNOdu6mBHW8OQ+MNBRe1Jl8JcdVuWmXG1QLvsJurlo6OwD7ugptebJd
elX5qIm1yWYpd5/q/Ydx8TrjI4B/OuvwmA6CiRWfolt7QYaLV4ATigzdyDao
JjO+3CUv7n0ZqNe2N7F/Los8ditw7SGeB8cY/7afouwzx09zoe4QorQy63kx
lqWWp9+UDYso5NUDJM1jBqTn6HkVdqa/TO4T5/6x9U9sxAcrr1pMM2qCKOa/
xKdgYZvoZl/+6l03iJyDNCKev9YQjQRqmvMpqfizW8BRiUOJkBvLiRYPQZxJ
rsvLQ/tnLwGqKYeEHeAZVOkEMO5Qirsil+nKj+XXR5b4OZvSULqrU54hCij2
+vhabb3208w6cy67hS25KDaOj2upZwBoAXRA+1fSCi8QnV60N848xRT0Ks7M
jbd+KfF8Gkjbyxr4o4xlr0mKmDwlfjx0R+1KV8KKATd4NuFN0hbZszQacUrT
nfkaCiuMuJ/GVA7cQx3sZ7Cp5RJv7ImOfXoxTbGmMqxC90rpTPDfmHG9G2Sq
5FAHpqHBwFUSs5pymHjKX+APisudgJcyEHUZG+Frf4+cn7PIwVYUaygvRkOQ
zRU7RfU1ew+qXg0UhYJhpRPY1ItLt4oIDoTcD5SpnYtV4tySj5tYYEshR8i1
iwoo8EvnU3HlozAzuwmF9ltJrX6tgokAbteLe4ZssaP5wRyqP0mtdywPLYH/
re7YHM2iaWMM0lcPmDRs4dc7hwq01vmWPfOASyL+LrXH7xf8lIXhX+nBFBB5
PIFkM5eU05alxepYEpcHbbTx7gtM7UTenHhSxbanIFiFEUZ2ogFWvDIA5qUO
otLoZuPXW7kV5oxKKbkQwywbWCH5i3h7u2inK18aaeZTk4ite+NAIGbCCzgk
zNusOVwaaePfVdVuX07vszXE4ZUw/4w68ojBtGX2u7QWCdDzFEj76WHNOgHZ
9oBBpAnrm5AbZQKmhoKtoa8u6x9UirvbLr1FKNoA4PARHLX2Gs+qNqBCnRiO
Myh4CX87q66h7zIqKB00i2dbki7Je12g8zNILe3VNP4ARNC7eLTkr/xCmeac
ZHkLuOv2bUctHWncrWCWCzCMWadIFxHOxNAO6ho86gP3IgrfLH/1/cpHzQVc
3KM2J8lsS/llGRsR24LDyUwFgg632SLO9vScVDX7X+5pfuvv3WPSjOJNd0Ya
z4Prx5NhYkc1a7txqNIDBtlEWFxkinCgMO1osp0QPTOgRBJ5oaaw0G1ROiTV
nCgbDv/7ikaGyR0hnjwIqxVlGwqvrZ5bFKvTRRjdvRpM8thwydJmwuVlC9i2
3wARR6gVlNgo1KHkq7WIaRBC1Pm+K+yynSoiPWq3UT9q6tkEOgGiE9DQ3Zrz
/vn+SS/yhALbk7T3Lk7AkARQhWES3r12CNCjAo8P2dxSQlgVvlbAHNFFGjX1
JL3YHgnyc5msoHsACkMedx9+bKHYKKPXUIZylXuWvAVcn++I6f7MAwlt91Bi
0GszJFfLdux2/grZ8MV3Pg2DYnurMVayR7OtT6XH8XjTZ8WqWpUzrLG3yOBH
TiVgdEIPd/MONUY1TmJpoLVxsVBQGuxxNVmHbRQsrrwzjvygsxqe9Xz1ughw
ceSvWTEo3MVqUaIVlGQDJrLfgzMFd8tAm1+v06nGp1uQo8A9u8unWQ5y7TuY
X/iZ3CpY3oojV7/R/xw9TNZ7bQ9ZpIbi6H7H7rKuziVLJXU8thJnZgjhPb1h
tQkCKGLisuOo2YYNO30rZVOCJ689MF5H3Ywqz2HvPZQG+JbEpQDp3ggfZPuZ
Q+Z1LVF9FPkllswm6OzUz38zS1OBuUHw9wvDMXnhHa+jSC2x0Eg9hqzUXP/U
qjE1QkU2h8YtZiGE02M+kSYqVzNDnja7JfOM0KXMIVw6Am+BZ4NFwF4cs7Ar
0ipQlx51EOOckkVf3nywyEhE3DF3oC+ZCBaPowF66T40FMY+xjTsKHfQStWq
MFhj7rjQmOFBiNBNGf1RDg30vZtwR5FQlz78hRJ3sSViLfGEMBdv/r4vmNGE
1revj+pTjUpWGYsrHhw41L+NRGFwb9YmZO335rIgiCJTmclH0OLdXv2u/Xm0
U/2WLEVWHQjnEvJpT3RbVPnfP6aRcklrUkWeAQrIKebAiiG5o5Im0Y8RzV3X
QMCReytCCwP86vkgNh0XwRFqfGbMplNZCEpKloWFi6hjsJzCSA1aA5Joum2S
JpesMM++wjkYcRSDbdwLeV/u0vuyWMR3POowpWcPv7iY3ubaSecIqHK6gagD
CoVgEnEPbszJ+dRFuM66AQBah73XMPC+gx53z2hag/MO5HLdCCPyulBisu0i
nzMatjHaqo14W/plBoGza5Udg1IxCoUsYfLpCPwkC6zUjg1Plg4IlIx7k7d+
S/W7F7zSYXQT0iFsmC3JkX0CI/HK8NsrrcjgDKIT6Ms6ZuggUb/loRA/4Ecf
S1CWwHyj5S+7F0QzpekCxL3Ft1XtPF19ydRYPIbnfxBb9bpPzM5PB5QggeUj
om8xa07Li+JcD7vOFxemJX59nn1nr2eHkhvEOC+BKJpBqQyeF7fbb7ZdGaCt
VjX3swMcneKY2edf+0V4cps0fZm3HwgZ9yG0+9mXvRWuy3BcdPdTbLJnWGzz
hnMBmSPqLdA8qWmy++YhPEht0Eko/DPuSb5QzW78vj/krqYTwcOFAbTtGUoY
gwiufb/TIsjJqr1KbgW6lyWDA6UjWU0Uc5+wErXX+glVHJn7Cyf6nO6zYQkM
YhfeYbdDEtlfrEkQvPZwsu8tQeuQLKxO0wbH9T4qyLq3+3EqFuJtn0hQC1Pp
7ZgZ8srp6Y2wQC27hPKprfrCOyMv160bmsfciQgDpPEdxXjP7yH/Sg+4AhaO
gvGfyj9xV6hJH2zy20dA/xxwNp/7Ksj4EFLU/knnwtAJjoMhkyIcmr4Lt6bk
GaeYuAAuaTOo0Z10NFUUNlc4/JHRSin9KBN9WqLTDgd8du10Syk331VfTCuo
eUovl0SeVSgUfA2gmyI91sTFxS9sQAckv96/2PphmASaIHFjgRZLAwtEXFYq
NtkIdJWNotYd93p4rg7x5ZLHezUDV49ijTnZol7g59gAE8YZ5ymPcPGCHQYC
84wVL/lEP1H1Fw0GZDdKeXMHdzkFEgJJcIEl3lNGUrEGdH2ky0etKuYJwFTh
QPlCIRAjjOMfnDjcGc6YH2Q73NM1vfi1dp+1qiRKPa2KoreSnVsGk+OSCIzV
FUDMeM+avFR0bn4U03aDU6U5G7n2s8NQNs3xrPHvNXn0k4yqNyjKylYU+rWr
zir0WNUxKUPEifGzdNx9z3YP7WfWXK4QPnOuAajZ81iiKmDncGrUvfn+dcY3
78dlYhi1I2amIWD33fEHEr5wigznkH+42ydt8NHDKGms9XOQ/4BwvbJK3zst
8nEF0mn99lH4QS79G2iQbmbLomQJl66NbeoUUiSrTtwhYsGRGWVe72p43ud6
GeZH9I8W24ZNEGLX3aUKiim9yQnIDAjVU/OsOGGkdfUjGpa3+HwR96S+c2xu
NNNmnyYqIdK6rezi1AovTfabnwXbIC/6jYekYwBdcZltkHm26ww7e77HrKkt
2f6+VAI3ZReE3+312b+L2zXr4gQFFw69fWjH5HOjvMN0X/eqprnkcAsUuGru
voCgCmmHo89Z+8vO+bKSTW9CtItWXct3qwr2VXk+O5q1fnz6TyikAGz1Ye4K
6LaEjqb4NkFuRnAfyHeCesPZGXGw/OMmz5f8j4xQPDPKYEusSBWo4A0GvioD
7lGQUBSZDHCP26OPJuKxDV5hDYx9dbiQltlJI3CRoCd9ZyFH5PZQObIttlB3
kaPsa5I0INhS0nlJSYUr08w5xPJUnZGhndxMdyn1RZoni99swXCmsfGY9qrc
fxZCm5fjIHVp5f/WPI+cIXT6rvDZ9Esmxqo6IiVgie5ZDvrZ91U8TWQY4HuF
xIUV8PX066isFOJpZOroMPCX0zapitb0ZOai1wBmMOb5LDo9bjsufvGNMvzU
JHIv3A0T9+g9WXM0n7Yl4XmQ59Nye1XTf5Ys0pAQ4V+FWjjXOD7o0raCujxM
VSWCr/YRgojqftif0162r2N0I+2Z9EdlWXjbDNBhd2RN/4YSwuAqeOfA3I1d
d3kV+ASDXRChTLXdwVMPT85SASVcRjeKBXq9vD13T8LR/TW85v+3NhvI7psQ
udfRY/WRK35LQAEIS0L1EVVZ6C70q1SHxoNHMpO0FC486b5gBrmTbako06xy
dK5kbB+z7IiPUySuumuVsk3wyTYQOFxB7X7qy9OakpZmyw8OI11AkKJmrzM8
GxYFHvNdKE8oiHYUGFqgk3+lSM8eKoULinv/4G/Bf/AKTiCyoZvbDwm8DQHa
811E2i6VucpCb5fZR1hr0F3zRe1kMXBPLE8aipjbcghecHGYu4C0PbLXIMsT
BnNO5eN2Sz/51z6GDYd07hiSCABRx/abNEYTVDpcWlN4BTO9MuLjBVD8sz4j
3fMNJc3rcn8DGCY+ep88UcEsc3Qg70jWrWK9Dwc4ZNkz8wnqyW9m1lzbAQLD
neTj/NPKYDfGPMQ+V94a9Todr2ry9OmPXHInsC0A29inVIyT5ltSBkMFbNe+
ZCDlKMGLhXl+BwHhHf/ahJYmR58LFqolgk16rUEhiSKDHPsOvKWUKmeTQ00Z
uC+DP+A/s4VLCKLwt2a5f32D2ISZqVOYqSuWKAm6GvVkk6BoI6EuzKMzARmf
3LZ6S0HLqe50mBwviD/NdTHWoSTBvZ9xhyVX5WYDWQduWiUzrLGkdjN9XoJV
R+JPFHnKH73JjbEZXS3daZdxKYHwZrhEclLqlMagYGy2D7YdFRKXlXtZYYhn
xgifNgU1fQkXQo/UqL2WDBYRA756/XLdkaA6Tde08kBVorJSGn4j6mIlB5nT
/Pdg6i7S1wh4aZBEG6A5vtLAyxtSoB0pn99vPEkws1AG5RPuegN1/1kJplgV
g0s3NvZKRI0i1x/DzuX4TaLaI/FCBL42FfT0Q97vUOYRIDgqiXOhz/XLZek8
aJX3eaA8dNJvFfdzNx2Jbt1iZfEokKl63DbU/MkthTflDW5Q2XlPMPRowVmk
RmyD0GZhw42sj7pfhszKdJUEcsgxmMxepqj99MCNMBz2jDfy+7NeoCE3ygZG
aTrWsObFe7x+Mb4d7b1lCJHn/toc2rDCV/vBcawmEigdfuk1W8TTr6VJ0bpv
GTbGYEL2gN/wzNpSK/ehfe1mOzSyXxaTvmb1N95hHHqir1f82/ncng9LmtkN
K+HxkfagBmlFvJ87Qw8Tv8/oHynbHMOrA1iIJL5FboGSrLl/czNwKaTrj6jo
0hR1hMAp3d02PQt4Str0ann36HsxQXmCNiv/CvDJNnufCaZPBzLCAF+jOnaD
9/Fmu2NSrZza+sWimjlTVrWtkhI2kj7unHbP+9CCdaQ5Gppo2DRJLb1bzFTQ
I2X2mPwOHBWcob6saA0xjPaxkCvWWapd5M7+Z4FDyKDpMRhM7tEqSA3QlVF3
m3CQVIzxaGtOnNR4/cQOe3iQIXCe0Pk9m+iSzpxy4Bnt34DUCPWcYIRhrG4v
W6Kif9jpfuCbaAowUmnhMJ6aQuoXQ/IxF2tdBGfxWgLxhQQU/jfUOO2j6d2y
JYSR0eUeS/vLV/MOO+I5CzfYHDPT2Mjx02rXPfUusBF7d832aqtkWjb/GIOP
dKqAMO+wHLdqw3Iw+fTClVTyXMlHUbu8J7RL96agQ2gA9AYTn2W7WM2NUuuu
1jQRvrtNfFXvJMK+A97eg1psDEHlGhc4kTFgT5tMA6XWY1AexEW9epkadJyr
gAJFKslWi3BSCbzo978esWFs9oOcwVMsFrkwWfw8mlBBKmVE9qi3DJ7yBFO3
1D5AtU3w3kWdUm/8C022Vf8XhDnjbR3m7X2I+95JRtoqD3o/IYOiJHZS+3Tc
ln8bpjvNIsLvkrLlP1IFDymub4ZjgbI1QcyWHYn5IYwYzl6P7KbiMzEv9C7x
cimG1mRywx2Pisnq9kkd1b8QMMKy0llbelkBav658ZWAxFuX6VOjUd0pPlIw
qlkOlaAQnfhcm8WmYXVNIaRyRuHZ5zYmpsk0VvWLy3i403OxlGMUgqZci9R+
C3Z28OZCCGMsw2bOM1ghNnweBLDhym7a3GEeDZdUPxvz4P3C2kVxow4HtSvW
Y6rvSXQwJGBk/B3NZcUTy7gD/WSKcyUGuftOM0shUVNCWVON7x2cy9zUvyN0
gj3adnLGnZTFQ8XAEUEzoZu3/n/s1/2SUGU/59GaKHufgXJ+qsuAvAW6uT0a
nXiKcbTBlHXULs//AoPzoFsvnNpRpxina9AEoHa6ox9z0g1fERY8rtPXCtRt
xXPbrokdS9nwWK8nCxfaQjWeaMajnQt4ky75UZdm8hrG6xUCekZuxQm7wQDu
JRXsyqOXmVfYc/prWwlEsL4iKhCyMZnwqpEwXd2w0JnSeKSZlEXRWKGEDTDO
WyK9XguChwQUx4IBUBUzNiulyZlJH3y+566nQfPZHfw3A6BV/+kUx+jUBUVE
ADGfgRab9+liPvNNW+izIAwn6BXeHFnye9YYMpBWBzZzcgVPTBxAvEDIRzeT
D1GedALQdR8wdkPPNgocg3LsKiuxwRvnkjMOVsYYNGSGqvCUVXBrlKIX2Nju
dQlUqsKNG92efMfZNjziOx5mUjniQja5WR6LUDXblaGZoGvZqAWu9i0BynbA
hurdvA06foQvEzfacXet+jjXlSJhHOB2VHpsrB3Mc66Gj6MBN/y7OBOKisGL
AVS7LeF7FU3XYzFhVaJunVFGBqlJI8iwVrZRYmtzObLOK+3Vs9t5DgQonqO0
0VC/+CyGpokiR43PEp384c3oNV4g/fCAoRG4ytIxI406Z1Kq7F9yczdY1ecQ
Xy6kX0iwSR8n0sz/Br05Dzg6VGDqGIUE9yf6m+XpKzARmb5yEPdmR2/F9Msl
2Wr5ER+OcMHRWYnIMg9OLM+exCQIkuWuGw44jq4VXS3DY3v5X9+3/NTxJg7e
7DRdkW0VtTCeiY6RwlXn7ARTC71rO9Sfz60t5cgWDrkwWXYWvROw3hVx5nlv
Zx6njlP5tlcOv53CQnOOpZVhTD/0NA1cXDibIUqLN59rqdGSpsmCVej5upcH
05czpmVR3vPVvNfG7FMimmfzfu2/ByQhY2pOfKXq6IX3Z+O7fJb+FupuSNus
kkhxH9N4aZQjKOl+DEMmao56I8mXbi6DtpbdyAxcKU07YICzfZ7Y/O9wUPcN
7kmJbVC3LgeuggjX+w0JwBWPkPgDAnR88K3tkBQtGOhb6nZUtIplT26AmgEX
UxPWDZ8z3Y3oKGU+GpIGzIYJIu+OEHEdSrAHvhBxpTAdYCjnvQyN9EPtobm+
PK6bzlYeQP9W4pOJnmhto/ZWcdLSaoWR6+vjs4YsSSUfYyrHBQolFDqCQkNU
fTg274XJaqj1wV5VSg30k4IK9HRPINu4S+qe0IFQ7/J9hPDIkXfBy8lfyX0n
TRBEHziTl11NJ/0LltYQN49tiEKwCiesKU1YImJvImJ8c4g15wdhTgCTYNoH
Lk8wkZUUA6OjgBDPUXHmfP4eGrB9VEDwQ4/iv8tLbc69lIU55zNKmaVSe0MW
QtQ062J5whoA+YfhDMp4dCSXaVahvNz/kfPPI7R5YWw6HgBfpXANO2G9HryL
Wfh2KOjVaZoXnThTCFsS8UwmLZb8oWPMlH6Ey9SriD/1y19vwpHIV3nF7Wd9
mjx4SpfUUPnu+bH7KWhVUmQwNRsErIh70rVvAhTWrgkDHm3jwaWmObyUXVQ7
evmh+QjEt5+kgNoRgGNbq8AlVWxY+ojPrOjTwssi3q/aSLtkeAFo2tI9GkEH
Ree0pEHIBSAclg6NanXKBfJx/nkblMvIhf/gXYqWyS0Y9yODGbBJcVcRYFRH
MvB/KmGL66qT54uLlgdvp263IXtUZ5+DoQY/gH4qky7B4JvkYbv3rih8FOsD
7/G9m+b3Mn3NyHWcIg6aPJVLdsKSh8LlgsyB0voKmC8x2rahTv6zDxSVVEZU
V0eJBqgAOVZAMz2PSCV+0WOc0qcIJmc9jXn2HxJFt54o8RSEjO5Zd7JXy61L
N6HPk1TjhG2mSujox2QckIJg4TRbRRGJi5xO0cJzg/0ebIzKrFqxrpe63INg
2AypzXGPkydi3k3h+wxWRTElyfvZHGAwWm6FPLFENsv6+omEJivw4Biz0nO2
AJIafA8g1XQ6DEl685/XdeoqQ8vyU1OFaw+GJBYYC5k/kV4npb6molik+d69
89xDmbDR+twGVEkzeEeWXN/tr8SJa+gmKZnQfLbsLnee/ed5uAUun1A/A2V8
dTt2PEZRMCefbAWobmMbqV+w8aYaK3qMYeqvBJVWq0Ct1kUGs4WGZBV56+Yt
gZ4ICi+9PboBt3gseK97CN51i73Ogoj9HoTp+AZxBKc7j+H9BvbsJzSHgL3l
vLKKfX3rm8SPTRk30CJMxYtNiZssJf9TqP+oSxgwhkxiVmEP1vEuz4DBv8Mz
t0wJTKVYoi0ZbMSF+JNryInaqFmA3mQMuKM/8+qxHQhCPn3Ojluv4QCQqj/p
2gVvE1KxXLzX2+2lBAYZRBHXD2fEuTkvQeQxkSRO9IlOFLpyUZ4s9JP7BQDD
/+ip4VDTBj5x6Ri8z23BYNb7adEM5tGZO+KLpW/IV1hv0XaeCq6lK7Zje1Yk
ZGrjAitSuJbfTOee/BHAnaSpJbIvTYkwnXdbi7m16HWHQ0paeX6nf2xW+29z
fi8okSI4vH9UnvVctBlv3Zl9l4buMlCvQPTBUHJvMcumXmuLKC3+A1504Vy3
6JGlpVerpAk+3g7872TlayGr6RojULCsZufy4+t+MBiKnMnDHDS7J7D0VCdu
vcx/JHLg5058RUTG67revUoAomm5PSxrctmmlYoyF9aFK3csZcBA8L8/CVCH
2nPEn4UyGpQ8quA0DS5/RidPImvECzux+bapEFuw3rTidBXB3ADhTPnVlU5z
EvV/iy8/9y9FxftS9uLeM0WQJ//s1hoK+KzSm8tVwaoROthaQ1cuNZnbSICA
KJY7gl+O12fYx0odKB4Sy9NYcdCl2e2lwiD1KcD9vSIYc5uUd9eH9L/P3FMV
HFsO2cil+xopETI2n6KuaHYTY0rdTqh4pqVIcIlGa9+hekUWaZP59Oxk0/Pw
yeoxNSDlP0zU9hTtmS63/2BrfY844aKHIvvlK9u6LOLAjZig6r8fpvjnXoEB
f2zOzW/DajjrOuQaco2ltzkWPyFrcdKRMsv8V3NM2LW4EPpDpqk5uy9XvmpD
nL9Ow2E+Y7RjuyxymvpRHF2gSJr8r4VHBl6diclLj/s3WHE08M+UpNfQ/ymk
+4s1SA+Zd6/Ayo9WiYyTOdb3bG6U98OKfw1gfWria64PSa72zXXyWuZwfAem
QvFdd7oxYkhMgEHJ6lsx8UtVsfVspEN6OlpEWC+X9YIA3SwjsCsXqqWCmJDv
U+bVyhqGADQnACaygMih4nWJkqu0AlgjKUtsXeobZ06ZgBI3fUS+/fQ6WnsI
2V1UCkK8pXDR+hYuGxfLzKpbgD3NEKYKYWGEjW3PzSywhK5272NST2yMr3hE
Sx/Tu6VUn1dRFuusg6Gkai6ukqgbn1n0iz9ALY91mnAAN8zBNBxtu6ylO3L2
4M8ZclFhizAfEPKUtvsymvtO7e6pe3c66oWgz7LieXl2Fv/7T9njmnx17iJa
WEE0BGiWslgh1LEzGdo1WmMauprOeAC0FMgHBe691ArLuOIxnFz257ST+RcA
V9QZdKDbhHm2e/Kfq5CXFd9S8ZMhSGGo7k4RskmMu9pHppD9LJ1eX1uKNqz3
W5n2pp6w7LEMfHv+o9GSJ6l7O7pfmAYmtpdHxAf/4H2rjC7Dt57Sw3Ar0LEC
rxROhiWn4oGvNysJbxcMvOtr8OcEO9RFmAQQqbsgL8Tivdy7fhrKkbQG//4R
Sxy8zC9aCrwDjD1bcujMKEfcrJSFUZBSZwRvdC8yREjZxYv0byAK+EAZQdmP
16xK/o/npN2X8A6pvEutYJyQrE1SjK66pGQxBBJPbBFRUAaIOW4KcKDRyPzr
j1UoDq+j3sDowt4uvpYkDXb4aMV3+3yGWCikEoX6CAZRrh9jPp9FQjHJlw+N
5BrIrwwL80v3vrHSRCzQXQIPFkjxHuLdJsQ94gQa59m4lYeacKidIhw00Ggq
TSuvNMne6C3aT1ScQAlzwwpkDdzqYdWsxJx3SwzFDPfJr1Be6PknBafyX+9D
1sTzoW10luGwOowWWAiH0d0v7sBV7D1X8y+fDIOPzHlo12CkatqlM5UO2IXv
gjuWOm+IzzDT6jlPBSq+lqqNhxqTmt0ir6sZixw98+49P1kpp9JgNuuCx/Gu
M9aNhHVLhqjXx2DkpRhvzcStl3IOkoLRBrZ0Xa3PyexFkXY3qa3hMWT2MuPD
AxiXfYAL0KgN5wSfbuVFX3q892gEZbkBzCdrM/iRgt+SZqYIc/sQRGdq3RFL
jtvYgdTebNqnqmnam+yuiVXU7963rXC2taw9MGZ/MbOXWbpLZ+WpmbbVFMHp
/35kFIA6N5wri1OQdjSIE/bwXBme+Izz5x1KjQwG3dGIeO4y27F7rfx1iRNl
4G+bSgxhK8dIK2MRp7KgEuUALAMP8MX2/WKdQ+6bUBHPto9bXwU14eFqZhrn
kMS21sSn5OQ312hEqCI1+oLPGikeKUnNbclSC3/DNLl226OVvkkh/A9FlFKa
rWH7Z7GXnOaEzLNS71Ufda06i+LwhPuO54DKElSBGZECH2H0ASox3ApCLM2f
vnSBkGtd+SLyMk0WDFaWGrRHvFv+5AdMsIExuUkSQg/ZwZVCMzse15QeZvPh
QIxTTRlBPwNxFl+isGg3Osa5LpEpaq84Z7c7NKW1ORQJe/dzIi48uRRxV811
7liHu0xAiWx1CPhkZsE/eEo51GvgAU/6kYkB6/UXkWLxaC7G/OZd9IxodbO9
K5Qto/tp9J516tW7bfrUsjqm9TMxiogi4mj7xp3kR8i+hAcy1HoAtufY3h+h
ucrmx5NawQut6dWk4ZXeszzdTAwHepABX6lZjGhmGIWyDDYYmPx+6aqeL9gx
LzrzzcdZbgrCijkTw4zmH/dfp2SggVw8KwuNloEi6pq6xUIUdljJWErI9ZlN
Q3q6nTD8vgitPl7m2wOwQHvrduHM7FsezszSWbZHjFCiYDNBk/J/ox9Un7y7
DJjSclG3aK6f7FFzuBRFb97jLirwq/U3xZu+WjTC02CN5T41f4XYlNCM8S2J
vHCmaUJdayeRJNuPnMZz1XrFZzSFuIMm0blxe06OQB5SXma+XJ+1x+XuLz9E
tF2S2LpzslQz5xWVyAqrhEGVqKaMVggcmYEE/azOHui9LV69cScIe5b+1EqA
U2nIfV7P0JTGyV5oeed9/t2c4pHyGNWCwByhsMXknr6JaBAqhL5sEIlGlfPT
CTxTgkgENwFxKaC4gHmy12aAz/aZAgP0T8kfAQu6fT4wDVWNwDuk2JSjh26u
pv4DWOvyBn8QuLSxVts53dbtz0D6j+rK5RT61ELCR2MFSBH+GQR+olaMZXF4
v6mU6WGXvdMWslZlLz11+aVr/RBHLpStJbB3kY3a5V3ZU2PhsM4uLTMfmBH6
4lRlj31Cz+0VAKq4eB37EbDDZrv3h12OY4TIIHAz4WZTJJzSIq2MmwVt604z
Pq1uSTtmpgSi2rVFDm37kUpBqwNl3fleykp0pBT1Wou80LqQykrtLbLRxy/1
nhA2jPlWcxoY+8SU9IANyl+et5stwv0cgO0OwVbO+nbnGQHxSMvzLui7C+LZ
QBnBDujQrwq+tz2zPmsb6i+okHDo1NVe27jjO39ayxP3nobroHh3iABCJlzW
Dnv1w5Oa2jXAvcuitIHAsHB2XLXi53V3PH7gVcNFQ/Vqa/4KM1v1OjWmxOKs
Le4bj2vLMq57K4+2cr08XsPoC1YLXsyya333ch7wTCksGDRozFs+WkncFgVt
0mOkP9blnP7h1Nijg5CVqqQYRSeJ9tIS4lzzIMIpLmRxUbCbeM1rYHtbvHc9
d1yl4wUaYz95SWNhWN83y2ZKGMTGqrQnW7G6SUwAtBBa4rydD4pvIDFfQGRC
DXf0Yu8JbM5tUdVJ2DfoIYyKl7YNU4l1pukSg540yT95HKpHEAndjtaSYufT
PZbodOYVN2vqlzPL/FplunX9gZerYuWcVepFrjMEgjh9QijT+bjrXkRsfDWS
2BDlIU8VgpdFJ469mBHmatdCY9T0cjsCTacL8RANVJwQJZURPvY8XBIgSz/Y
QHVfJCBZ5f6+7svnoRbRgNj0bouD8aHVNsIADE/v4W62gNxne5JxQ+B4uFZ5
jhh9syVJIlsV5KS4YcMTDT2feOm2yUwpcZTD9NXNMwfca6duD8pBU9shdHEL
sEkK03N8MPIMR2tZje+t/xNJiyb/fHNZ165OoDLqaDn4bfmY5fFQNC/ygZCh
sre/ZOYUns2x616EZ6rEmO73JO8UZX0ikfvQ44796oKdA7+3d7rfgfNwt/Of
POCSu0svwjN2/8q0D65Z13A89dG0xnyImazV8ZAYvhQBagcu+qfLmaKsxOlq
+T8Cuiqr+lK14rODYeRt4HuecVZobxWkznz1DR66euFGcBo+J9Ecn+AuHao0
oiQoLNo8FcnVuqs6a6uQPjElWwxINExk8xre5uDtBgCrn64avPMN8Q4uRo84
0RHi1P8M7enGMmjeNJRMvKYvAjerPQYRak6zqC3ZY9PsdS9n/5fChBLTIOo5
ZZZAg67rY6u13mG1iVT0PWNUX23z9LMlUxqih7tUkpakbEIK/bqXakkLLDBD
DaMBQ8RME+ZC98Y7xcqketfMvxaveqyizm+Q+pz+2uNpcNxy1yPd4AkVTO7r
xY72Kn91lnt2fgNWqxwxkYfhQ5JDvtxhAsTzk9VTB3mzS2TVnvfUPwaG1m7z
61UEnTXJ8HWZr39nsqd3N2mfBDCBR5Pp2JKYBawgv7jOpsSPyYWexLcKUWG1
DabjfgqbDBTDWs9r5n8ntTrdxrLKfsPQ8NYyKp/QZPt6LxXiXH94ZyTWnAwN
DX9BYUZbv6vhGqLFhJpLu89Ew+hxkZYqvhGM9TTvRAS3D2kzk5K1E/pgqMGw
dszTlNoUOZl4Q0CDQCfedoa9fVR0MMoKiy4INbzMZqZKlgS9cIqo7uSRHAMr
BJr3c89x0V32LtyM3PAsZD+Q7zlIy/UoFCiDa4/FLGH/qLSCIeisVMfLagio
Gfu8G349A/0OUZRowpyi7Yde9gavDSWtRbjWK2PRNXHawN0X7OpEouhmfrqD
n4w5obBnNSrf++E0Dtj5jY8R8RgET7JRVgv/7pjXHtKNCPOU3GvLJ2l8S9M6
mNl9PThvu5Q97MYQ7505X8A4pxfF+psKteoNgwsEx7Pz/9aPyIuYffk6MLem
POcp/oKO/Jx7yCnuu8six1h1do4D+srNf2cC65hNEFzpSYQP83D7IPTDSOR5
JXcQ3bCPi3GwVGal7jO44uzmG8WaC5CDg96UziaqKBKl8+ePo1XuwZq0vywl
x3rtXV9BhphIeloHjUyjSYkPFz8ZPdxXlrK39ThK2MviXDtiHZH1FRdC+qlK
oc3+ugy7Gaq3kj2kQ8yub6Nh7nNi+hlLyzBCz7ikwwrXhfKOqD2NPVL5ZwSx
fZS9DGYGt5NU/SV9lES7uzl982Snkg/FnuXg3O3l+AbftzlQC7YMe3s6MF2D
gGRYI5e093CIRDAjqRr/buBl7QkJbpxzhEnE+AnsgB4p01pa/wO8i91sDqu1
uw2mdN6+yqSUCJt6UttJT8V4fsEROkdiGeT6ffJfLoPO5PD/Llhi10/uSTN+
tIGkloFyT4FOteXdSoJN//vVdyEiE2V9W3zCOAenFAkupmRy9oo+uuBgdBoB
LpKmieRNIaz+mWuiMUhiUsR3E8WfJa+sTjTGWyPtRl+BN3sFHHIkgusdX2i7
xM9KnmFjCfpley1ng5o1DUuri68gBMdIE7Z1FdFbPIeOQFUOvUfGHMoSPHxg
ySFtga5R3dXZfhXAs6L40/UcoR3sK8utAvyDoXaOga5Qo8xbNC3+rncRrqLI
vwAm1qqMNvjW3CrUn3FtDxW+RomJxEv6rb0VRmHCdBYy0uNbEpTw5aPYW31f
Tr1j7w7kXmCpb+nRXwGai3SivJ3iXAu8QWAP6SXBtJ1lVnnXcyX6GrQCAYAX
StK40omn4/mh9JiwM1SVJBJv+hULkJqfXkwW84FXFNQB+FJlCbZno9uBoBtC
cLjZB+94T2EO66D6r7dQIvW5ZDLE03EnS0entqg8bJ6Dfte/FPwATkKsBeI3
Ge1uKrhHh6MrxDhNomI1eei1Ybri0fKBOq2fN45zU+oaOm0qlAhWbUAs3Ylf
8jrARAxyadVumAK65x4QkU7mN8+/hCDxnDRr1qxCVJ7A/tQiF0iXU6EbgXfD
RitYPjbzpUB8vWpCB+bJSGF9pdaeQ7qI+LwOJQfS2Qy/PP8WYsvIK8mjdHEa
cXBidgKKh++tlsp3yLLqNd9wQ+RXj9ehHrWxNV1WJHo3gCnRIs/nsjH7eC/I
A04q/ZrPznODIAglu6qTihp7/4q4IbXJsKwMwr23iZEbrGCkg58AY/dOnWpe
LdPM456jiSm9UPKf6ySKGmDBJZazCVQymIr6tbZ/CuZWXf7603REsl/Ok6H6
DKvJYakOK5vxkEgGLR401j/XYezM0P7PMfWKSSB//ftuhufXRnQinPTACPnM
ZDPtLhDqsjfqqFpQ5T0FQoBrSeSBES2IWECGp0dp5LxxLmpDLnN5KiEmlEp3
cthpfXIBFFfgFqqRiuYKhJ4+1m3MZ6iKjyxTf6u5Wajo/tG9cdM8ZzCOevmL
IjoUJYcWLWvpIfUVOx7FlpqRVFBNLsY6BHCLtiag4FGvx84ifSRqIA0aVWlu
TEH0D0MEyZ8bSG+ihWObENLhZ2RGI+N9wdDJzLZa88ipOBJDekNFxRbewVs6
ythbXj33yT0H8daQ5680VJoTWf4irfU/bYJ/sruU4nD1+rWs1sQtgefdK8uT
lzq3zOElF9HoYaReK94FbeYjJxvOlMeLIYW0DyqOJgZCt0C96tiQeo5nVJ9U
xoJzUt2030BjAkaMCr0TPfyRVEgoEsE5vftQOt/Z2zakDh8zsPx6m74TO5/G
f3phYorLuEOrwb2XmBtIGFzj6wlweDyzQSuVaG6FkoDUbUEIuLF/cUefDlD9
MVEmUmTeWP2R7p2uPoK1NRIt1ujymly4Ga6+FK1OsRYcyah5QXChmy86mT+T
F+ZV5N6skjMUyAreSQSnwuWisEcdJziOqjnaMmwBvoeo15Woboil5vwh5R2V
dA2OFGHGTJzj37sEK+fWiAtM6U+to5spQJA8Ykf98k4j/x+Pd1HyYUFlRa27
Vr2RUeaa3VGz0nMpvHEJtjmk/JWYQ+MckE7gCWxmXDrrgs3Nr4JDetZM4pgP
ycL0AIkgK+i1KR1Uebea4iC0aXi1Kt+Q/Z47lQoJy3Kt+3QK2NA+NDrym5Kr
H0Yq9rxzX7dijubvtSevaF2RsL0m5JK4Nslro8G1GG55HN1oRSnE1D6U7H3D
88STmhZc0uRnfHEkwWGBIIj9s6QQbm580jwPPKsG1TOs/xive9rmSOdh+JZL
crLkxnJwsJ/m9EIsm2Y/Cdq/8zjkF/hr3d7wWqS4Epi3dcZK4IZ1yezvE2k7
gFRx6zUuY+eeMfVYTtnEUK+NFM7znuNBJT580/KiWE+yUdRBBjSNIY3VqeCQ
VwrkR11iQCJ9biFaGQpQnC1tWNmpiaKz8RB6ce1NLonbJ1dKWO9JR0FNxZyO
qly91EuXHdo23kPl214NG6ozNIdXXQnUV0WVjc2dCC3rNAxYXarwzm6HcSjj
N/yWDUsf3zT6nCQkfDoG4gbbp4MiT1oImMIrV4eEYC6lqhucoE9anxbJhqMn
K48Udsk+vCHPt5AKhKB5Kv7fjTG8Hfkd4bR1/0LdQOnI03IYMRPyV8/SBgVL
dVYP2XCPSs4B2/I141yEyRbLq+EKQ7O/wamT2XnqmAo9167u+K+otj4MNcNy
sH2THz6ELAPzvkb8IAqe0coYrG9TJ+CphBZ4NRR1mo1ExXGNbV1QnLbTwoap
P+FetJv7iUMIMfdvB42j0Hv8U3ovPZFGNa0yjqPqWKABxxY1kZ2TI0LXbMVO
DEVZZzleQ+vtlW7EL48Nr6klXEuHgoUP+1dzrYiQwnx5tJzGfwlvB3GAN3oo
aQUNXxF7550B+QMRSwQd+Zd4eU8qDwEmbR7J38SR1yC5utZKbC4Qtlojwt6h
vgdhHj/bNW1Y6wO6bmEpcipuq71dodVwKkNZwvfRdWZ/ZT0DebhfoDmtdcwo
+KQWbk2BBQTigoaPgOoXkADJ7xfh9GAlmMqPMj9oFQuScgVypXYd66CYBRDn
OQ7RwK/lJ8jtKWW354Xyfqpn7vNA1DLBJHoYbqdvDc854IfDbBci5DN9n1u6
7OgLcRccHE4vNwQ36t6O5l3eSB6S3ylqaZCyirDQfHO62Gr4yMXYu+7HWTVI
l4qt8lLSn6IgAek9yNAf8KnDRsoR9Vuw5gTeoBtixXAzyMGqdJsz7AgEze7i
l3gSFGksqXoKRw92hY7+8iOOJJRRQPIiyzmw8jJ9lwoZg9e4zLFzKbfthYgX
/49i9qZsRcKcNAuPJMdvDOVtDKjqxbc9GSOLmlfBhCIfmIkI/mY0gWpjWRk2
KoWsd6kH5DS/Wp/7QCF407sR70CihKLpJ1zSW6Sh5hx8ZsAn50F+7+IUPQdX
A5p4vl0w4B/+9rpRySjTQbpWOrSxYSX8uiUyLRupjOXmpVoc8HL1DuTBo5GE
GUPRe6Cokn7jasF9gohGvMMsyLRQAKOc+kOYNiS+LIwP0H3CwVWyxYhZDY7Q
klNJPehG89xz1V7NaYTyBXxCmFjnwHS9i8gCiMHguBrD486vVZtkn46R5BuD
IGb2+RslHUpiKRSCa38KgBzECr7BIeuhVxF3swIpRzXEKKGFvjMgq8EV1YGF
lcZ0PM25hCNTuKbI3If79zyGrmhnXv3O0JMR01ohwtSOeMVR4yv4/DKc8ue2
isOWFRfkJyRXnEwGBt/ZR+EBKscrr8LZQRe4EBzEZiy2cu04SkZXk+7j4l1D
WuBjGPiDXZLzATVX/Z0EaNerPdi0ouUE64swQngF2VAauJv0kCD4xuNCppkH
asSRetGCv086pWtRWbRqle2TGxzrXLTNLlBXQrsIUNZkd3uxevdzieUq4uS0
jz6jFJinREQ6itlhSC5eR1hTL23KP0JWn5TNJ14E/mRpG7gwi9BdTBn2OCQ1
763446NtfHQlQaWYFI8P15OI5S2TQkgw0L53j65dFDmbYv3I+2TiAaL2hC9W
p0mQhs4hU6NaiEbLw94ISFmXBV/NKdaJm+fhKEsbDy/MBs8TaVVim2etYEGZ
hTzvpp0SFQN4TMtIT3e1erb1uKhj7ZfxXnnOCMzwnf8kWF6jBhz6zvJIPi0l
LX5ofvamSBoMrQ+NDL2ikr2dNAE5ZHltpRl3f+jJ++fAPQHjtUMyBMCRQgQf
eZ4hb1qCIGegPsmRo3sXa2ISezeOkcw9+ubWoXz3IqvlVhQWfLG0VbLOaVox
yGaGh27iOZlA99Iv37VAl5R6DMkWkb2poChCbblXx60k+ylTnH9/yY7Oayh/
9rimpB3tWfcM2Ct3ZIkSSQcQDBJO0BDwNqSHRc1Uei4ncyWaBARz4xKx/JZC
uye6DNfnM+wwDSvl4Gx/sJW/cXaVgdR00F3Z4qhIbg7+wxHjb4pM2JlHaZNc
pA0hM0kIHzFGm7TT/xHug/2Y0yQof/anY8TVt0Kb4Q4+BvDDEScpCRDbQJSf
Ny4MaJ+wyTgeKOgqjRvFjU4CAAwyhanmdo9VVyYad9vRB+3rMiWZNVGUcT0x
inTYXIgQg5Fn8FCDzEHwow69LcisxJdjuV1PEU29JZyqI5cxNnjTnIyjl+yI
PrBYP9L3LwlO4IIESl5gQqez0p4UwhWaO0cXcBqDQNkAzWS0z5BTHN9Xq1On
3NhsyA+bpNVs4d/bO+KusdtL59eV6OB2MVWV00UeSf5mWw01WE984s6lT+Dw
K64B517aT3fUtpJLEpsQAybwwlga8CyoCFKz3wWuytbvBD403X3ib8hqEbYZ
pKFDg/iN27wb29FAUV1FYf+IKEeesfklHl+6Q/DFMZ3JbkoXtjibX7xuhO8R
EfZqktzlGqOICjRZ18m1JXCV+0XHydRk0686yDyyakhawv/qDMgPvxRzPbqw
xKxoE2NGnTKYiNwR4IBDDi6p+BoOT75B91wiTudL/K0gWzRN0UgnYOR8HGDM
vWw4GJHhqF4ldUH7sHVFfNuoQWy6WOanw1cesALTBwJnAXPxZaS7fQ83N3EY
Bqu5KySIEAQilCo2qu+eMr1A5Ca36SrYBy25LAtD9Up5QEl/yysTnf/KOHjw
d8IK9x5u06DwEDGxHh/X0m30b64cWuzt3KFSqZgDgKhcDdVDgjykJsJErNlh
RbA/0AAzwLugsLizXbqoGFRMF23gs321nO1RVR4VzvAvvdevAxiJJ98hsHvD
r04N+yB8TrNTX0K8HOezzJp6pRLTO+b68PC2hBOW+Vxex+qMPx2U80jE6pBR
Do1G+xA0F9yETrKlCuhc+WQwSH6l4++8C8uOpnkg1EXAiCxVCs1KJWyh5M2L
wYeaZ++3dj0r17GpU1+KZASd+WCTE9iPX6vGATC4hjkKqX0kprJzh86ilSUJ
urPZH1efsJIHzPDeqX9wWJbyOtnS5oFkvtRXt3mc2s9rhyWEhn8NzWxYnxE3
qjaLdhk0rYfdBP0AY9hEEEIH70sZBwJcsQCb/kQRwTBPhGjrT3cT3WJ6/Qv3
8wNTjXbsWkrj6zR0+k6Yuzwg6AS5R/CpQG4ZpMVxXWYqkZcDOgTNYWItQG8C
HpOtDQZfwurSemq4c9q0LBrXNjMyFBP2+DxhjgKRTLd/hgE+7ii3RUyQaVGC
kGUZzHs1GDd2Z6UEuoGNkNQOfu2YxwyNm4Xk4iQmsrLXxutTZi55eDWQGDGl
4kaRmlnJYnmgycaTQMZo9/ARUcH/4Eev4swQnydIMoKGVdWrO0u1Rsg1VXik
4pklxvDpYcvyaWJme2z5y6+xURGWFwDMT8oYSqywafMlWeaDvbfUaklC8L3b
ToPUzDL3x5WG3SlVPi+zmJwUgULJO1g2bxC6R+BkSk+UjeUJM4XI+rF7t7km
33u9sBrTAziPgFGWhLaa8AzcPTlokOY+Tmr8zoTTgmqJ5AHqjDWQfluOGH58
erKFScjyMW15n9VgrhkvuNHeUvIxHjwj/BXjH/KnOW/vupczsKGxm3IVaHbg
h3Bl75FUm4UF6eeumfl78/07lh+BZL7AgHpZy6GjQBKyFAVqbc9K9TF52h4M
0Y30nngFnznP87Jx3vZn3eCYnOFFtVevf8OKnupAb6iqw54+mY+IqCBTTspm
wKC6fsqB7Q36X70TuJ8KgWZLK7rcpppZOKH3Tv5MmrD3cEaZzTqT/Isy1Wxv
PM/QoHh7uSD9DdTO6m7XEaafaDKhlXdTz9Gu9b3vasDHqoRERNErtbd6DZLS
DkSOl/FK/pxowSKN50uIWiBw0Ehy07lWLjvUfMRtW4uUmSTFNrARFLcInhCf
BAF0AsbuczNt1fbo8wm85leLgSCyZmyl8w5+F8yKAMFCCRlVQckvWwq9PW2p
hH+jrwxOcSWbSOu2AhoN9JN3cT/8UFY4Daqu7Fn6mSyNhKK+KlViRxjNtR2H
B3DFz/Qs/kPnRgOU6VmgwvMnepAT5qwgxqHvL2qdxQX3R29+RiI3V6so7ucj
owFqqisl3hEu2zyPMZr87zlcubi0RbesTpeAO25eptmDv6l0eux8ELyN0drR
9XaKBlCD9JOf9wi5LbM0hxiM480peJxBX6j3NdZh6aPELDjKb0K0Essi/6de
1z+qwCkd/+mlA85bJ57mdDDs4iWu2Lj8xuT4m+VT1wRyscfNI4WoIc49EJy7
N3pdsrv8YSl4OYF96sH1sEEwLBUhYW0IPXbNgtrlJNpVWGGcSjPJTvGs76+X
/Av1AnhS2xw5eM060u97pCaJbc6lk58mlfp5nHGCYMUFIEWhYrU2LJj4sWd+
9UZMc+snCAO9oj8lc9lW5/+VL2/30arwfL3mVTMEs2rPcm8coUWWkTHHgGgw
Vgp4bNrwU+PdHcyTF9JPKYHimxnpHv9qajzsvyWL4VSKm+JMPlJ/tW5AwR36
gD3Rvl/QzsifljKcGAvmqkvHOd6CRbLWSVCqBs1AoGt0ZdBxyvy23hfPNlcT
qAVhcLPrrgyoAJ9XgPLflgdrSDUipuJBhIouwT/sw8s8NRGof08zq837hMVa
Dyu5wYTMhgG5HzV+11nKF+ejzTUVbiXh5ehb7kzZ+Is3lHjNkigY66dG+Cli
RTLWMkfKZxhnDxI9IosPyIKygToaNuYztgcduJsjXZEWMHrHGStgGyE40Rn0
IjSl/RvMWyAcfovLW+x2T1CO2EM3uyt9AYLk/Mdzz8C92OS3nnRAPCQOCKrV
yz68BOuQeNZGElwCYWdM7GGZT60P6m1kMOQRhln+p6qqz9igLz406OFxVanF
Oae4TndaII4RXX7TbnzZXy2OX/wEt+UBBADtLbK5/VlbdYL2xaryw2pXbkPg
htAv8KEGAVB7WtfUInbmU5Kb+t746cr75Mku9P04OQsrHStTqR9EkdhlQ0Tk
UuEFRHa+AGo/vAmpn+rWLOqdhJ6YC9trKUm4GKKodb969PtIrbquLJm+M8Qg
6VY8cGAc/wVBM9My1HbGb4/rknFskMsiKzgDiLnb3PirfnK032Hssyd696YI
8sx+BKvzaLxKYMXD5+093LyG3lYjxNlQnqixjlgLdiH5MipMqGvySKB2iTY7
KHEel2Gv+++JnA8PbExP+0xxkISh7BHRC0vHbSzKBYxBaYhStivUFTUInyES
COy9vOg+sFSndyvJsquCBMyz05NvqDUNIujnnngdXcKPZYyuSXg3xa68qvED
xDDWcNxcG6SWg68prn3GlpnT/q72PbwvdNRnRS+hqDHUbLWdWQ/YnYv1cAyu
JUeNwyX58KWTYZfXJusToC1yfc5aAChm8phO3snUdkQIahP8YekhfupyuQ/Z
DolziXK+14Nk8Ao8pu9ACRiUVMOcPGXQAqsCgqPHd79KSJ67qM4ozyoKsz2O
8WYXOv90ZihL6+XdZCNokOXe8EC0wZa3hT0JPRJ6Whe8tIpBYeAJbwjye3f9
HLUPHqyRaVa4jmr+FX/tNANa0xcBiVenCXijapT6oYOr6N/7/v1WUfTA38//
q93/tCV9w7ovZlSBzfmhUNItZmtLdb3mcpjATd7Yy35xpZFSQF4jMHJJagBi
xBHR5hm9yx7AETY9TYFBjT2wXPLrSLbakQYlExJ5nd4H2LE/iKjlphEKD1/j
jCpCnBG+TXy+7iTkuIk+kNBQh6SnrY60IXa7EEVVrI003Q0RD1u7dGqFAIes
EEgPKYkmnd+4d27oT28rcjJWsAh/i6hIev5uTNOPBOnrDWy6McgnKIF9PgRt
/9ZMO4K6aalU4E7ddDwYK8H364Rr7g9AlpyoUWtC8ZhJyuZStoL453KMvbpG
vc/7m8wrLGv2QlHCzX7MK17pW8TKRWIwUTRnUvQnj2AlRmzi1MUXZ5DnJ2kZ
maYicmdvG28ZsBtaGdM9S9RTCoxtjcFqHeAJZX7EmCA3PGbHMbjBxDw6T0fJ
OJOdWIglGgnOSTPya63hhpwl+kEBVs19ZMSP8cBYhWI4Z4PHMImWze65bSvj
WTPU4VVdlWOu6oinyVbIbdwhZJFjEU9jtSgM8ndNwgL3XWFKUacgX32l0Y7k
7gzDE2My56v6fYKTCKKY41Sa3Pb3RuPZMrgTiKXG/RWxi/C9EzBSYeNKgbLZ
h/qi8EIZusACRyfWZleHwWcbSU2oOMAspjPDNg8Hy39l8q0k73+EujQFmcn1
sui+Zb/nBJSneCTi1Tst4wJwUpwdhwl0ek0Y0qoKN6Sow79W0R9Vtmx4hyax
bjW3LfnLBwYYDwFQC7zb8/lF5N3dxHKDvuo6/68WT9rFpFFNnzLfd7dZXygn
25ci7JZIfjnKQCh+L2UvZX1JBvI+HgeflWgHKukKP33Gq6PBtkazj6wiL4BZ
dKnhI+2man7RBscmxDEeqWPmIMYfuYl+l4PfmqK94jmh0gGdp8+3Fxj4EFvr
Ww+5exqfKQO49QUuvS9P2BbkT5zDWvuh97BZeqKAKkE9Diiv4+3Fe++ioMli
NpyH20Tbj+hvOD52xnILL/wn1lZdBQrS2A/IKd7BwoEOxXlwC/gTkzGu0nLe
/U1XAzPxqlywwPx89zitjD5qCMEf1/yZ9miGs+ArtZMNyr586WosRiqUfJKA
2ErLjiMm8A0ZVhmZ5OpVnGRD38BxBEja7a979SJ6RGZro/tttFYYxkOJ/V9g
PfBTjcrF0aiTj+7fEFkdWjr8M6u/qgAJnfHss7yRCiRrwyN1M8rYwTRy2a8X
oK/SQwoDBWS2TVcgP5iEkO1TThNNO0OI8bQw7Ko+a0i+FR82TDboqM9eggjL
3ZqQFZFuOB4GEa3hxumXmJHJGv59Q2S22HToWiVA0d7zXOswVejxP6bOPKos
KCo/06zRUhUBHDPh6T5JiJEGCVzkyAo4JTj6ChDF6XmXcIp4b1V+D2j96HpZ
GEc10+hmuug8uKew3jel+EoooUuCE8Tf0YCUdvJ9yYegG1DGP5yx1zX4+dtA
QSwOtl6cGQkJTn+3tlpeLs25LDU2QLI5TKt2EZ1uDwAMfxi6JS0RZc8Pk7S7
smJ3W2Hvjh61MWgSO4zIPVyWSAbMAaYzaJS4dS6PRsQ2Q2LRbUsXrTCNPo/X
LpByozS8RJ9VgxpxO4b5o+Wg4mJ9X93a94H5w2Dg2aav+wPqX3RrBJ1Me/f+
L5kM8PhMrcP4JHLPc8FwxGZ5+inbf2RQd8F4ZdTr2CgaLszLqzy7+f8xk4jO
EX30SfsVYKmzBLP753xnjEFDDsFNZL8BHzYUoGKxdXKJGultxXJ8l5wYC5Ow
FcZTLRlw3vZJUzk2XYWo2+u+Ha7B6D3BhRBE8/oZjA/JDOsSeaoODx9s+gau
+nA0vFLRZPUONo/+h85OIpWunY0hb0GFvZthXS0LLxR+u/XyNesi7XCWqVAA
uZob/w+jU7cqHljTNzu9TQzZ7xMDrp7tCeFhqIx5+qt1Or8mBZELsCx8sTV0
b2vsgJNvi8IhbwQ49F8LjIO0M1FliyNEVbkr24CHglKcABueQTcTU4tk1Heq
8Oafv1kkgnAoHBCowln9j1dK/NtOiG4nrm1vIC61fnBp2DnilsiaOAZnqxE+
f09ajm3eVPAVNlVqH+EXEgE2MEezyaZHIuA/0sn5n0q+jZLK57H+wZwlwWh9
QMGcviJ66mNkt2D4cR0lSU3nler3aAVeYLoSr8apDUBFbCNsfQWHlZ38HtE9
7enMHtzTyGRzc57728SKWDQ5LPJ2NfAT+1hdVeuPhJsyig0D09kaL77wwW5G
JsEY8EJWxfRfhmwzqbACZg5GD8OF30XGx+XYrqgahYw+doMWQCk1Doim0v6V
ypNqC0R0lP7U04xUp4iQ0a5hghQn3pIpKNiqA+fsRRfjmAKImDpU8YVzjkQY
nMsG6921hhzlermOuAu5RjFX2SxTGtMrd6NYlekHXtcV10TS4kXF1t1xiqj+
MRwMwPtU5r4TbfIkOvYIe1277gdFcOCmmHXsZgGTqdVfUThBGRrTaujjuC8D
1y31Dm5FCpnoGg/hHV0hsyHF0BGnMixokz9UsoeE+bWqnN3wVGS05tBL189L
LERwM4yTOyHW52pgPdkA5h7s+/uQqChIOdmZ4fGrMGJRFqypyRl0GiCHlxep
w0xpFe4/k8pfitgRAfQlVpsshKWYXB8WKtkmnV8xI/At1QC50fazoP8Z6hUm
suYW0Nc7vFBWUvgEVZoYUdtkIPEHr5nSlAvWPbte1Q/9Vj2t6ta5Zg1keVrx
at2oPv1z6tdWLqUXgxkUPzM2acZwL5LjGTEefAltby6wp1gNy5ACTK9kBgZn
hDVkgcSEXTaKys2W2ByeFljKPMME+A5OSilI6SEIUAV7dYzSxEA7F4HIoimn
Q0Dv7HNJlOgXycGlWGhjbj7wBJgHbpIcZQ/uYBvOrXe+/tEfQPQWI3pWZiNc
ZgEpLQKxQ7+ydLNwED7gU4MDRTBkAj3m1mbg2pChlDFR6quj4/d+g37YPtt9
E4yXAGPuf9+1XYRlBJnSwclaTZG6Fix6dtsBDcGvD9vKpkxWlNWeGHlsJVJB
WZewXahxSnvQbOHZGRgh3gtbKuIm2O25iB3uKs6KdrpsaYmCAlqpDdaUmkS3
wflH2sQ8RM9mykekz2HeiaKA6ofpB90v8HTga5RVwIOM8y+vUnuPUZrFluVG
51VUi2q7xfBGL3orzr3ag8py8pmxt5c9ONOFOvTSAZKiNudPJrsimpMGBmFF
gs2eZ3ZbOjDX0JsR/yCxFn5DwQD4ASdJHAHX6KVXOvOoM7bc/JHA9HWRWOL4
N2ZOtAke810j/AApig79pykDswkeIKYw9KxdT0WQgbD9jjwuz9/bv3/6uMUy
YL24F19PRXYhPiI1Q5YkskZwXHnSLg7r6c89jFcySMY4I5KS5Ha/M+9CXjyr
vZyswQUY/C7wZRJTnriIDw8C+0rukasBAenQ+4tfLtSTui7WkVbabwVmStOO
WNXyvuZimirSP7riLliQegcrXHZoX8xlotc4l2XyEupKUHDfX9MJ95Dq+7Ev
OV4kGKDNk0Ixj7zpWwFfSBgv4q/wWsM/D8KKR1IVbtAZ0cQoxQ9tQcOUTKMn
0F6GFWhbTbKtK2giubdwrWqUrtpndTCh2oYLy5y2PR1rPnSlHgfknT9iBclg
HTYviau9Sg0nDQmBUHfKTQirtmFX6xFRnIUzS8cCRzuhm2aILqbAxubQyChv
sUzMKQbWax21UpylAUa5kv5pU5VTt9dbliSf25xpSluNdRhGy58M+MrQMxn0
aYlO1fcN0xiuzJ9/Dfh0RlMoFPOvQseUFHME7NoyudocHwyMw4tuTHwWyyia
A8FR3Qt69pcGU6wZ9tu/vA4ItC0Ouldsp6mip6WqQfcCzv14C37c4+vnukh9
nA4n3d2MUdMUR0sRDEe+MkMb2Acw2g7A26lFqhRu3jS2BPnYnmWxKt9Pukm8
XbFxrVUDICucsdxir5tJVpsOWZqDFEddxrmncrmiZJzDPqqPv2j/QkIMktTl
SuArHYefCZYG0R6AdF0LomraUnjNRb0kou7Ql+CNdshCkkKHB9vUyyD2YvEn
LxNkbMlv4NVxSTfFKl5x7saOyqTA4nfiKWko5fWSGWQIUnGEMWK9xCnJNqb+
5CERurf8qKKOC1ndaxcPVRAy6LQFuPlEBgDIE/ZUnC2Nrfn3czqZIjsgPSrg
bFWu4Tv3LD+Na3nvdUOEB9C0orCNPSbG80cySBPDTpsvxNCa1sM8zZEjxF8k
Bz/ajqhhdbY4gOrVglORxAUE2rxXxsbVT1bsYbCDTl70o1+R1ktpdlzT2PZ+
hv5ujMbSMWc8Atju/BH+B62fMnC0yPS+MoWaru/7+eLVawz6y3C6sEEl4bNW
fy9cy2UFm6VTcGwm/mDfXIYJ78dSz8qzwM8+2zeNqpTdaa9A2zbZbN/sYkIi
7AYDL9U4bVxwEEs0skHZL9UubviHOUzOmG2F78aD53wvottgpG4oo2FRaQOe
jupV9twukAh3+kTjyeSOXHZoL3qJvXJvDO5ipO60EXmyo2+it5CqM6z6GkcD
0IaVl9SjoDwc3zII9NGHzEQLXRfTw5m6mUjP8zc0vrVqaxKClynXyUXNHs2g
0Po0ExSWHdZVVqaxmW+keh9yodBBN46f3FxR0Zb5KBWInbN31Yi3Fn/3yC0e
8Vg7H20LbtcYwstDKTG/XZpVlYXeJHMJbs+osGCNwNDBEGvdeheeqLiy0CvN
XDOyE1UAoYzD6A6j856jFWDqwEa7bp4uLQ/ilu0ASR3gJdozeXxWjflrTbXx
bE66hABTXnD5PbB/H+GyvQ5mvoSSBWfWg71kPLsCFeuWzVOSxLVhY0PfBacW
vwLkJVyIhcMJViWlDsnCuTV1kvfldhdpg/whs0VfPBguaFmZeFGM7LyMx6+I
wOWjAfejggLKcRl9NJr7/mfz+xdRAqxHmC3jW8pLmQ8Z78oFWd3SRkEKgJNk
FgiKvSnWGg/Zd+n1rZWsBbT3/wIO6oVsSBr7LAY6bnDVDh+28+Wo49J2dDmE
Wwf+dRX39ttdHKLFs/QyAWMHXSiinqL70jUtDqzCmksJGvEY+3VWFt9YbJIX
QP482AKFkaApbLGRwW7EH4qdFXdOoLTI3/tMnFvy1jJF4JBwO8Gsl0iD8/Yr
YhMOZovCKc/jZztvhd1jXM31o7sefodTlC/X0q6iWaBglu959qYo0nLSXPDC
e5vHHNA8MUYn4Or0BgVlzOcdVaGyPZWve4br8ZxqiA8ytARj3S1Okk0DVqkp
xoSf6DlR+R7CNH4peBtToQ+2oi0fSpIw8Uo8Mpvymww4M87AotOtkgsualTv
wkoZl/D51wshpfPwnnjRp9dm/BzCSz3N4fAFkmWNxAapel+7PdRlx572wLcf
yIuS4of5ZqSKUiI87uOM+DpSZ7O2AwzkLAYWfCGYzyeqy7J70TvuOkxDNJW/
RKotZNHjRB/0YcqwhYvvYYOQYiqc8pPBhNVIGk8q9GupwHl4S6wPPvZJj7mz
5LHDP8Yajy4CdmaeKOM5YbMM7i+JZ+KkB8/V5H9eBRZpcgNsLuFoZyngj6Xa
PhDX/lexr89r6u/cLhf8HcuQ1x9ywSfa707YNRF4R2UmeJET4g3Jh2osL51k
ShNxvrC+dfw+H67fsIL1XDtjat9toJqJAV4LZSbWsxK4RC9dD8EZCmeqjDuL
H908dyisGASfp/Z0A0pb0FtUMaMDh6f+FlPyfCsEvGzZH8e8SbfFYT0/fVcz
QOeVBJLFYSSxOunBENg6aphPXZNUiQ/UEkJVEY9y8HDK83snr+24iiof9eIY
ABjeJULNBsNU7nq9PTnOA8+6dEO4R+N54wQA9ANJ92YEaqMaLUQmjIUHxv/Z
vqO5xCMtT5i8yl9KCNqnFuBYmWY9txzVmWp/ua6odamcMJAbEOw+Znjqq9Xn
Y+GOThVAV3ZyjiOWZKbarmZHFF/+sldOe+C1GpUvy8JpDRdQVlarNuNRBdBh
uH4el6gWaw2Cx13IY1ztUh/1gI7iCp3VMay0sXDiHMDLNPmc6XNXVwmTQoTw
cUMINJQDRumuKpQpFTHQ1anFs7rCTBMpZBSAVikerw6cJzMiqCnR89NQw2tV
AkgKWdqHgutgktZb7LfQ8qwRJUgWIqn/QkhIgBt+GFN9Ee4YmsiwcNi3jBrH
bFm9XJui7Ijo7EmxMp94Pe7N8GcQBjvDtjroKctE4nZdh6gRkzQDFVX6orPR
ORfWftn5w/cibSuB3p821VvYAuzQODdEyRAhJk7EEUN841o6fhPOZFz+KPPg
eD3nIeD0WdXX5QiSjvlx0sfVFvyQTLFfq1Iu9ojYTfTTWnkcwweflhPyepvA
U2QD5cpH88vBFbaORUcAkSWUgCjIXSrTkp1MAKYEYbM0KDVlSfVB8ITD/stx
ihMW0GNvnxOmcR8PM5Fnybx6sZvPg3EnuJDI+NI+4Z3hik//RiXUdNOcWLWP
D1FGt4fnWkPOoHHSd2eyuR2Rp2wcJe10sRswKhn0mQbbbn1eLN3EGukvBxeO
HB/CoYHHGzEl4u4i3Ur/UdFA7y/iXOgqlENofh9FcJ6tcx0bvpaBSsGZ4md+
s6GEcFb/pofVxgpGXZoPf5WDOzIQXNjlZGpSesCmdumD8AxeUuTbIgFNkA70
dSWD/HvKlkDeWcFNav3LzJquKoaWQDrC5ugAYffwdrh2sDNgnY3XUZV4fm/S
PV5ZuMaDKKvwWds4k3D1jqsl6upLeyj0K9QvRgk3p51Irj0JfJmopa1AU5lD
xeQ109GSkKjWtU89WQWIX5PA2eg2nTk6/lGBFvJYxRjDJjKIPOUgEp0OgEVw
AWPssw4ORN1mK43YbhxAFHXxhQGl8gAbgoFWuqZzxsbJISmURYnI1JNv1ARI
vaOPSEJeI8NZ7ZPiK3jA+lT1Q5oj2w3aA8K67T6Ro9z7NJjwbdn0H156NRv1
HCzgf+/QLaBGK2fsdzGFmgqEFhiP9X2ZVihL7/lLdIZuOvBgRD3R9CsB/xCH
NhlxCyGEMUMj8MVKbVmim1oBh/PN3vhLgTXMWaj8qMjfLWnHRopWWCScWU1Y
LW2/vu3iCADQv7gjmpHxEpnXJef+vmlDHIoSnZ4c/mnPYyTcZloJN4vnDecN
WlzcrMdCki16ub5D9pjAjUftjW730q0Jyc7upGJMkSctGsS8ojK85VvE6XYv
Lsnvr1mqeQdX+vo1wjQt0awWzqLyzhFFJWcJ6ycYygRviftB6h//ucUAcakm
T4e0bGdXYrahLITi9LwbAn+Cuv/zM12OHR/mbn7b+m0UPpkwJ72jA9F7ybl1
0oCmxX/VCk5u1Sk9frLm9SSD+dJbCa8D7GeDckE6FJcNFccXrHa61QLlvx2f
XYHMwkWd7gmosz8YokBVPIO1Ae0YuCm+1mS75E7LQ5DJF35fndlO+LqNBSA4
5REUNbwV4DLwQUEFsiuasqS768AEiiiJ7riw5Y/PPJIbJCYgitz4mKEZu1F0
EnsYwbkQyY0TmHYiGxk0LAJQgKtwPXPiXR2uqg/fsjCMxFPnJGHLMLRRLpp1
FwkMxC52cW/5tmuBuqb4ZbELgd6595T68fKnCo7aD2quPg2eFYYidPdkQ5/d
HUxAWWnQdMVqxa9Jf/NQ1+emXgBLg6d7u8VxilYsfNNoEvhoaGbqIfUBQPQB
rVJk9j9nmaP3Hwf4CvXlBNj3GiGxkg3TYkxBIkoIio50A7sDv3Ydfk/8jAWc
KzLMVHVnlM0/UVHD2z8YAWWkK0gG1Lfw+RtyM8lHYus9Knr2SfViLHquxlYW
AW++aGjj3shvkP4gv6TVdOHtCmcY3zmQdYgOUxDHJktQBYAvLR6M06yxpzwq
lJ9dNnGFEeSidohjhXxiHLksOuMUZ7RR81usLeyhQ8epvM8Mj3FMH/reZN6f
NgR3SIp3Q27esHgCsq9cCznf6hpjpqNxzh1OPs+HBTkphBP/o9m7of9zNfQ8
+dJkfSR9x2+pL+jCOyU49J/OvSzd20FugY5B/kdkMkZUimL4Za3RX5QFwrtK
rzxuG8gNyI1nAuboOzMmTC2gpgLcHH2xJOM0y4Bz++eeJSKSVMo7ZcIXRGwx
67JzTtIXbwj2PhXQQYWFgii1rYCoSQaiBUjYWjH/ZrU8oTT4xaPjJ7KlGgzA
LxMEP1AMn20yoiww7/WVCfuk2Bu1HPOubCoGYSQoceiHAGDh/8R7Ejr3fGoG
DsApt2H9fYxi5UVmheA5obyKi0jzd+fMUhvnuBgApCfxA+BW5V2EsZ2c1q5w
gUuXEV8Wid1/3sd+maaWruYqTyrkHk7DBfgDSoeKzq+C0sBtka2mOG4Xfwv5
y+XQ6amWVkAZ3Jm0WW1dELFWebXOoUjAZn+fdLKxnqSoJk8i4EdHutvRv0+t
pi3G/tmXvM+DCnWhNGsZFi1SmsdcG6CpTnC+3Eg9vCQ+iPfbNpAmOsaAUm1t
QUVltqowL/bjeXNvcPVLoL603XOIfXG8pO9zMMlFyWRCOJ+HS//7ml14oANx
XQLHENQwYGPLZ+N8Tx+TLs1lqYG/F50BEJ9cndtRWVkATwyDPjGqXw4ZzvxL
67k3ZPowwWPRA11Vc0ajjYk5M5fmKGevUG8rWb/MaJgugpnhkn9ZgybXsNgJ
abzczdEMS2dWgTkoiaMPW4YygibUvFn7L8qexx1QHjFByhlxUHQgbGJLZkVx
r0TrQ4bVQxYFPjBWjHP87qcb7CEMjWhHLE8+6BA4WFNTQUrD6qatWqEJqV/y
Fng2JiFqiMWK7wbywzIlvT2Mkoxm91j3KOmPxWW2J6fMB7b6zqs4emfN5NhI
gRN2RH5C6p7TdqdNma4j1pfBs7eAzFZSj+Q8IDgiZd79Dzpn3u1YxMs4PmE9
0jy1x6CpkU0IHB+hlPgXZ+FGOx3OXKFZbzQaartenrwiOmJRSCbeCBX1oboD
d0VAlKYuiTolFYNogyssEzzPnvBmH/U48Kq2lrecbIzmAMRKhGO/+seFIeIW
3hS1hD0Q9N6+8utwkPBFO7gheL/9maVXY1mMfaLgS3c35Ow05oJfTJxPS6jL
ZvNHbD3Sh6yfvUw9ldm+P1tL9f30ulEb8RNDy8XLTZOFAtURPNWhizD7mEAU
35il0HhD3SwLU9AAr53Ya8c6Xj7JlktsWQ+BH5dEqrcY7gAc1kpYq/8vusg2
mtRWQUvEM/xxr4E2b9Xjm2nUK9nos3PzQETRHtO+HHHZ8CEAzOo3vDW40fe7
UZjvtbyLyTzUhLpRfFLa/zkdUyypNpTBCrZggfMU0r2c4EIE5xqRbsvCYPfk
2q7gT0LbJEqBAxbV728kXeasHzkflbLV2nbqw2zrI3eM4GZwYvdFOFT4Xfr6
tzHi5JqOBB7l4DtqwfNf2OmmcDgmD85lfT0+/FZOQWQCAB/tPeAxIbgTqSa9
A5HZaR2rB7p2wJ/P3wGacddth0Gddy0PS7YpHyo1iJI0B59QgiIg6moMTWG0
9MxM2q922c0O2FdIkpao7V1ZdQfrTZv71p6bacfWQAZFtwYD2Cy9Il8KWbHJ
9gXQCO/bXKcHYB6qbikHgHKsq8X8efiW3J8uHIFgTi/vtS8ykXAJa0WNdObl
rbK/W/7FachrC3DLmQGWZjkY9ptTlNlvB1WKTmzkkm3Tn2vMJtLvaEVkSZo+
u9dQBIYDU3O7bXyVDzkGnAHl0BktJj7IVIqs1klVuc3FLIsXn8+6XjOttzJz
6yjZcKUey5RAwVUkdCjx6mff3ACNWizePeG1jp4PpTDDEvhwfTA7uyceYNAZ
rOP4niV5/WC19SHy2yZu6jGFzkxbd7QH/u/aLWbTIGL1MHXiJLo5im69dJsU
7I4TaRIFyJW2VC5D1UsIZ3kZcNPiwGPBX0JwljZwuq1rELYCwUexbjqQo6Yz
nzCU2kuj0ZF/HizOYAnv71NzvRL5sJTDllowxmvbnIRWKfCxpaAVxnjuiK5K
haXBj0Y+5FGl1fbjtCTGgGEqJ5yOd2sRCHbZ0tzK00kt+/+CKabvjrvUmooI
jUn0Ixb6r0OgObJX23Cmz6/v7THEQ+jXE16FaNPhh5D1gF2Mx2VZV45tnedE
AUNg2C8UM92tjBzHWnbjzitN3Rm1PwykP/GRaJWT6E/2LIjRG6XfadcHxAhX
DaBA9fPYMib18vCO/v9otf2wy9J1GGkb18lxx77oaR4nDO9dI2l2QuzVkKsw
QGDFiG7ax3Sn7CUlAURKAy2oEDr2vLEwlyC2JWp2cKMmqakpT3PxxkJHGAg2
nTZpcgfN/4tKzV5I4nu/gvK1yUCTIOFDYwynaI2wAWNfgrs7uXUz296iHU4O
h2NvyH1z5phxyLUPqCBuuk8a4aWQ4yEKR+qSr5dhwOF95NP3YoxHkTW4eByY
P1Ny1iGoMPcVtw1CFMTaG58onkml9hxNL3yLNBi06uSv0nJz/D+CVp9N/yVp
Q3P/NOYUpdjuYf/r96HaQ101Szv/VWZ5eqCsKXyMTXR5oMSEKkjPxw7Rc4J8
5G2pYAm5kmlSO4K+PTmzi5fthClIld641kM6qpgKM9h/BO4AJ6gazbqq8LR0
BexZjeERocWr8p/NAdIqAcGn/4O6+cXGPV9tXXp9mPRSYaVsEUpFt9vhfCvH
qTQ15I7YA/EOG8yV1+kOc/SE3vuCAl+sh9Kz0EFJfYl1x6Fv3vXyPRFpniqi
0q6wwFLf/+Nuz6V1V4Nz/C5BduF3G9mPAWx5sjd28TwSAGWnngM1rcVdGNdy
jzaX6quBOhGkmUwtFW+4uXY0ApLNCB5SzlmhgGbqvm40HVbv6J6FUG1i4Ima
Cv7u8GpI4Hc247fBPOdDGKLRIifAqLhQmscvB7/pKrd/f4ILT8sJWEs9O/La
B1Yktmac3QWXu9dK08rcs22ofpu1wyJwO0kurJXjCrc1JmWf7Ba0i4fBljK+
FAS+VSTHrQjLuZtZuWpJxl/p2p6FpR0yFYa//HzjhFzvmS90MZE/c4KdlAdK
b/tjxcIIja1H1H+qhtLvKbqtSgi/q271aaGiKpLomjuV/1F2BcPvDk3v2oT5
SxNkakQZT0xGC6xM7j/XcjUkwZOeGpQsazNIRYgvQ2SSrhxQQeKAsL4vvuEY
8XOZMHxidhoZm9DWZFAGpkdyuJ57bQJdxgRocljJHl8170oAwx5MJuYyymul
9m+otdIpWV4Q7AaBMgEcchlfdr1okTWf7mjKONC/2pBEsQEfMkBjNj8zYS84
LzauL4NI7KlTKEP7WF8jQ+luYEU4F+POpdqsxFabm8ryDwRw79hdlVGrMmfz
frkZesbaZSnxwbQxNNn7bpWHhyRyY2GxHNCHi1m/lCMv8VReBmNYIRNkui22
8kZcQgadrqd9cUdaMiMdED7wVkuUemPs88Z4hNTgXzhSqnaT98nzdzwrmyjP
kubw8NQ3g0Pf97d74UEhV3rg0XOTMgSlG0I+qaMAWJm7viMLygSc+3A/RL5W
JVsrPUqxhHrM76NbxDwERA96stuiIHGZKK6mlAv0hrF602bsCPL/9x2jmPwM
yH3091ZYLHNAM2M+4rzZq5b/AHW12Tz128Kj1hBw6TsemqngZsYJmAIzQ/Ym
XoCu1FR0Axjh+awwLdtxn3T6oxElwvHnIwEX8ga5PCiqIHrN+ffTfSAyF5O3
x+VESLMm4BX8wV4LRpFhnF9UxO7qje/50YiXBFlKX4CvIj5IybaeHEbyhYnl
StqpupojcXAmpW7W2dhXA8vf5pOVRPPKLlfl3OR6s4rxuKwgJ3f8m2Wp7RWO
l+vqf4GY8qbT0S8RyjH4ufKe94R0LSZdhkMZeZGf/MkHtmqTuvpXqHMQJAEH
JakUSCLqf66RpogNcjk7fopw76fY4gbqTlP6840K+rOSS1O+mfteaRpM4ku1
PHP/0jBoUcyQ1eVBZo5z6HmN0UjwDGXkD1ONp4rkaaxcBhpn2WhnEjfwePog
S5sTRJe2tTO2dLFmdXio0vlrRkoPCQOixpXR0AmEt6ljU1GnOwCYLFFRrMKU
A7j/g4fZPDUhIF5OxIE54O6jSRK8HdaKWLKtba+7WgO8yhEHp1IXx7F7z9qO
Y5Fj/wSKQciZbkIPFofs7Ggfg4fDcontccK30Vo/OYPCCVDqbAK8r/PNQL3x
HHJVnQN4AOE57DqVUR9xw1AptcygP1ylM6TDPQkYvU/rcsdvg5sAB+5zwRHO
a55ojjBrIn1E+2VDoeKTynRo1LYRHfeQICLmVuXFD/8urEnB3iOz7UId5SUg
3L0ZmA5k0VognNlUsexXlHE5kuG7IABNX1Jn+KiwV2zMzpxpA64St4LqtU8D
/lTpMVJH6Hqr/GJrXXSghBgK8zKg3q87G5rQqLnXNq3A8lx83hjUm0lKtU59
ibZPhultXFLTAOosS+zKV6R9VAJGqAn6w8jOnWpVN3w6/vGUQPsL1Dlxz419
GN01rfDFSOEhPJ28KNihmrrKWD0GWixahXKFkzQqMzaPlnZHyt84IvesA4Jj
hlq69e7+NhVwIPUQvvhf1/Gtqmt/rJwWWZxdhyJqQa2FXpzzj3yvhmMh9I2+
E6OFbl/p+s/vgzovdQRBSD7YgXZUubpaYiYQotnv7hMTMDOLUupuG8EWNhIx
U0RSkCE1ysucw1alwzMoyGebisdhNc1UhtUmiiwhJgSZduxmNFmr16+wDRQ3
MYIJwYYkrXa7P57nCoqfchI60KswJnmgmwq4Li1Jb84EC+gCuA77El6HZ+P4
rwEy3nrbRJ+6dSBrZ0lnz18mIc+ZFMMYoOAAUmYR89weKjCaHVFqlobNb66K
PBzQ/SBGwGGOoTV43bHVp7L2CuR0rjGLnZPMs1MAg0DpK2Oy6AXnTk5fNRLy
GA7veyPxNGHfrEf2rc077F6hZH3VfCAcPN1apgNkZoAdJyO5Fp9SYWkT+H6e
YKTp9LAonQ43i4ltsK8Uo+WbwEY/J5Cj1xJkL12z32r+DakUBye2FNaFmrWy
rFLg8OwUGmR35h2Dw/sL7h02LLdjiEDYd0xTSTY6b5LbJRb9ahz+aSDBf31E
W+WHB/mFuV1AhY6nHpeKVorcqG3xLbwLinDr1TSJ1Vr58arqS7m68ysh3ERL
+aCUk68X2WP8qbq+XtRzuIjzAQrSifrpeAaXcS5g07YAVAjUoNYnlKjfGIIm
YE20QiE5C9M8IKArlFJZwFypGuxAfYhY1dM4zd6Hsg4flzjmbu579nuWMAF1
AcIIcPU96b1imghR3IS1P/82meJGESofxqx3LQagfEdsgWdiHd19hbEOEOWK
26VVLHfTu1DzXN18GE20JF3n655rEeynEVrx94U/62AgNVgYhziiW/myxNhL
gjjC++qiK/kO76Yufetukibyyzw8Hdz/rCzg4KF+0gpVwJT9NTHExzV3Yq+u
JQ0MH2w6Zh2t4QZ/C57xmgVY8uzby1lmNBNCAAl++sDwaeNAWdcb8oJsLmH0
2Nj6YOk0D1RIzGcea1G1SXf89nhdPo/yrGjRf0BojV2jANwdLYLxCz4YnZZX
zGPc8+vrRFRdrjTyemQAimL81rD79vEmzKiiVSnCa29TF3QnXo0YQ8imbUs1
Cm0gm1T2XNLpUET2Xqni1IpdylaiRHfTo9UhVOQSEbP8M2yReNJ02GUqHTAa
YKU4cm1gLhnlvIzvpFHbLTPbL0ebaoE/lEPQK16In3ccXpAgy0aHztryM8fy
3mvsvchTi/wA2outcs5d3Ts2mUWh9duRCU/PyWwxeKwdO7jqRpctOx8RVy60
55ymaVOOx65gEEXQJl1N0KSBh/c4APkVdpTF1DBvvpjHCcisd9TKP92DpNdM
ekBf6FekRuUofyBmIFh70/QyLKwdhWzvBOCHJ2tSvGXfkSyFbK0XLLbO7xf0
mIYWUi0vm2Ty/I9PkxfnMKQK4z730UuPfCPfZ448kf2NfnXEVJ9Wf2JPoj3s
E+e52a6WYr+40DfCY6oemcRA1PxiNGzwY9JQcGKxPPPMgYTYCljNTi55E/Dc
Dd4964fnrBzG6Q1nEDBidDk/svAyOXCN7nThwpGJXJUC/VOyP09r1Auonqq9
q4kcdrks5XfoUFxMFyJ4tdem7Aq0qkF8s49kHmBjWQDEmsbwU2As31aKhQU5
3VFJeI9fQ9gfcvPMpwYYRSplZapzH4vgibomWIQdWIFnBjqECDg9B9hZLmt0
k9C5HQmdk76KrNs1xoycO/Y/LhT88Y6fCP0BZUl40Z6oaykpdySJliX6RiIV
dhmHiXfJMMCb9btgJ7pdYyyn87ji5acHyxyBKhcM69U26RCmjF8hSdg+b5Qs
zuEsIgp51swg3llNaEpbGYKyGVxUnPda3ZY3OxGyO1IsMiGEf3nWPZ8Ca4XO
1o5DPN4O90Goa9xibHLpdxhONv9rah1SA9m2t5zsBxDToSUddzdEn7oLu+3B
Z9wLXdHZGUOGICKdjYPnFBQ9FS0TIGDXx9nc3rPYwPngwUEeqTgHnjRtieMM
1RVdeharz3QDK5OMtRWYpU+1Y/vGLw95sJQ4j8nDIUAgRHQiUTTAYKHpXDfQ
sakKVLucpMON/UlMxDXlXjhn9+cHniP5eYc3x6VIy0ZEDoXGWn/ZCpeazllp
wVAb+UfNTlO/aEhuZQSJRDEi4EA2O7bR7f4Ksupom3jDoir34L8I/GWSY2Yu
os2Vc9XteoebBZUx/RDCgZHfEVgrykeqi5n+Ox1eBchvMtSJRDlQapgAD71R
klpYZNpWheYhYxZhqbVlZCFDc+997NmSAU9h4MwaHjIQhuim0BjWT3h3ItLK
o5eBINRvtkj573JrgIPtQim8WhCdjEFF/+JoASDR8Osl5XyCWKFDnakOX+0G
Bn0cTD293aXyUuxeR5+NVkg3/+jHyo/6FeiUmjds5LA8VGkDfPsfZB3bB0Hg
5nLGE0pYA2CM2CrkhYMl2ERS/ihKp3tgS5J/aycIrkGONwca3gjyzaHq8yho
mA0VAQqGPMcD5ldkF3iqmUzUROVb7pXfSeIpSJvGi12w76L/H6DBKKvrIECf
UjxosQumyhHn3rqSis5bASjPsjxWdJpNsmsp9gQuJ2agdCFFty9gnG/+0QpY
Dik9LQ5HCFzBlO88fujVJp6G3vP0OW4zPsuKFv+x0wHO+kaTEyPWs3fjLUKQ
ZI7DCIhgFKzXXrkzJE39TuVStJNHHCzQe0kssCuaB4tzAUxIFDtqrXjpkIBT
Cd1mhoUBMok8KGMX2nFgrpfAIgwwmo/HaLD2IJUfHH1A8TEV7+7IF3u7v1BX
NZnd8Lx5JAch0rSOpDGng+23OYnnRzv2pdVwfnaUAbtJT6tTHxL6q5nJXDuY
kHTGuC+Zy1tDJRmmaY0i4e10twEqbufqN7dode4yDTmo1ywAi6mUtXfA5H7/
PrR7XTzMuQ2C1eTn8gMfzZh67kz3W9vImDNKMelp32NN4qoXlaen15OUBzkC
Dn9BFxWShlXJLvTbBpb7wLcI3J5qcZHb8z1FAsRDa36SuYQj1Ca3gqUh5g6w
I5NzUr9h0WBcs9dsrAzw3guipY9tKY7lTgyA3NEr/TVnfkA08Qn9grJ/0ypg
zzKlDJTtiDk3iqkRk5FU2c+FMFfda4bGfiKP2MoTYFDEVsXJWvCYlHQlHdui
iQ1wDDGyjvK8wtakSUfxh34L8WLHHge1T0m3QyHMZqG4rKBpXk90SvKJ9A+A
t0iTAW75VZMKblCL1nyr+xyl+pW7ZAUIjzlumUBm4TGR2CJ1rThpY9ejgSWR
3h5lusfEXhYhZc2j5bH2tct8OuNT/Xia6xX2nHHKqs08I9p6nexMt1VSKB/U
jWQE5vmUO53yn8XMb6xosEGoT4gQ1otafNEkAOHZN/8ZlZnOf1XRLLzU/LPS
IRBa3WCFiUFZzGC/+27RcLm8Mjqjyn0ypBE8z41i6/yPv4nVL9LaIa+4feQw
QXmg6rSmA7iVFROb+CHq0cTt0P+b/0uPHixrdStckwfC/D5EPAguRJnzi1S7
9ZeRDiQixnUsVraGntmJVx1ACOAEWFGHuN0ubh7E4HIohcFrENU4mu4opS07
zjRvXKI2YSE2j+lZX05CJepgyO5tsdzhf795HlxAI44Wx4yvlARcNO/iblAU
8j4iT0piznTXNnnPotIq4deevM2e1QUCfkkHBxAUbPXdzAqBqVoZnccWEkYw
sXe2MpQjPC5bu9vo5xQJn+gQ/mypXOTsjLVGlDdfRrJLVkHpxQ/J1ZLXNQaE
Xir4sT+aVUPXQbRK4yt4rqrzWd1VVT7LfyBnjaEDgUMVn8D/oVLrheK/cMxa
vEfhKo2Bk0gAOcN14sQFCMl7YbyVLFZK9evY+b7Um9zngRoIVv33E/Je82uY
O29Ix7fFgwRz8NhaYqwtnbj5rDUpZSk+ME1gRtFZ7vv/B3LPnHyOLyFfdOLZ
diJ+lPKnRS3H2qy8M6qvqH67MvZro4/BiUqcuZhQX0/ezlSGfe13p+ciIEKO
e6SBuOMOgNydQyZirC1pMkQwzajpPqjwonT0K3PM3lDbGVBBOU/W3TMiLPCc
FhTX6eDal+atKbaelD9DtX5ROss2CmPo77/a14amRppsryJ7qVkMoGqY1CM/
5UKyizhHdWvTX+ctyDUj6wA99sTl/sXu9gb+z0Tk2kzkRbAVbAxHcRmMChgp
rWztpRuQcpwb+LqQaKf/wAwW7vpZ2bqwxJNq+XiH8wSwKy45D1lLLr6CJVxs
s5gJ4tgQJVqCwiu3ZUgrEkLNlH+/lOjpVelH2PQk9wvU4usWrjdWIWyP1RMZ
tPsGTtr8kw6dZCli1J/SQg+0OQUH0PSO+3pG7fJuTw1HHaHDqJJ+/gPuDhMr
SeBTGsutPfCsC7W09IIi7ViIAC4RNczNe5sdNCNaOu8qBQtZtNQyZhR6C1sG
X29mgPd1sUI6s8ansKd3bziesIY6qnCT+aVm9AR+F1XpJn1sLqYLjWnw+Y3L
Vi/OBidwssrwUwgKa2ES0AKpG4DxJ2ZS9HJHqAy9dLI5pTHTNH4MGPJwuG39
KFx5euKjGNa/Z1FQ4z7LpU9n1V5hOrLCOvod4RgFFa2cIPDQpatM3I64xqEm
PPtcmPeBoJLr6nXoYgrbnwCmyC3KtliaD0wU/JwqhD/lH/2hAgSMiEjBbPEf
UeRGzMZ/SKCS+fSE89nai+RH0heO3cjDjFL4eGxG3vEdpXYV6EjdgfJc2zkI
0gvXeAcMvCswXaoqIJk2nWUzEJqnpnAZ+8NSxf687HfraCxsCDzdn/TynwIW
y7mLMmK0SPaRIpRYSjsR74vL6cnEdupkYKIHJPJ70/KHuh0YAaYz8tcE/74r
TUES47aur/LFL/J10X+yxuNnyEJnX+CmC0LEfsM0DrB4YUUdC4oye5NMDAvY
BrS19iTvlCMvmlHYX9KP1yF7p/kPWI3YcNiaAodDb/rIMyyFzaas80IV4e2F
y7pxxVDX28eLvjEhIRUH+W1B5g+MmG7bMzNAb+EZbws7Mb9GyOpq+Kxcqwjn
cCl8lIoj/l16zMkScRW26E+xCP61vjb3kkUV0dg/noXYOIJy1KfgdHU6oGOp
A/rXDfwG9Fr4aBh5kgn1jhpO6EHoQchLxPiCxW9ZbMduE2OU2W+GPbzLVAD+
61r+nRBFVHtG+U7LH37H9giVOfUpu8fbHg2qoXJzvAZkroOR7SRJ+Kwfc4Vw
bAjaKVgKXH2sl8TsGxcep8kCB4wsA2Op3Km5CK2hEdFa0ZJmi/NfLd58KHP5
dTyhQF6p2pKq7cYqRtjgFnJFLwnrwNIwTEn70uqtg+8BK0GaHll7gHygIajP
jHJ/PdX2aKcqsrPIU6s9jYIX1MJwO2skPt54smvUp9hqnvYHqOQB/pjglVZ1
hs2vAYn3CHg5CaL4S+q5iToZ252rgzqYAndkrryAUq6gvDmq07g7lnvEj+WK
lhxWgFXpZCGwNhQIJpUelQ9Y9hGKzmMb6oHi/SblaSi/XII63xS5BNmYEIu6
3L1LNWzuXZqI8eCYvUXMUYFr7ScDLihK9OZG0yzZciGA0+n3BWxiyMyc5D0s
mw6kxm5/ADrNCmMElz3xmEC1k2F93HDpiLi9h08st86Y5+KK8XDQT7LxWpK5
lIguZB2ntr7euxVql8dN4BIk3YWzDfy1BxJrtaLwIC3BTACHuAAFzWuCBfHk
83ZAYLH3pl4vZarN4T12aELR8ExGQpZtgNRQ8fVpYMKdRca2yHKD8ncb22bU
zG/74LG6nbZhw4kz10iqAlw1SKVhfjtpO+HUXhOWaGrAycEXE7yN0ZhE8XoY
Y30PVTr+K7+vMVjjB3IVHxZzOMTCxGjW/89ItNt1ZT8o7BMzzJf+7q9yV57p
q0tfxGkeG39fZWpKjC+d1AiubzjBqOpD4lfbb4wEqWvUsTzB751nwTx0gPG9
DunbdK5QNmYY2tDiEhuqpYbutt1bR9PAjeUBcJOpBvwqrn/95gkjCbtoY15u
48rY+IAk3Q4Z/bZrevy+h9gwu+IWZnUP0ShA65djxdmWZjahwqbYb8KTk9X7
AjileCjMzcBjRD/J9x4gL39N03YvBA5WdrUlmR0NfXd92jpAfVq5CZDcz3oP
ud10iSBhV1CIol9auBVJyaAH7MkACRKjKT1MpyRAkRu6MpmKlfO58CvjWACH
XnoQvvE6Neu9PHdc/V5FWZvVgwWLUrNjz1hRzyEFRsfDgLHpYSBjfmrmAals
aqAcRWqApK0gocIf/EqhgbzOGxgiYNz2eiynU34oPwJsfN2pHuaDzPQRtoD/
BYTvJjYXoirWuJ2A/lCx4WhU8jofBOu340aDJLaVUyS5WSSoa7jKXefftgvH
E6c8sNOA/mHp864zO1tXVjyb8TzPRJ7nNDG8jgVFh0+IQFUuX/YXWrGagwUw
44Kvb6PVcCewKE9Cq+wKTGNhkfxIkYku68jYkyqU8NPPef+0r7tlAmB42C58
B4MavBGF6e4RMxc8tEnx1/7b1fJZuiQGHZSmtw/n7vbLxtEjH7zFvpADxmSa
mDOn5VOmzm5ldPEXrS/M/6S2DbwY2oNzhCjTBOwShRxD0A/GH6Cm0SliHg9u
wrYUbMHWSmCplZtnMzQ+hjCUSFD6o1xguYUBwkl4DGgttFss9EkFxbFH7XUn
KDuJmSpnNZp2ZPno7+0BiORvy19VHj2EzQS6tp3FkdEk8AQgErr3xnZGhB/4
cmb/tuUzvl+P0j79fllvGampjBHvNBNN0H/yM0vhiSrljvzcsQPifnNh8god
EvGW1Iv8My+7l/nvFSgwr8Ep+cNzBlceOhBZVNVkT/P9JHkjFGjPTJ4mqYB1
AkdyTxTsSIh6JIb9veZHMxULl20Z31qD8GzGFoITn5Tc+9J+rILyGThBOnfW
wkbp00vv1np4YL/1zzyeOdIm74STIEkCOCewLC917F438jYdy25KGDU6PGI8
9egaRGsLZE28+48jJZSu8CB7Qdm8ODb72lo+cLN+y5EGgdIa/KVw9nA2DUmB
u5Urr4Gb7LLkcffxC+NktCKNQj+qS7T8DKMwsCQFxileXNZQABRj2TcqU66l
ZS1LaFCvet5wICBaj+6wjypyrA1s8lqcRwcPBXEYuf7OxO7g3dq1uV2QXIGB
wk5WBb0aA1i7Mzw2C3B5cnCuwLm6rUgkHX1j/7i/87kyPDyCVjpVr6c8w3kJ
GfMNmIhG6MroRvD8tPKCC0edzrvTkwZq3j3NVegMltE6gkAHREEvqr1n6Clu
OY8A7CPN1Tf2/XZnxppr9KtpJz5YylGfp4bvfjM4B7vJWy7bCWKRuonR3WA4
L2to8gw8Y40QB/kYZ1nTrqlct2xVL2yWCZ3gfk6hv4w9fsW19kmZTRrnXFEu
RRZvBTTyj1fHvh51UfmF8B4r1WysiHtKB4jnfxBCX+Aq//PskKjeLE9NqR9w
dmDBcq2PAMJ5Jb27I9Lj/HpPf8gnBXrcLldVGMO66OqKYl6KXtX3qEWvp/iU
ZD6L3lxIUoFZBONi1cNUSSR6sGNr/tPBcKCL5jW5gJsMOfnBA3o3RgupiCEL
fWJPehrBCY5aYLvTq8UopWIX9Slj76K7E2DOChtyhgqe8J1dcgcIaGY5qA1Y
wcIPzvrO3OfnFBXaU5eq4+ngjraTz9FmDGF8LNVe3Ny24IYhLpLtxYzKC8zi
/Ce8S/sF1BeeblJxC+gVlNrecDhc9BTVk4G+SAErPeIW3SkNosYKNIchTZOb
+UB8sfUfikJ13vON1COEjwxOlOAkWXzKQCT6Wrh7fA2PN8XR+8sHRHSnOmhX
2xHr9qwA/n7jcPhAd9+xD/SmEJsLNER5yu+EjJE8LS/u8+6qvVjGpfDrTVi+
x3RdaYYPHAKxNOKXsgdzzt13t5zZPjm4ZOXKGSAQiu7qdQ5ZlUDiJvk45gR7
9nnv4efBJ+GDe0iHc++SIjyAGUswdQe94xifpM7Bmccz3oWhVNgkme2++1Ar
ZJ/rHdbJzGlAITuS2ZaDNY+eC4tL+AhKpVXiyrWXmGDrEUa7ByGZpC/r2mEx
Uazdd4UWX3ca9EQKfWFH7SYAyL5iJwSe7dwVNFauwMnXdFfswYmTE0gTvD9k
bMvIAmp32acikTE7i6YiJiwmOlxKQyoGU5RNFP5P+7+muu7Gvw9ljhmMWqsT
P6ZBUbJ8Zf8dWIQI3QCBuQ0pruK27ETdYWeBpA66ZfIc1KuYak73qaxo/dMD
JDVH0t+qzIycZfnStRmj1AssTXOuJ8ao2paGQiIZgUQJ3vzrwL53fzbaDTb+
BxzbcIVEvwkis1I9ZLvJzaNFQ1AtTxa5Z4f07rwGFxhALhj7jUB8VD29A3/a
zijEGP4f2iXSb83PhMemPSa3OSH2M5VXMOOlJxz4H2BTTnlskuvxNZCZHWzn
z3n6qClcD43nvBTVzDxAoQ+TpQeCr0wtEKRInjcauCb0HJcNJk5YDNG2IXj6
dQeG7z0BMaQ1TNk45QiQhk1a0sqrDmSJZRF+2T9wJmJX5bJZj1la+uLgBur4
DAjuNS6fzL89tGtieNn/61jhmNSeT35tKBL5oNx+P1+cul5yQnNl0LOowf2g
zi8J/6u0TS+c6auZaZZVNVMG/0oJ8f2ZYyf7VuYZeKQxZGMIM8eujn9D/amQ
BMDRFfil32m8TiQISMEDKe2+AfmWOzHhYfwCtBhnWba6ytdCV3jm2UTTtFpO
vQauiLUQfmVf/zc7ifUESNKM7RDuYjtHpqgGzUHz8qtKm+W7MysF1QFKMzaR
A4Qzt/iV0Dheu+VL52L8VRmNltU6pH6XiPnmtaxQ6QWMNlHDtcJz1paAHea5
xuU5gONHIYOPF+LRRr4b5Ew4htLWDiSH0xWEFs7eKyPIjAs+4rRj12PHCBtn
544ZgyUJ4zzK6R6YA7JCR9c5YC/ocmB9JBHC9tpRt/YhnKipWE/Iv+n10XIP
BSMrYzHlfhZR8SBXvXxi41RmB7DVOBmIP0CdIYptf0n36DmrZPC6jFVv85eZ
zDal7u+JjopGbkvL17t9JVeBb/Hxd6j7ahPeI6vnznNX4X9Nt61VVwICvLYD
gTCJA0IFNX4RYgm2Pa4rQtyFdmey+6H9fElK7xokNLRprJbXzvfvfXU/ybSE
VKEmYmb1xEvLpiuvY1PrhtQW98E6+CYhnXHQ9wwoqp8NV2vgo6kXnwTQVxWW
1Uflrr+mH55/2AMQh3ErIxiMcu63YRuLT2YrT2rz3rgMCXOIV5gfvE+Ivowa
SxyTIrek+vcUoa45OTAx2EnmJicjZ1DsnVNPiwIoCRlOEyKk3gb6/Lg8M1qi
M96wq0uP1LB3exdwKxHLL+e1zbpZQNE8quwGOCd9RXoILiQX1TjbMjYZbLuv
39A7vNYTE8xGHzjR4QemsTMKSW+yk0HHUpNRKY8cLV9uTDZI+V1G3iKdZ4dn
o+wZNLVjHm622r2uIFPlX2mP/3Lcd++WX9rFkAOL8vlVGPrmz8K9vogP2kYz
IewLY0euEKU2NhfF0ZGobIZuAgoclgDXlkGO92kD+e7nNAoSNj/tVc+LRAFs
B9SNlXnHXeYY7VZ3SWhYlAmtJBpMF0cd8Sls4zAVNNuOg/lcezPMj0dHerkP
MekfvzzebjaFZXwSUpzZExWzzFl6l7JVV1bMIYgXCdE30SJ9cNnTWlfZRzHg
/mjoT9ZKrLSNZAjZPGqokUUwoyhN9858UhshunMElBIjJA21mk5bXEREpp+5
9p8SHErTMrVGjSDmR7/KDkfO2fy/zeSZZ0GU+NPVHrdI95/aSLl1zOYW3RKD
TUNbGWjbRpH7vh34TSxRr5CRYPzbq1dHq33g3LsUA1ce1XSulZSXqBUeJa7T
6Rzc/tokvUo8hh9Jv2pP8XWLssO1R/NztYdCb7zr0IV/UdEpurd6ze79Kyzv
Dvm9g5ke5fGEDWCz/DOIH3yxa9WDHMeqqSJjn06GL0vzThV5s6tciLsFra4w
qZQv4Xp5huM3kK9hoFFoZMszSFZ6VmTsqsRd2Nfn3e531JYsh7fBfQZBxr4g
NqOgyVR3z9c5E309xMdgj8ij6QWeeuE6LmlkDRDhEAj+cSh+VavsksJ3Xn80
ZGWB4E95fGD3ENoRcm18CARv4Bn9vzInz70arR8IMevc4WrCW16hDhhGYP4k
paGyByeWo0Zy00X4FHuI52Ga9yamIRUdPg7Ww/od46KQso6RwxhFbJ5mfZw1
rnC2xI2gPNAAwkvRRSjwNE+IjoL0vxBhrTziSYn2Oec4u1AtiR9h+qm+mgpS
S1e+4kkZtgTwkoHAvCKJ97OA0bya9ik50faPrSxI1l1smQl+XI/z/zNV0ZXV
c+QJcp6QY+5qeRgXRzMiB5W15P3xPNa3Cw2y+pdTV9TydGd0yihkpZWA41tc
6br1VEMLCBTR6PNpEMhxRHkbMJghMTNHE30ji6OPV/v6KOy4wfJ+jw/LNjm6
mF0Ew0KkEfUOhgM0aD4jl09wyxdHaLDkGxd1xSPG4EadT7bJZ4KE1R/wxrWO
XsfQ/G5gFQEe9fVLmN4nvPc2QdRr2Y7e9qs0b9bOlzkk1EwySgh934+Ndf8P
JurC2PJeIsUvNmXOT3KStiJ2AxWMzMfMS1oDZVQowwjTt0QI8pDniP+k05M3
lx54EzY+0K2Qw2SLPEEwU6Okm6QoqtMXVP+R+jFmYIpAZgORSuNyPSMINJg9
ZGs+a+y/RYd/1qqD3Cxdw7wo2G5IVOKPY9Kx66yMrJTfzWk9cvD8ZoZqlM3W
shz/t2Udg9oUIw+ftg/JEvsRUTW55P6ho+oXTSyYpckdXgnDn1OGtOSrLovX
RdmcoTb6/fYnZB/TcyfZ17cL7sVppImrOkgTDXTUit1xSl5K96/DVD1Hm1/m
62G8RLzvDFL+rNJ+VS3AER03cDhKGoCZ/5zmWzaRfn496bfoOqGYvtmOzSvn
h88JjduTxU11M4B5hKllbPgXRc+mrNubFyDgI4Ri/BoG0VH1TgAOyWXtO43i
VdpXHRIr5GNVP7NVKaxfjiHCf98JffXAia0ZWsOCSQPCWSJfHi4+idrLyzm+
hU4IajZOW4krxmc+QpMFSdQbClSVi0PWy+QWbLPxgBIIal2l+SvN6GWUWWrG
8Rz6sqTsDQy8g4NCp+/npmegQLUuk8GZI/p4EqhExm0cN9r3Xu7fsG/vBI4T
c6PNWsDNmU1d4k8WazL3jF+3lcnfXZW9nB+80VXHyC8S+pgzBxj5fBvRwSaH
ZECY7TQdsVIdrjAz2iioyxko0aVEkyfvdQYd8A7lCLcJL9aQf7pRe+A6pYde
m9FD1OaIm+pPcltwwzxn5A9nXkcffCgDxHyme7U94oXRSlHvAqKyHVbDm5FL
h32TphRiMSx/pFGq363gskj6xR+7LIfd10Im290pegJTq8Q2quwTBwEIau6a
ytk4JNWBgXXtu9h3wnoFwswK7XlqJz1atEqSpPUgKFBEGl/ZWbQ7zzNwp+vY
g7ty+cAaZuaWzZFWaR/YwngSQt4bRI+YAz0ZjKq2oN8NL4MN08anbTj3D4hY
yMnVsLOypIMKsuSimgaHxBH0/RH4J1u4KZmUSdKbmInIyiyHF/0rasAUYoMK
c646GnPfHY0UlcMI68+8LOJ/EE5TPUJH0Px5EugmBYsDTLTcKVXqOxw4W2DP
2Ylh+JYw7YNelBdux02yzIHbpuNm8wyt0axc+Iqpbbb8HPJYITmxMXJaC+xy
NUrXsMUQ29vaH50yUhVVph/Q7SfVpGaNumfCaBWoG4i1Jr6PYiuTDwOwUiZx
7hwuuK7vjZLc3XOANba3tdqPZ+i+gVGDtPJ1vVmjPGdb4AOTVpUD4NaZ5lUt
yeT/Bi9+2aTkce+XGfn5TA3BOTi0rjGYKWKrUNjpdyDG4ZjlIGRPUxePiHTS
Zz9C/YBtpmJwW3OfvKMRFrX2NEkFQlJVyZ21kX6/eF8UOBWmFfX6dmZ5Mw3c
ePMyujZMFJlicmTZG9u766im9f+2dkIaso1r6C0N9NCcsuXsigVW+Uwlql5N
GFWvcn01Ui55FJJLzVtqzb1mO315wiIx3EZ1Qm7VLD4NuRa/35lOHhX8ImEZ
5TexHbVYoH8W8RODcukXGBLN65v1Fv6DDh00BNxn6vHPtvRrR3uLmpqJXyAG
YNeIf9B2JTt2c+z8rchyDbYvYSfZJa8vcxdSa0QoabqzoBCqMxNgZFdESRC1
3kbgTOFkbg7TcBZzBBcXSSQ5SOYhl6/MgcgktKXzutOaso2x4sZIvxEpdzzF
mCZjSyKe6YiPFo9nbjFSLcuL00T1BCjcBNV3EjGfbl1fG0R8hs+LcBMSLLmH
BObfn8w8ke88hALeScQ0wL/cKxLIcHPvrOZVnkdqiRYHlju4h7eWlAXMYHxZ
VtZ7uAr/hBRFd/yevpQ7WADR/mDsRSz0NGew+Spnr8DQBrGOArlXhGsDtshU
dEoI9kIUuSzMwYvrjc0WN6sUpVNeW8oDD9YsmW9C6NpN2xRNUI8SznNlBeW9
hFdof2FBbzRGopmfdYjDDF4QapSj2rM/zIJ/Pepj/4fdCyWzGAEN3JNrccWK
cGIJQuxEk7tp3VQJrDoLMYjjGkYgposDxC0lJwjyp8RBhFXurJk6WPb7DIfx
3IkJK1uvdJ4msCu/tCOw5i5hcHdR0zsZhdzMQcihY7TXCQjAAQ9KNkM8UfTF
63oWlJjscCzmLCicDoU+NvIRJG68ooCa+Aub2NAV/CnIcwdxHKoiAtpGlP8R
T7uLg+jlGVN7p1HzsO+6jRng4KasZFwC5xVIfrd/y2AmdFJA0i81BfrwFb7g
6qaFq4nFrtiOFYoJ01xuPhGKEzy3TQ/ELMDBM+xVskmYS1xW8mnPVlUHmpma
QqUzox7lw5amexNBTkuf52dHVTXATg6PDEIMNKKPA1G11zJD/vGwh8LGGx1S
+YYmrV5dtouxnoTIOYhYSta7qkFfGndbUC5reqrnpt/pRJ5JkBDu5o5lMz7B
d3pK0i86HNHl4EGhHsMu/hEi6MpVpGTJ2/RDQ2ZwOShNKaDgS2COql+Mxcar
I0z8CysXDjNbZGu1mOn0ei6q4iLTYCxXXEoo1z8fhP9LrQx3zZuCFxlfrDFn
NseHOrjbVtawT3BlB5H8Xbz+UCrPTjREil40AiliRoqoMUqsB3jDjpivLj39
wGnchdMUJDtGHea8aV+kp857EsIU7rVqYu5SZG36ejb3jnoe2faumK1xGj4s
xZ9j5wnMh4JBsEtrez5o+Y6By8ET3gmhbFafdWoN3XKku9Hl/4yefrMcMFbw
cwvnkFXg3r2k7t1VNs3yWXjZVhkNTxJBt1U0Enq0NFnZUWs/E9CcqCdwru4N
wPuy0n/VKnIstA4QpQG50V1UBeAoqeiP2DsE+1JB6+WTOk5LnOM50hydNDeu
+R/dtI+N7193slSvK1c9PRqT7u0kZ1hFw6nmc4PFJP5xn8ybksApd7kcNGtO
2uvd/QrS5P6fZHjBgpVzSjP6qQGje86gmkzRX58WMPgp70bPxZvBe5AY4Dxd
esE3NIVQxcJiek2TdGaALqqhGlsmY+NYG50xXPwzyFWIEcdo5+d2M2z8JDWJ
tXYDFaFnAuClNm2cU67gie+t/ElloDBk0fC7cpRLxdENDd/f1kFtt8ko+JyX
nbn2pUWbTF9RPcRfDF25ik4L6oxgvO/tVXHYRM8mjHsYB2nCyqUHLm8oUB74
vuI0ySm4vr7W2R0tNAVcPuPLPza2Y1zbfJd6IyQkSGbPBzIYVcwK4jvKjw8U
KJCZ3XH1VC+c1eKgbAvBnUOvi5crxRqZgqejiUrp/HV4dGAnU83MvSGxbyk0
apzF+OmHGVSaHwyJgIXUiRzTUvE3TaCi/VcKQUcQw4LNuCX53avmbPXyOYC6
6yRq2p3mh77N457k5AxcH2+3WFRwSdvlVpT+QvvuRdKqe31dzBKkaoHg09XW
hO9WfZ2CtUPoD/k/g07NF2FiEgJirpOv76lPgHcEzj9CN8PDieB6k+fbu+ho
F0PShius+d9XLBQTUyGBCXliBboxZWGJMYejfiM06YS5sBqH/WeWU+WKJDpp
DOQImZ9rwHig9CnxK+TpZdgGwSU/dP5697lppNe/T7jHRfRjJH8kHjkg3/9N
2H8KrEdmTuujTLXLOKTSfGghloXcrT9HwugYo5g4os+M9BFDPi8aGjDC5hxZ
FoWwV6hZ+Rplhx4bydS3duYAFKmwxb83APBmsOca/rmpBRNU9a2woNbfa5et
i0n4IMCGUCMVzsKdxeQ6llXg+/Tj0boo4Vyu7kywxguhy8BwNVY5DyOpZkEB
OLcJPa88BmPyeuyiQdzc9bWpAM6xX9RYiJokzIjeEiy5HNinsQmfxbvGqKPk
509A4ZrQOG38CLeNKQT2e+oJcU3vpSzvt6UPehb8JI2IM9COtUWlf/AK3sNR
K7AbO6KY18B/EGnNjjXYYl1eT33tkkNpDNgKLDequuSHcg+XERnRUCipY6L5
wlHpH8aRyV7hmEI2OYlgqhHcAe//pSiLY9ckjC6KtHFTkxWnxoyoSIBXNOZl
m5OQliWhCHRj9FAHdSQUN+x5Hboh0mRkhh0yh7zhmoTKXhuxH0WnJWZMYlfs
RgCkTbytYQtuBGhhDUClGIIeO2/QjqfVbP6h6GIujJaPWzYDwfLZ6enSE2Uy
+r7CGd34ZIr6x4M5bZ7vb9953MD5xzWkYhJLnh+9Yd8bs66OvuDNX5CvxRwM
WQRPjCnfzs+3pMq/QhHC5K9C4tmKv3UfUU5o8HrnzSHPWDhku/HU66Yw+WLE
ttYX0kxX4jk47kYq0DC2113XCe5hEufU12oK+kRGOMAxfxIroV8Q9TwHj16a
Wh3BrE/UTqTNHBKdZdInetq71oQQUFeXqtUs+VM5n3vj9V8V+GO8RS7rEnZX
hBz2LqlDQbsS2/NELA1c5ACXti49DtnWbaNaRSq+ggoAbc+pxHbhL03CjWMz
F4CAt1BNhppcfYcMtzIRpCVWv6viJjK3iROEC4eVFVhHqc8lTzJBG04jZc2k
sMFzymay2UF9hpHwaXSswWXVEVv/J8dJwf8AxClA07d4pBgpRPTGoms9PhzE
bxcFKJtBZP35qNVbaYkvf1OiJvRh6Z+GUJ74cjSImwFXY3S3cy1kiP30nAnZ
qwiqjYm0kupZacorF1jmEVKlE6jVEvSJvWMQSNrfEUdJuVYKQ7WuukMI/V8A
6qigUsNmCsj9/8XY/4mrYagK+QdY14aexQ+Z0GwabPsPeLljjA+l3rY33meW
mtxZI6Toha7maRTT/C3o9eclC5gt8LViWGMMcvkr2zuuDj1ffn/2QNq5n3Yz
S77KxCiCa59bcstKdrRgv/N5rNM68nFtHbqxdEcgtjd/MULojvneXOFL+3VH
BLn9eB27zehsr2Z4CBdYBYXD47upNE59QHzydhFULdX2K04ulOEr63DaC8zl
HSf9bZKKKKKmbUgKnvBdHF/1UouNuQnJMoB6NvKA28EWaD6o9gIj1rCKaktY
49vLWBAVlaguRE9GRbb5soq2WaJL+jU22WHR2fSjISMMk+L5+CCCrGm0IYIg
VlzxYhiEtdHbDi0NZJ15ZvNPwBUCP6AJLGaWqMj6hkHZYBJACAy9gAY3vEhe
MpotBWkZB7ELDlnuV7Xqad5drW9r4ZPD9BYNWU/CkEKOOwQyYlUTMkFVHkFM
Sai56vkXhc4an6EMW9HDUbo+ZrjYVetIJjgLe+VXvIlMjHPvY4UxLpNJJhr2
M1B5AWQFkc7MEqWJgU7fqqbzUkxgYoesEOYyeEZEWtdRBCKkEtpKN/B2ai//
LHG1GYRxjAlF3sxPhxzRxcNuR8r4S8Q2mpiC0a6gvhGRh095e4pk1dnpDnQu
9HEknYchYBknbAiUa7+TEca/0VsGRIMsloLkHydrNKsdwgOCpuHKUgNgugvP
7hKhZQFVZFgFszJ6mMrj22xdxfJLop30/M38XjMWk1+0kugVzm7rE/NbSwM6
xD1kjHnA4BvjJpIajFacif8w8bgZHb95PD32uK/D4tvWPHaQnV+ts/rI9WYk
FFcFSJSftXEak2bWOdfmtUHc1bwN4waDzouVjM8hE7rU7EH0h0Ks43PixCt1
2ACwvNoIveO1/ula3OWLoAnvX+HRo1BEkGoCCezB5Hs21l6hMprsiLqs8YxQ
YakM9cLga3CqabzxgtklLRkzV6HwlDkYJ1xPcY7ICZ52RR+WtltFBDKw8QRO
z71/dqEjHr7ai/3ZmGuQ2COibdHuvWxTRYAdgsmW3wtpUbmmVxKxu5+VX8xB
5t/zW3YIyrUwhqwxH+WyCMW03JN/SwRY2rQM0zHsmyfIlMUS+TNf++Czwdvq
vjq2akicmNwJdgm91V6C3hT+2T3rjnCeBoVIRLJ06lz/cD296ViPkPpjZ/is
jpnFY5tQSOFa08i6X3++blgL/Bw5YmUIRt3y0hOnU276RSutsraGPZ6OJcMi
l3I9At6BU7VsRAemBSk67X1QIhoqTE0jEo51Tn/KlNRBR1VGzUgsumsJMZlC
UugH0xJcNTKmGAaFLic4LfwUVWyuj6veLxUDFQmXZ7arRAGOl3cgrqI8pokr
W2ajmBA12tsQ0VcFv4Bb+y3tUshswrmm9HRf8wqZgAP/aw6QMwQG+ABqNIIX
onI5LHXE9laSEPAG9Z9qr58bRQRKMIVEiF67xf3P535R4Z1oM+jBZEoR/wLt
1ufcm//TUrHdz+GiDBnpuB6mFw1NaJw1iTgA1+o+bTk+ob2eC+FEx8hGc3Mw
PclzMvYoXOfHab77Y4ve4sTVNa614UVUR7szLptIFHtlL7FRO/bjo0QW8y4m
emGlYdM+FBQZqJ7n0A+N620fUAmS/FJRwBOZwiOL/uw3/Ld0w2sllS9Box5h
qgWEOg3Cogk81xXOqAHtTu7HHbJeOM0asa5coiY+kWEduE5MWolssyGx1z93
//6mexCQD1hWHhbRVbN3ALo66ZQjBWXMkgp7ijRtMWsCCdCD4Y419zTNsQeN
c4Z8K9ACshTrBnjuC4nANngCJssjwzj2CWLsYx3mH6BXyBvOn61iBU4v55eU
fvHi228wMGXTt/4Ft82z80uKQv5kgvOe1AGX1C0bpj4dlZaOpsWpAJ4Z3Ivf
wDktvNJv5rghWtzCOZINwpuZ9BeDYfTNEtF4Hg4iKpMz0LB0K5+BKYAnrtfM
uzONV0LLeTJLMLOBaRA4mZGtvjT82mQEkXKtabPDA3HrJ1cGoSVKOvhvDiII
dMjFAiiIMOqCZ17Lzn+NWbGJ9HIkBdg3DEvLcFBiggNMEWDYMKqIcQydLJVp
BKbtC7zIGkAYjaY3dI9rwvlyO9xA/bMQqC2QCY25xk2YpS8bvFLArs70dfhK
f2kjRs1Hazo4Dv0myhlqB/WibgNLJyBBUCLdBISSyUsHo+jjUx4YbYVc7Jc0
lkGwpLwT0IIiCSimLA2+bfuufqonAIX9n4yjiXAluysKP+b+91oidddh7Of4
TRuyK/zQ42UX5z1u05FkseujChnU1ECtgImY9UYO3yzEM+gUU4z0rqdsuQxM
J/bXz67wRknSsIaJYOUDDS6JoXE4tAPrXQiDpEl9iCk6Y+PolfTK43AUWi0c
9it/cSWdz/sMKy7usAR28XYEK0HWJa9yUGaFKcywLxJR/sXI/Abuk9KUIsaN
UVc+zPeDgGx6wKMB3+5dSR8qBv7sUB6EDGbmYfX95XC76KRBnR+RzuVGwvSY
QpcsW+l5pXgsEj9+5S662jWYXVmolE5P8JWfDxOHMN2YU1W5RmVTr0CxQk7Y
e9NTkd1l2OMVCdVC9hg9IkQOW3gur2j4hKrJyvZg3PaGP54THiekWHp4cMAl
wL96k/+VUf9I1y5w7lBRVDPM4tqrG7FJYhsq89isihFTpoCpDv2u1fiGgx0f
NWqgm+bk5IXpas7L7isib0MEGziS1UVNIgZ2wTbVFdTkCtnij+PUlebOozKZ
eeY0KBqpDMQ1pqrw3POfu8UFUrILODTMnIgVzSW8orx4hM5EOwlybQlQ7dYd
ezn+5m+BEjhymVgWtVvQQ4IXoYsoGnSHBi77C5uBPBppnGg23e/IiVgES787
x6ZH2PWeMrd6+qlyhAm3u7sqrFxABPOp7KXY0yGUheGCKZUllYGnT3ijpgwi
VAcWpukvFvZQxdDEsaRBOIxefFTBn3p7E8nZHECS7TqPVb58ZyjpduliCZFP
/WecTj7cxLXnSUU30lV3t+PQ/cxjUKHUS0567y46mQX2aqpva+CFe66RKxE0
1IGCBU1u6jL4GZmPD0SsVxph00MW5zVu8eR9kgdOGcri5kVlEg/D84kQ0IaZ
rREDEgbdKVAZik3A+KOro+oYJPwNNnSpoox3iQ1EkLpyyL1IFoN7wdoenqtf
+tXrnxmZ/BmchpcfkKFH13C9VtIjYntOaUrhwtJP8sh4kNfCMY6f3+LV+RnK
z1SCfEq/bITAYZiLFOvFSegH8HFnDDDzTALGOnHXEV2bLXJNjTwcbXU9KTlU
iLpXTD4O+zkoc9a5xfmplIyISSCn7IqbKmW067n8OMER9tidxXWgLjHmx8U1
pWqyZoIQs6CnOBvGpa/sGVAZLBMxYXUb0YyL+x7eDnXNkT6Vxf2iiJljzexq
D06+1ikn0LrTPYOehmDKAtg//3kO1wACkVBKo94S7ibEwwS0SBJDy4VI3sqJ
3JrHcYC+fXPPJHu/brvAylPGb9Dzv09B4BgIK/GPWTmNoopfIR6EFUzl66HX
5lq5Rpp3k6xWlgIwcq/HybGmlkT4nbKJpBQSnZV9ZFvTZkTftOvHuSnu04ob
bYINz+v8DwN1Y7DlHc6sussTFj7EZnm7PJfz1BCbJh86Hm8sXxTo79RDcifq
3v8EEiBV9r3PKj//HmxWRGJqpQjI5bMohUFgogcxhoqX+UcUSohaamyokHNA
3/81y7VcKep/lhlz5dcCaFr9kyWkZMONH9J97CgfQ+pukj89epxRLGXCGWYP
VgOnBCDYm0PSrmiJMslf3GsFzlZIi/gquy/REgn75WMlkION7Nyky6RXjDmM
pSDYQKRm4/hlnbrXggrmG1kkt4ztO5ZnoqEI+D3O/WHXo28pYoECIO4h7Vhb
h3nVzG7+zkvLg/CqdRPIC6eLzYDkcVlHw/sBTrDoznDfxLK1bkdhqNaz44vV
CeQZhYdN7Hm/QeToY4vBs103lAlXcfEc3U9RL410tykYk/5Q3mS98AFLlOPY
DLR4VmcBmlDWNLC8WcpZxKA5oGQ8xOKzKfHv/gnL4HfmcI+YN7lRou/U8qFh
Z9obydTzMcZuC8earpjMMWRCzB/o3740JvFoSCpfz+i3rYmjvM715YUog3Nr
Qk6Zr8qlT5F9XPlPf9EDB5HPxcIJzkUK+6qgrrpoErsc9x1wKFXzoQ6P2eJp
X0Kzyc3gf5AtScweF9pAAM+fPUVZkMMF/+uu10kRS837gUpoVjZglDy2a6zv
3q46VWOqBE9lxuVAnTYnZ2y5XnIdcfcSSAhBlGIRfFXmFnCQIl2revE0jHuN
CqbMzxM9/cIjusJIVZ/PRiRJbGH/Q5XF9vkNAk3lSFnsM9/iXNmMEmP4dEc8
Sb+RigoreoPYIspkhT4LFLewQ34mGsJdvBG241djYr4bPoY5IHWYJVkxs4fA
cjfFyaMU6/kCrQnYBPx8eHWUMFsOaJ7km2B9dClxph1RHYaCQ64PDnHmPzdu
qupl23M8jat11BVObbCIp7FKOyDiP3ZWs4+KZeWWM/d5/umaZfwqJQaFNvJ2
VjLzdUoTk1Eqkwvk7d9wB4c2UDKIvF7OrBDCjtqAkETUEEpMZAeUafF8n1fD
DXiJZwt27g6pEcmoJDXICcQwz7HKobbAWR7bimiuGqc+WURVnFns+uU6pqvx
AVbC+MVOr9oySu4o4DmFdB6ykjgjVAlMXbw+Nxm51Bx2M1aPm1OuNAFkXVXf
RM0S6TbHGNpB/EOApioe6eGk51aw8ZszD3SDJBosjn7U0TJTRXr3gxiQ1bl6
6++cBw15Y0FEBMzKzhPiQIEk9ShL/vXXnueHCp4ZyIdk0NV+VYrlOcJ3L/tG
i0dReiMRvAYBhXutf/nCdn7mVXQiBeYoaeVsD8nx8Sb8Z/PZqbVoTqZBppJC
3EVT1qVyXVwvx/i+kIDV5BvMtbsJSiuUoZtm0aEfx++Y+tzr5+ubdzVX6Pwd
xbAQECKXoxgnLwVKdCCbug2j94M1nZypUgeQSMPd5V6DJk+Il45HFzIiEJ/v
2jcmJQF/vfxCUku4JtYEIrePnanbbgfuUukZB67YQxSfL8+8LSiMz3flVY0s
7ZPXxpWmcKa08YLITD5pEqPyLYtoxEZienj8gcF8MHUpSJ1ciJQTN94bqOnS
JuIfCbcctu1hdzEw19fQvTe0Ig9bQGZPiahLuzrvBNSYwEEgCi5VOKAgtKie
CEHk+YjKcPiq7Uv1aiu0zGNankuAaaEMWSEQb02cMP992Ll3TtUxG+sVYt1H
SwrW/iU5WdE4JXDyTIwsgZSFiuZmeJdH4ydNUXsu9jIp92xvCnXBpvhf76p9
aAcMtYw6mGWuTrZx2mmbMeQ47v3V5dTJAmmcrmpRmHULMrUZQ/VOalIBZq4V
GeTSZbSp0Td5QhEiqiA4ON5HUMaPOFf0+Ch3PomgTdoDIEg17EiYoK917sM3
R1yahCoxnHSu2MarkTaKT19pVKSOyxhJMSyi0H7mqNeVdvJuigqBmg6JpPLS
UsvOcRzc+QlvYziaGff6Sq27YtlvbYIhh4mr7E0OfbEKP07zFQwjQrKsNDqG
PsPWeUkcFIScFzBuzeNfyHVSqZqRYaYLOvD6kAxJpajvPrBB+1UJvbzg0LRp
MwCDVrSfQAWobVgX2QNHrB1D/vcG6SSuSh7OZPuZMLXExKXutBC8jAeq1Ywr
uzucHzMTbksOXBXaGY5S+zUX+pKaEaWrRHptsgCnh3Tb8pVf/M5PxKue7Dhc
NnF+7TPnCvJEmZ5tPavBlH6QIMJpdYp+GZIvgAeSIDwjV0fGcqto1lUnxCPK
gH5cAq4gqG8rsz7aa33kCeWOw2vg4haIDMMZJY0CpavxHaGNGPGn4upTRiM5
1t+albvIGVDgLTVKrkjUEaRPYXsolMn6eyRnBTHrex88aDrB/ROPhJtJ76ub
LNHggI3AiGEzKNttJNhu73ASHfa1K/DlhoW/Gr28aiYIXIFvoXhv5jzddIOb
oe8YbTRG9+u+YvSdesIxdF9eQ2ZY083LNqstW98PotNEDD8UcQm2OTH2U9nK
PRvaxuVNnr1TJuyJRb1NSXR5JKJqcQ9311U3c+kXJCGgOoIlJaJ8qF/oXvDk
/Hj3lD1nVN5tJXW0XPjue9IGzohRLpFoNPXu2oTf6FbbZzo4oP5Fh50gC6q1
8rFjeFo/fMUvoHLpb0njCgKUfxXJg/Qn7egiibVLpg6QIIuQ8O3AfyPDaqFM
376+v6PUZRJWVqco1WGVZf3UhQYAj2HWUXh6mPfmOVxlEEzKv9ksM1LbZQU/
Qb45NJT/Fm31HdZ5Z7hs/Qnm3YeP2bS5gC8f8FWt+e1s8D4cFn19TEVh8rqa
Rj1TNtm+1pJoUpmwN1doGueDyR9iz42ETYSHh21GP62ERwTq6UpDRrfJk0ZS
qO+n63lrOpIRvI0LH9YfJOndLlULvbHwRPyceGtxZXfBO+12si37NgFwq9+6
lpTymdfQkJ84jf4uJCORUFBdRotlLvnDCjF2RNV6fJ4DifmSe7w3Htt7EWa2
OZkK/ah0KGYDNieH8W2x4fYpzbkqZmNXVvrNP3Oe/aDhCiqgUqdWrjTdRCbZ
cyh24qw1yi6zKwFXJ09RJy/PtoTtxaiGjbqKm6IKdhP1Ch3XB6R9pfO6oT0D
ZlkQ6e6LiHl1r/KZXXN/+Z78IWcLitqiVcmTjghNE3N7qQlVZyC9b/wBU2DE
y7JioPU1G1h4y60Y632hVvynN3cvVJ0szgiwTv+hCYA3Jvz7WDBWec4Q4Hr5
RqTKNxLBauCt4SFzrcqKYQOFBGT9PZRB3UihGwqjQREk8DqXEyeh8Ut+d1Y+
wzbdi+od7MvXykLTLa8i8jw7An5BgOwRXNaBkARnoRt07pMYIVD53kyQRPR7
5+1B9KcYUo8HtcBPoS0pyfc30r19wMXjwxFD7fLDb4QJgk63iKSS1o+BiwMJ
lF1z6wA0CBxXzIRhcOSClduii7y3g0P7kcu8TGPjJZ1i9cI329sYuuPj3hoC
yhmoluVrSlqRqMKF97mhNM1zYb9CxsCkcG2HkK78Ex47bPMGhXwBOUabGBYj
UYA1hhXlY19mh5DdIspgVIanVljsnfxz8JdjFRwfn6CodvAArzTzmJEjYjZs
wXtPX87Hz+jNzYL0kDFBuGVJKYcrAJr7Lg92eutEHyqarFWhqmsXGVQkKmyH
9au880uAuM48afKmaftTtXvuDMT7lzqZnXpjAskOEZvfmn+Eeu56nThxDl7q
ptQFCU/n0iKJNG8msJJ5oPdqItJKdK3txSiQBwKxqoLMNSB1BHQcRXQgFAFP
qzf/oqY/xH+SiBReHGtXApXxiYFI6buu9UdoVr5tJqd6u0ey6fdOSK+xs5Gb
TzBSErX6jKAXBqf0oLA/1PbM5UQ1Tt3pLEejE8t0ngbHgPILuKYWybD/XNZa
GQJdSFuxki4Kw/a831WSjk3q2sECR6LeqNB5qcChOFcT9fi1ZBRCrWG6Fp7M
nKjjeEx9zVacIe7K+153jex8LipkIfLDOIap8eGKQuY6krwUd6jsJerFxj81
LCVSQvFa+z89a/CuF346gz6hlaC7Jk5pOla0EWN6LNETAfKv+b9UsnEvsl3y
ktfBdRi0wgLUNAW3pYIHPKKpwsNvCGXi5TUH3fdlL43lc9wbOFrrHrYKVXD0
ukETYJn2g+nIuJ/xDy8vIP9qZ+kv2n9j/SbiGeT/xu96l9gTVkgIR8Q+zGEL
MW/s0ET/0+mMHVM11qZO7hYNNPyCGUBvt5RHyd9W8SfsxGiMh/4EfMPQGdjS
kWkI0APm7+MPUf1YwoSxWkKCDBo8iQ05hXCgxtkDtHFnxzPpbc+AIoVHRmr5
Z5U/lDgwrTpUfXMnphfxYX++CWxwM6xowl+Z/nwI+0bgHy8osm8kaFZOk7vg
lzBT0SOceyTZt+8zsgw+mjf6YxmnnagAT3FrLh7b/US6tvN0GuCz38riwo7l
RwtGeCQNLmt9Q6wLWbzBefueJE8KIMHD0Qi6oy+5I5Lize+IP4CtFXAFZJSp
OdWexOlvOFSHbVwB8GjkSmtEDTORPAQMJxx3hcmUJgkou8PGEjdfD+mJO7Pz
CO3g7fWrkSCe4WUEXPUNXf0cS6czaJRSEZt3wTw1Ml9hDel3Cgg47OL0XNbc
WmWXtg41zDrrC7SA9PXoDZ4Vzx8jDRKntE9p9mvK/ALx9UGUIaGSsnQsgz0m
eKBUPTDLPJLaYVIvUs1mH0g8/eLOMwv67Ck0guBkdx2Aq/WFx08UbfAv4nwq
c8bGAwSYkE0dEaZxajZW6DRNGSHqnusIiSDb/l00yk6zLZMX0zpO8QYlo38Q
Q8Vj2HuJd//k8/2es1Q0QAbAqC9BdoIrPqP1Z+rxxRF93IxBFVNxou9qtM3y
rYIyHg6qUxWK/lB7wV4W5gN5R2Q3OlGt5kWxtBNkWvIVJVL8Nzv/kIDkV49o
s+oT9QhcY/ZY3O2Acq8OQz+bfM9zUFHmc1hChGTlBOPoI92rv2ys0E6QsjFJ
LOjCSBrJsl0dLbt/qY6bnNL0BNp4Gbd37fiNhquepePKWPbLvP91u4hZ1XcC
6pSPKZD0SPUI2eCz+plpxMswlFmKwyMomcLuMcWdEO59teILVpStn8HA0jAa
hF5lbvotN9sgMeVzUmkvVO/D6kKp3eaajDJy28hVcv5r6Ob2FgiU2n5kW8vm
3qfLJfPj50TUZ1tEfjvAn/3iQ6vrqw/o1RXBWh5UZYUo5H5moMWZiMr49DoW
YQSnrRL/q6XPs5dZJ83zP3f+ANjpl9ApJiK3GSkfYNerm0vcujC6WtJyOq1t
EigskbKjIgVJiN7rg4XKnTnsKx6DzHA3FVlcryRYksVdexXqby3Kn2RY/JGR
38wzXCvcNR1owroySXC7yBnaM4Y9BUZhC3S3iA2KcPbjdZfl8Y3fM/36D4NQ
vbTVZqkG0PmMavySHNQM1ZihX1kkRtdSQBT9HaNs7tz44CH2VO2cuszfyYJA
qs5kuVVH6UJcSXPnbXqAwDF1MomSQMml3CYQtnWu841TB4uDK5GsF8pZs6sZ
tmux2ouVFfWbokX1vNmCJLmp58xgIO1ECb6tVAv1sVvpp/WaGOc1+RpskY4Y
vpyAbFHOUP7uMZbBSOx6/ktMHFgjIB02Voh41AmmqlLrVMg1VBfcST5gv8uh
CRnUcOF/OdcREW0gyxtCV/7FAJRBlAl1sM22dfq3+7TVeWdRfL9f2gttGK1X
Z8XG0mOGGEgBUPWcXRFxw9Fq1S27V+BZb1qm/669Wwm9F/AZBuRvF1MCMAix
yrF7nbGpwSZD7bsChKQhJIMpQ1BijgfaFUohNPiYHDgydtML/bA2Pl3USLQM
o4Y2fDlKu3DTlMoh6rt2DhMJY7SV7KN783CfPJN0T5bPey41+3ucbJ1vRX7h
olyCQEbbZQGOwQ4/i9Kle2LglhNjAWqb7jzW3aagSpIC3M3j8py5Z+ClDfUv
uCPRu7MPWsZmi50JmubDCOSXsWRehJ+pMzsNtb89u7TUo3/1myumuTQoEZkE
+R0ZINNN58b1oqV3ZGs3uLbvpuuNRWRbgnedMaBjAzafJbSUllZ/HMicBy+Z
ew5QX5v9gqm59j6lYhkgNuCi9YMsEmVCgrvIkRfvFUa0WOxmc2Iq+ZESduAS
3aJ/JbTUSDUKbYAMicE8QYbLjfUU3/4dTmy928K6AZjFJvYjYsEaK6kl6rUy
c36f12l73P/K7I8orL8px5xf5+amVYFmXEmNemIDykFQn+zxA7n+CX7jUW5M
gPztuckVCc+HPywJewewY8i6K5alozdNOG5By+pNfNmafcF+E/ybJn8lDjHU
C/iC8oJgijyn5+Dn9basny1gsf45mdZUi3yBxDrrf8PgUMJfDKv4u1YbVUsc
fRMo4HGNGN8FgSs7+rte2Nv4vdZTWoB6k8h/p/K+NpTa7Pj/8cHMH6ZdziAS
f/pQ4b7YpNMCIBXNFsIFQsZFZA4evv1ZOmf3oo/e/VTlEWL/P6v0PVtiGKm/
Mv1+stoBuYVvLgOU9w/e0t4TDFRAuTe2U9xZiD8ZyH4MaYQT+KNFyTagm53/
rnYNOVemFA5pbyrQu1FGLkLGcfrGYHqhs7szHliF+tPQpR82hOAjvSkDv1ma
6xCxnwBZ8colDaCuj/QdNgG7zcOsc/4Li7qWwF0pn1vzZOHbIzZSh9VCjWIg
1DjFIHBvsxpNndMNhdI3iZR30XzadA5OSKzN4SH0/HyHrSoAbQra8X6H6Bue
vZEQQYx2tUqwy7lHiq8VGiSLgCIV9942Ek4uegvClxmvwUZ305oW3iSJ7orI
+si4qpVY6YRkJ+AwFdMF5jtsOz7gyfxJvzD4Z9h/VhXOcjyopcbgWldvptC7
EdgleFA85SZaWuMF4HT/GQaTSGo9fJoLKBPa2RNUtRhpKog3Jb4bBgRzgZ2I
fnVbZGQ2s15ASYulRF1CZi0S5OnB9lQ++PB76346D/Uf/DV4hqYCLziRQHu3
eNep4+g/fNo9PNeP0jCq22iX7THpm9yqZVgOFj8fG6aiocl5z+ELkaq6NWIY
xTCc6aT0G3bIw6SlbfNIONsdSfSZqj+TFE3TAXpJjQPCriLx1JvvgaE8kRoq
x8xXGnUEFibTD+0SrGri7kb3NYjIOjLxxWSLzRt6eDqtPLq5yHUwBJrHutuu
3zqZcorivY5wSbLq23ng5LaRfB7Au/lPmFn/HsjbMnXbdccaMJSrWWb7jOIZ
0BDaDXZW9TjfQizfEpWkoxhBjasx3SpwRrKbhYy7NgTlKAsKapiOqEpZynJl
2OCM608SZvA8QXnPphencxO6zBwp7UPXL6qRP98Llhpx208QMwHD9MenkuQZ
OHGjlOnVXNgtkp+RqY3H9DmgRTqiBSm7b5b+a8nKa7QdsYewVYHPBHDbRPgR
I/o4kGlOFMwtpDmlRLnkvCMQSNZlpHyEaXHP/BjhIImhup4/2XyShR/vYhba
kvDIeE9RxuG/Nc/zwWJRjTBqtUM9AdzcDII1z2Ok/0WbRkbx3yMzkYcZViNv
gVAnnrwoAsItsRistxRx+QYZ2jNX//wuaEXB3vNW6ngggvXHqbukFeGzz386
36QPEWbB5+5UeCv1f0uxUeIbxxSRST1u0TriyTPOfGduvexJ3CsSfsmMml2j
XPhxzwuenEjUYTdloVi0lFGwXU/RxpvZM/jVI5/yOTLqGkoKVilLvcUnNGN/
gIlOPq+EOwlB369toOyjUBvkBKxJvRPNgNKUIFLh8ThmCDTMOrEjVEyKPmqi
aQHZYgSI+JceOhUIUPbgzlw3cgVFZfjM/K6j8EReIdVKsXJzUn0YA92hmoim
0uKkwq7DdR0JoWCuM3ZJgEE3lnj2nGYkITrT5RfHcz+7e3BcuDLuIzLjd2yx
tWdbdDEq/3SGcfphrpWUogrCqH4YXDoMm9vGLKfwoZSR4tJxhKx3xM+wKZid
sUbE5wBXetLCekGVuTKpBgPiDhyGAdDHE3fCBCcCuQeYQKvawACoeeQgNQNw
O7y094hglDeAaPWGfvLkQI0I+UT36mdlOjIFnGfF01WQOU5XxRGh71FOu2lC
Y26RaD593dqrJx4FblLQmal2xNlkKvVYT361y++yZKKr9xZg0R03l4gs5J1P
R2Tk0j+iGnRow6VjVps+/Y3tVswc9ZbWrvmj+yjclNm+QeftFirAf0pVb4gT
pmAlAVMoJmwqnTdXGoF1YXoYakBjoF38iBSgsx6JxQae65qmfQKSWABLyRJ6
jLDrO62MHlKkjTRIw/754CVs+UT0lISKl/6sR0NOoWg6vDkqKxGOe7oHR4yr
qlKWj/mxZ67AjuQWipZ/KSgG2jw1q5U+db5G0Tl/d44BHtzmhh84zFIU3Ba1
92f9JyhlkEru3byemSeTYRKUUG9muuNKJEdp0mf4d+RJvom/6A/S+Z4azUXK
c09RHkJ2i6Xze0vgoM/g8oOY7g4X9k+f5MVkx5+1DDSlsSJhnCcM9ZjgwaBb
tL/QRq/Od96s1DiT4UsZjp10SdKkYGTyCHd2s/ryRWMtBTpcPtcNQ2oGT9FD
txBjgONeoqM3QPy98EC5wrpH8nXts1dYCdhnTa2876lPUlUFhljNDvzkW5FG
Y48ofuQRnQ7lrN+nx0uR+6NXRa2b9Me4SBdrHWSpGCwtlc/lUr/YK0VZfP03
szO/e3qK0DZK/zjAMeBXjte39f9T2w3cStJMGfIEZSCKWyvAlxA72Tg7/kBd
sA2SjMRyS7InqK5mKl2hxv5GwTXW22DldJiYnCWUbGsGvma4vUjLVBViNGOY
5TZ/p6k9+JW+8gEaRaGpq7lM2NHkoMcuKFfd5T7ZKBtfn4fFw5h5vj2ZXUmV
CsNfnmaDL61odag4h/L123ahkgysyHXNe+lgWrgUSEwkGpCkmpl1aR9VFXuo
J67//7pqIx6Vz1a63vx8izXTCMRWc5OlsjztL7FXDNTt8YB816IVJmYtbEjd
TXr/p6qjSfKtoqCRnEI80GUq3a2dxM5UR37/YVz1Le9VBqAcyc8VMgQZdQW5
EpTQaNMjzrcsRt00y8uquxzcPuq0ZDMbS74W0FkRVSdEgDVKGzvGwhGpbSJc
WL0JWC+Z2qDLrMwqCSQL5sph5Qi47c/2tBGkpu9KTXbv87rJLuPvXgUZWc2i
SNSkdWH1k+/cBSN02XUSfDt75dZyhqMNE50dCvzWBPWBcb6qvYze7rToDS7k
7/VFZbCAr0pBjmXMy9n620bwM/DoV1NWx86w+7uPdqkPPoT/UjJv9xvTzhaB
jA8qUTLYOObrPMtL2plB/CqdxFY47a9nzPH/80Z1QFpTlyO7nOnvVtyshJyo
mbaZtSulcnqBm1Z8Q21qPQYH1QQ0J+u+AZoxQyE0f9/72CXFv4Xp+jS3+hqc
ACzBOUfjm3ENFF6jn/3BLvDECSL7nC6HeOIFG65+WM/7XTh8itNv/2LJs2Wn
gXpjjhAEAFD55qml5yD0+lQmYoWxrONj9ZxMriX7N4zneXq+KWtGjEVE1Cwp
Ej6TomTlxXF0AZ+0T7esnZd3OeonLJVaXHVBBldkdp5FMqFcIc9OPGTf2Hde
Z7UZmD1/r+EJZvPSdxZ34+uLzzjLxSI00FJ1AuYPxsDyNh7tv0YfPymd2V8d
OgjYDZ0cX8Rk40mxqFOURt7F4vmf6cmvEWYLgSjhq/aWjl/nZFdQJodb/ATl
OoqiB9QdzyvDPem7AOkJ7sCSua1H2kXjulHlEhwfmR7ptoUOXd73JmjsKl1X
LZnnn6i02g9MnxuakvJ+g/6yByJg/Ja9BswkK0/220TcwWtlvh5Mih2aVTJS
Jku/JoZPau22gfjBKmbUHywOUzJBuMP/IgOk0UkFMG3SkmcKl5pJxV1xzIrG
5bgTCGQmZfr2HbmW4YAQYNh5R+v6DJ1jAwzzE6tv13wFL9RVzWJ0gIGfLcnQ
vyfxBDKBSYcmTh3jdLwX8cHg1SacmSfY04yqjmoPC9wu5fCIZ+9NAPgByWFc
yBd+k4Mus/TfkYrN7ACWeQ1yJ/8DqCfDLb39XeFW3GFqkMBH/2e3Ad/omDqC
m+FgCGCAMZjPtJUfgJH/Ah+JWQpnWe5AZL97pj6BYkQJPINPdo3CTH4F6FwN
UC4Knc9JiqagO2NFs4LHgxk/Om0cxPEfrzF6OMEgj6BTI8IvyoVRnlXQHJfv
hSDmUBx5ksc5JI6PyM+v3l0qu9rFs2CD6sX8a3oKIyid54jmzo6twpusiQCU
GCRsjrUP7frtS+74J/9S8H70q1e3pxtu9QvG2HhhpwSPYKwkuryGRdlTHUaX
a+G23IK6iCypWX2Go7LcGDboDtIFd3coW94jfsVTdFhDykTBkCNxB0Zm3rwu
eIvm86SYtUz+kLcAypUDxSMZ28rpp78Aut1ivsJFukHx59n7fWJCJGDyPvCj
gs01JkrfyAZO9wuHbtx7p9ri9P4MfCD0vDJkOG3amPafV2UGxnRACobhI6AD
ASh6V5v70Geuf+Lv/DugnDkRj6MBWCDrW6QojIi61JB2F/1p+Y+1H5X2ic8U
RJ3vchzqvJYxhQWDW0zelQXG8fpqU4jrH3prhmRRdG1oCFCoVoZxM+R+pYOm
TcHVMow3EAPeEUesxC1vmL/KkL/sB96Q+LzMpQJlbacsvbeLFEuzvym3J4Ts
naZfXcqE7Sjx6jPgFpqorpvrazGj6YHTpv+lYM2X1ZzET7tyEsRF+DpgLtW0
1jliquml1h8KnSafYMsmK6P8tk2Hl3KPD4LqpZxs0eG26TD49vN5pabpUiai
WJzBVgR0MIfIST+FEqjjHLzFAnSNVawZqKIu9rte6IhNe/rT0V3K5skU7iZL
sSpVqUZxXvRhdU9uFQtZjSbaJkx47P+WSqxYNabAJCt310BhTJOD/4/1FkMJ
T9Z/PHVN+o8GlOMlSmNADe7zmEKcMlP/aYFTz4yfANcl0RRUuIsxAAEVxRpU
MXW+K3OSlOJzaRt90wMj4usiDR+AcIkRm9OIq8LsgLdCDTK0qmtG2ZBykgEE
ydQ9NYTMNemtnhPK3vBmDYktmzkmMwVHKF68lxOfBiTCsq6cehrJIwcff/+U
mPsQVE+J2UzzZAE4Wc+JvIH+6JHGENrHJ3G/JsyF9O2TFdaS1CiHpK+iMCFy
vvbZje9RFNv1RCZLaLOXUMzw2gXP3rxWxw0UPVDRpg1gGvqUtPuX0AtlDaDb
zaDcNh2b4ItpCZ/H5wq3wJxmkoEqt8Sw5vtq8ca+Iw+BdgybzGIMlGaXasx3
QEWrUrrVuDTvbo/bxoj/pWd0bDSuoUlKrBmzUbTKrSGsGGi3rBJ3vKEEdVtw
uiUURkla05MXD6NCllNUmjNZ2ryIK5LZVIvyZqKS9IJ7S401BH3WLiffFrzr
f9QQj6jxIyyO7EeqVBxOHOQP/yKWrPKbcYQFkcbqPCegNU/aBFKh6iFufB8J
WmQ+kApsNuyuzNeFZ3OiowohxhS1VUIFCpZPdQaom4V4VJ50eb2pyNmrIN4Q
/fhx7U5tTZcs3S5sj7aTK0Nk43QxWqAa9WlUViOK/ZOsacKI9JDHgPYFZomr
wxwr0dCLQtS2yWyVE1Q/xs6LZOyjqsgQQUA0CNWXp9eM/Z7hnEQ4U/zEtl6N
awIWsMZ8SM4n55urcp2pZw/yq5EFyz81++U+H0Kv7Mgvpw6ObdM3ZDyVlgyh
9s2usfW7Jzoa6i2QN14Zln5vM4Z8bFJco3uYziziSXJxAl7ztak6aZA/4hl4
vpSqNoNQ0WFPyhEBxg9WsgKbeRXCrvIo6Q+nsHKXw0F/kQa6yY4K9HMP/d4l
JeEqGwXauzGmvqjb7TfTHis05F80VCO3fhWJZKSzhlA1SDJAfZnvX+vvsB0k
4wKJeAWeb7FdG0TqjOcXYR5MjDaUTFCV+w/Nk90fESHL7NPocEFFA0e7tVsX
tFDv++RwIlHMfjtRo4MHMxYmgG68iZX4PzTywIESXRFnhaXnvF6SDX/04eWN
+jKAgBvDooyGDV5+DM2Gtoa9Rdd7gsn5t4eNTCblkK943ZotBmFU42qO4n2D
T+xud7PBUbSuzZxO3DtHEMhASJe8ecBzMJ0szjG+B9TW0N0KEUFGztlV9Bh4
MTiyzqToOLwMoUa1GrBaIpsEJYlvfj6r2YoADVxPp0ZEa6mcTiCdAXCclO7j
rU3qilnohajam8lbS2q2rlKR41jOL1gACEXL/FiZ8fTGsnekm1mpQLt3EhLK
6zlhIPwLPaDwe23pxDRoUWoZ6RVpHcXUjPI+5Yd9BiMqPsYUslpQotuAHx/B
gUVOtsYTHkkIMPnKKXvZC0YxFHq6+sBcIrbOS1DGI2tLgits4J3Ee+/cDK6g
97eT9FCzMo0vIK0LP9jthtSBB60aTXDiYX8LU6kQK+8f0RxWdy3qm9+MkwZX
/L4ZzSlegWy6cJtsS+caBSRTkz6SgolQ3vvImvUJyA8Yj/sGMvavsC7FlldS
I3r5CIvmYyNIk+NCOuvfscNqQZnP1igflOSiq4+A+qRAeHeb92BTSX93x8eM
dLfXG0s4qMSIo0ciYabNFHRg+Rq3Wd0VjuKhmiiTJ0ahaZP9XHfX/O242K/6
/sZ5qUWFFTwg0MsWbJigHQVxYotzMMXLooF5pQhs1a0l2DID2SGl8Utfe73n
xTxN1MGbAAprzCTg2s7qgdVj1cHhoDYA2Sgo6/4e8aPdIJ6IYyD5X7lF5npe
v/ndfTJbts74hcwa1JLnDUN9TLvZKqC7jJsENLZ5uvTgKc8Xdtj8FhymTqah
azKjVSuMbAXr7ybAZSgCKXnEXy+7u7pp3ES3DQEyr04jJ+mYHOgm3TsqwWd0
yklynWjR4/xmkYPt1IaELPBrZD5VUFJa51rAR1yqW2ybPkFpRBLoRLmop/ip
VM757/awPKXKYRFVuBiMAoplLUcIWkgRlvExdzhpaeWSVHkeR7vmpNBxP4q1
jRKgpYlpPaQSDjp+NAqYkc+N2xK3o5yQfuah6nGUHOBcztiHjgZXL+wAm7du
y7/HOUWYTr9DbEyAygm2ooc4Wz7VGNp9OcNCXM3Bn5tAmccp8ANzF/cQqBNw
zBWNCK4/EUZqC3UouwloWmikIb7QOimQyt8Ay/trsmqLNEiOWbiLh46/uUVy
DwHDQ2Z8upJ+H+7P0NelEzPLSXZca0hykHvytAOH5JSBoQItmx66Ijzhx84m
Sh2EW/zfk05RGgLvRhzrxBhP2aOTFQ9+iA/9kavAHBDV3VQgLoAkC5ZZ8tGa
CYgzq4tgYda2xbohv4I0+ROpVLGMs8KdYhEns/n6L6tqbwbMBA+UhC4RdIXO
WFXTYjj2QrbpTwoPB34Ey4ebtV6PcYjk6xBwI0/nMi+9lwSeJDRTY7DFTxdf
qpjvLZgpwtipRSBloRfoBxyz/dJ6Tg2gyFgYK4AlsgzVLSIuQ/UqccJpRyBq
d9rQhX4ZueCU8OMw233827wAqXoJ1Sf8rVWDAbviEszThKq6n2dkaD72+V12
ZJulM0FGVMEAF2tHvCyuSxln6TzPLhJDKbsTegZlEDsXqMJlGeSsqt3ALs88
r+8hMuFrDTWri68aTQ8JMTEEIdzkTPm3X4uBRchRBVr9ivVpaDKoL+1RP+ra
xxeobcxTx/b4dJh5yF+uKuB5CVPHL0QupJnWMaEkuwXP/7JrOgko3ihDsqyE
0FRXj2Cj9Dly+P2Ba5gxS3fylOjyfpwpV7NnbNxR8urEA2iNTgiRSxrTUWPZ
ds6n9MUt5FMHkaC/O8/ijkaBQeyVaJjkdFWP54i4NnoQV65PFxX6JXeH/NO6
U10JGYYWnRFbhRA1FHdTfHQE3dD2mefsgChQJJRepUjdNVQUl4HpD139PmYx
dG0cERXSxykw38/5OVPAuTMU+O8QIWJNUL1liGB0Xzg54vbHenT7QzvIc6Jp
bc0/nW+YOYFpMov0fqd6ZXi4JbCUywhBGThFS7v5wocK/yF7c+u48HsYnRCp
ybEmmVBS5PJB10GrU2cZ764FwiNixXwsZmZVyBULOzsDgF88+kupvIId/u1m
oXuX2oFDXNdSqiHyJDtaMFY3pKTBS7JrSXULSedrIrz7GV4+PCYOhN016Tg8
Fynbl2lTwbUTxJeTkv8dbparXqubu0pDnfoGznWGAqEHOjzbMGRyuPurJX24
i9O4XeB4cRmJgIZOW3GhfxNebwkBEPlJNcA4tYa2Top1hJ4vFDjddloocHYt
chHsZvcIq9lc6HoKCX+dcvY2JugCO/YTlm0EL9Gw5dIHE2eeqWRpzKs960Kx
HkX+8YgsBvlo//NokKKrjTAW0xfJ+wgNCNTb+U149DTJijxsXWOC+yKdrMLR
b3YuKcDvQpLmatGvmPBWfgZsJJN/GNtmsMj9Hju7NRNajNJLvrIY7yTwlQUj
ilV292YhxVah8S/AGIR7sUQibfsP+fw2q5ifM+7m7Kula2Bbpo1IrTxnYIWs
4J2KbmIOyAI99qsmmURmxGPoMd2hpgWlss9QBy42Q0OF0Ir7vV4LNfj7SOdQ
RtYDkHi6Ka+UtMoJMfYYumoFpkp+iZB/0XKJP19L5Q7rnUZBm4gEtzxBAiyV
FRBLmrAHiBDHbw5E5ibvWjjGz80Ln9vcgo+HM7v+eE1eckjAlm2zTFRi6AqR
DRB++3XfpHqqR8aqGvkSFwmIzwfi0qo8rA0giOw0ZBotm2Z4Z03I9K9I3ITu
Zoq/oAf+5qs+ogRspkRJZdNIv24XO/EBm5r2df9SDqqWraJR5mKe6P66t3Qx
dtqMZ38kcx/06ru9Wj7M9wl5xhqiS+DEN4ihzesA2x4THKmGf6s/vcTosFwJ
jagMc5ro2FEGcH9kksnKWMmdQ1E0ISVyJKfYJAPizlCijuyK6sRotsh/Wzau
oQ4pWlfudXc5Jw0ERIQEi6ZImhDVwkhIy+jvA1g5vs6JBUiaGeVTawhIY2hh
lz4LT+ZU+9WvdABF2lceDiAzSXk8zrjPkptc7jcJlOWNIe9oar9FYPxHa8hv
Epkl0bxODPpVx5i2Y495KarauX51diXxyp9SoC72kPwY27OAjpMVc1vYM+GF
iWpJDNdWr6hHu6X2RJa3bUzMcEH7FaQuiNLOPF9Fw+3s/dzLNBJ6P1Kcv3xk
EUVmtSApAbVKGrsZCxNaa7TQqFb8u5/kg48+sQ8a5H+6xWrqU24EHC4wfh2V
uf24AcnHusYnBnerSFvpfeuEwPIz+eHGz49x2hLJH0MIODDH08dmpLsFIK4m
ZriFHSIsHLFrhXq96sgsv4vySRlxqA+lgmAEK1Xqc8lwxKHFgyhjQRAa7Mf7
1JeMTh3z2Jp40nPMIC6YnRUM3j+9R+SoqjrWiwXE5E8EkPilb+K2pp6cEXZB
83OFZgTP8UO0AJ+5ePbpACpXydvdfPh8PeNeNHlL8w1+6Co1X3yWPefdD3R6
rEROODuPUIkScZF35IxfMw+bQwKEJ+2Fajk/lDAnUpLWbzz0vSSLjH0uJhIo
98/qqG87Eh9r/SosK+f2yxSzyjZN8qA/HoSTOq1+NsBksOs5hDBHf++G9CZk
wwKfavtHzMiiUy541bskBmNzTW0qe91BOKRUNZa7B+Ql39zf6uW9ZK0i1xQs
TdpaLNscz8cmmOPJCd0hWahz7/rSx4yn/F5I87jsAHi3rre3Dkx3j8RoxCm8
2thF4F0bQ7z++84b+oSp/RnvODeKBRfwKlvEuPRTsq1q8EyRHmEVgVVvWQje
7+OUQyXBTw+A38d1UC8MQvdCpepyjyuU/MKkLspmw/BOTdwlD0KbZl4EYe6K
tvCFVuPzbk+TUJL9oRhM0lPh1MSJ1IiZ6q056RIz7eGN+v8YCAr6HGxVffCW
eO9gwfiIRmrth0L5FCQB9M5uG9NTH/3EzOHEr144f4gx+rK2qkmvI/AKAEhZ
XwoaA1rUMqMarjbvRLCy49gLvspC65o9EHxlwLp4msodrDI4zhZRaYPm3MVp
MR+x5gRvuILeUsFZfu895i8AQxyYH2S7VuAX89NC40KS/aYOdZH1+gFZBQhr
CMoZKZQN5yPjfjTB7RU1iA77m10TLQjg3FvXlyZn0QYwtzT+g8TInq70ffIe
mVRhtft2MEZN/Bji/iDiipV0kwHFagWwAmxpGinM/KIHwORTnqQRHSMCCM1Q
LgP5oLl+9+uJZdjD+X8X6xGG5wKeVZoe1+C/4tY8mf/dQtM5xf+62r0UFlD2
PbsGDtufwEKIbgJNyUt30Kv2M1/B3v6Ecu/OvtW3mITo8CjaV8cMD6rvbEmF
F4yPKggQtvtR/hgzrs5zCVMsE1FC153/2f+MgJ4oPOZLMW4TZJB0gduU5sSp
RYQFDHZPXSuj1/BqOBQtHX/J386pYGGSOxX0qJaSunzr9hkcB7R+EJsNtxJC
DYNOSXVIpfJYhJJS9Jd6QVCc7ejVrIAdL/0Cf+21+cYxf+fiBHJYIluIuW87
bXK0L31NxFI4GWpfaKJADJukKAA/dDT0F/kqI7fKCPe41JaUIbERndNOeVlw
KnNkR6axGbNRjoF+nAgyKNtMjRYB7Tc6opkJXwpS1omwxT4ay2g+uGwtpV/5
QYL+beI8KgnJhEQ6Vs7q+lbinov+vn63DnKGYSII4AAJ04gOz5mdLhYlRKY+
pARn6dC1lNDWg/dspIrVpwBnFBq3Ldy9WBWynZeY514O+6j9dcRTx8c03YRC
PGUlkk/s/55/uJy05XiRPnKAmaPVqS/QhI8J4q1Xg7Ru7UJgJuWTB6NT448+
9piUts69EIRTJbbg8HOgkzedxYkUnKbV+UuvErQa9eDoXBpf2tnhjPknmEG1
NejV1ep2eCzdmIKwSqUAa6/9f412zzZA4YaOQXQf08RmPWODJm2LMyOukiWA
VZ0ezdNtiXRDBsvEWSI9TEOoj8Y7at6/X9IrLlzREcFmVifx7vVA/iPVBkN+
KqQKN/OCSrryxudtctBIcOMyZRqUv4nukVPFtIb2hl/pfqYEaJEoCKhez3Dh
2rhLD7KZDoonvJrL7EVhWU2mOQbH9sdw+c9Bl8Pa/wNnWjX2bCTKn1CIpYPa
YcIlGSUgD5S3Zekfn6AN+oVwA1lH1E6KABBUHg3gwPUT5aTCl66/e52LKe0u
nsNRyIF+wI9gQ3oFXNlNNqjGvfi5w/hXDK3YJ2nM8Lk87IvOHXTOFP4Zo3wT
z8Dm3HWxGa53InMWW0RC+fE09tjw51QuEJpjwqIqNLl1lbjsTiKx9fsDADy/
VGAJ7h94XkafQngjAJhvKsv9Gn8Onb4+Z5paMlfZym9f5thVr5cN2ypkkgNq
FQTuanwqxdKo90GP9OV8owpC2dXKasr+DlPsoxsMdbFkYXShfz3lCc9ab9Z0
GRgDC0Ge68Sj28jy/RKKIAbtD/4k2otx8MSFuaAudwRm0clXrmWW4G88dkZH
t00grLDqjFPP4v7GKrjR+BK5QjmErQ97SRL7UNW9G8gvAEcbS+yQyOiPTrue
IKTzGfwpPlnL86Z9WyPGfTxAjMlPE+EPOaWiFKCNATVN4rxNkC00r4CMejUM
NVDIHrSundTFgHSj0wZHpGmSh5Di+M3T2SOAqLCPzcxYKE+6fNoC4qpknW8P
GNPZieVnpiuNol4brUemXtoUhtinww7gCJ4yhg1qgktaAJy3SEWhZt/SVqp+
eesUtUsdgW+e5KuOwZnpwFyJSbwd6OMSGeyVEeLqKIiP0R1G5sEK9t2IgwzF
YCZxa59QZHrPTtVjPvGomwdtlLgg/y7/zHOuKo0OuL0YXglyQDLyPXeZbkph
b0vBdVED/zSW4S210WlC8i4wEGwrffvjX20m1wT+f9sx6cxYIqzIp9M6MO2n
8hKM+I4FcxhIxYGlqWr7CuDwmnKILBndMXnDADIA4Uwq6TlMMqWcQjr9Uex7
Z/vyZvhKFg7vSyL/7A4ADYiKbvSHVgc+FOamUBRDEm2wQM2RhE93vuafLCPr
HRGr3CrmFpRCSyVcTJpBgrsSUjqaqI6Pmi2OaxpFrdl9TC8ITTDNmNPXrHXW
cppwmEr0cbVC0Hbz4b+WUvHOLtu1hQ9S0Qlcrpl3UdiIatb3Bmr4EWGU4XSt
JGQpTnZcfB8W+joLR2Lx0j9kZCtYqm4GBuKF9XW8kbkt6dLvhz/BUHw6tvob
4orJJzkrX4iGTk2oDrF3UxKECDQHjJ5Tjfpb5ty4wnq93QT+Uz7a4/Yu37jo
H+Oti8glr5nFIgGSjLscsE8jCISQITar881iAdDkbfutbLfF5rPIl2qJpATp
vWlLEhDdKZi/ki8ma5RTISVyUZDBzaYSkHWGdkL4gN0DJQ8bPFx3GyqmfwhG
Q+dKU1CvCML5MN58Dlwr7lgD/CiKBG5vgtWogvfFsjg3TNXshrJysSBU5zN3
XFT4GZ8AxyUt5DYQWMTJcQar8cROR/pqCYvwPf1lbdRc7XhIPhGja0zpAxHv
Wmijtf5MK5FjalxulcUAbhLQU31StAcRO6B6gcSSbu+7QO49ox704B6DARwm
HTBdqV6US2us1I6PlqU9p46xWbj/hbgHq4fRBX/wFHbOHNzmtziEpuIBHbPY
BwK8tCxy4Usc6XJBQPvJ/yxv9mfnQj9dYzELev8gvLGvupNEUFgWTeYgZR6H
5/d+71jqAGDnhQZhTH1W+sg8IH3bnu9LWrukVtuYlY9O+WOcj1ukQK7Wx2YX
N78Ff/tH/Vzm34Ajzjslcr/Rm7GA9mWKcsE4Qh4SeJ0qhuWncgRvsalGpUb+
L4Pp9YMYUcedwj8Rho6aL5ieSObTMYeMRcNzkgj3Gf//cWDdPmcY4Xh9HrV3
7c4fnYvLH2ITdcJpcELwDIqJbH6MM42vRYj7KdM9KuarEdpGkR7e3MJNBsyt
NtQD8840m/vBeRDZtSDExP/HYm8qsyhF6OpZJfjT0j+GFfViu0bJ54wR9IOJ
1uG9zAYbyRjS0NHAj2oW30Ah2X7RA3LvttrZSqEJlp5qcIah/EAL7uTX5TeU
jny9ndPOOUhKZWmEOmrN1YKFUVPpNMaBS+VXxktMV4hF2Ksl0jgCSkDDGnAF
dQZJF79SULBeZ/R2YRaM+Lmzy+04yfqM/Zd3gXX8I57fJGTYH9rvpPEeakih
lgNSohe8+4Yiur0YMtgFkCP73o7RpFT5sAG3d7g02XQd6n2ljKEEGyY3wxAU
U0dIHy8Hdu0CRa0vgFOKKRNTkQKb9JO8XhU4fPRhtjITOcMg08LwJ65iPS08
GphXEw2p+O+sDN0RQpF2rOhjPXjry2uTaw7dw7ChsYFGKHqbmv32E6lDD1As
puy6dIhCJWkHpDygUrKNYjZqVKykz/pid9QITHXHcw0XfCBp4w7+cngPYnFz
59J6Xjgdv481OdP243m8ofwSihMhZOR/rG7jkWGBJugaxGt07GFcooWTZ4Ad
iUzMfHjAvDLpbfVZK/m5ZxmK8Zu1SSeBn31fs2o9Q6dCLcMdxIz3NuRs4qqG
/pbfz9TFsjv08Fae8y7ReIlTqd6gQShMyIlKtcvHJj2JWQu5aSI5A6A0RvMB
me2ZdQuQOr5MQ/UD+vsFgTI+UT4FjBjGlvgxecPyCvxBl1edyA7b2vHvAZ0G
MCerku+MNtULIBmXHeNUmRW0JIInh7JcMPB0AZGryrh7CInTSqUrzq4WnPPP
MHkyX1v+K9Dzt1rz7Jz+AmMubQ7a2Xr2xjwPTFA2F3RmsAgcgOuJIz2aQC0H
pfQyeOoyo89GyhWiq+KwcGHNh/9zIt4a4B1h9Txg8HLhEs71ZHElPkiWcnCh
THvlhUtd4eW3k7lBNq8JpenMYlphosjesoUqSCYDyJRZMfMI52NgsxtBlgPt
sQhgcXrR7HSeOFP6g97e35Tcg76coNnhemmJIUSUf3IgQIE9Oapc8tG8fNR/
a/n+T2amuTzhoOFveuxgr2RJvth6JRoR99e4B4N4Ys/6ZR1FPFPjQT3tinqs
I9aKHwSQZce5NofEzxSpsYYMNnq/Y2lXz/5C7J7JTYDbn7r+226BfJg9G9PD
4wccg+f8JTYt9DzgeQC14L7N+NQSQjaFvQ6rHh+uUvLANnwTXh24qhXTdAfm
5UKOu3hJiZr++IGziF54VaFp9U0f5GrxfSSKSOdhd6Blgkx9GmLmqL2vXnix
KUPMCxJ8A9kr3m2/SW5FPvO5JKoaYwiKzYaGhTfukbMyhyKqhmjuPst8Bxeo
/eR1XKTTQbddpahJxftoE5TuMuelnzU20BwdgLxLe6TR4Xon+EwzUklBCj2D
zZ1L2+6hiLokdcFo23sdCmVC+rWiac3KD8ammTxC/nddmz5Tk47UUsRahYVY
TeUy8KMCJwalNkmJSIT+WiWTj8Y/0pmChf/CiPsKqe4uyQeHjRLdFamDK20v
vP2TgzEwtj9fcpQbnl2i4jSQUts7Wfp5qXLuZysDP8YwiC2QUgdtnuh0musf
b0SUL1eut2htCRnT+PKaCVw9ywHK4YmjuHFEOM2xoBDqqT38mx6TDVXaoH0h
2SR6o+iVgoRGdrndk7mKukfvOk5gAQrg09K4EFZD51BW4d5IxQaPCisHdToc
ukPNyFvMkR4eesS/Se8r9a5eNRivOpaPJBH+aHfe4PcYyHyv/+WI5x8NPVzQ
GRMxmYdQHbLPm0HfvKeu1fmeIkOCFzjjvugvrA7pYV5v1msenEaE4HoUNfo3
RehqJWwAidizYEbQsmnCdE+BO/dTRqzcUuFfRHFE6VTbbWR08/xAxFsjBo6X
NBqZcZrACT5zBK09jHcnDldEU6uadQeZV1xgD0kwEM/vmt10uY8tOCe1g4L/
lBIX7NzBM8FXZV71WtdGeHAUqxOiQEjW/syvgPPuIHXaOBsObcMcnNd/DaKd
DbX9AYo4Gj2BgiR3UwKfKe/mgYFx+D8vRuI4mqjNo4nk/VISVRjr+XuPe+Q5
F2RVA851M/CJibEdGGllN0bhDRRO644QXAz/vZi472mH/eiMnKJ6X5ZFfzir
stocprL768/fMAhbME4C6U5L6zQNZcp7gLtBSgPpTnfyO61hp+g1AFmm1Usu
BzaCqaAQTKydkjhumKMizgQ9InDiHb28ZhVU+JmDy+bDed7wG0ctaDv6S4LT
MH6asTFC+fm3i2DAHjb/f0fqYGBMluFZcl8ZPNarngfMCjvwXZhj3KVAfynh
KmAHEMSp98dXI0Z3qmD5IeGOa1EQZoAw1Iti5/dK2SDIZbbwgSu9ePD06+2H
usc5HK2UOQsdlRV47CdGyBzH5iz98C+fVLVCvWqm5wZ0qmIcULygEH55zKFi
7Fel1PYinmaR/pdCAa/AGmmcYiSLa3fUNcNuQHF8EONC5pnGeH4IhRFlZkZY
DIS++4CixI5JabUkDmItg7ei/x5E1rDYc+xaP/56zaSEwhenF731wG8GmirD
5VXCu6bDCfIgb9w1xJvl+ky/uSwETP9+7mcDCwTKMceuya6NvbqjCRMGSrRs
gb0O9cnQrMQzOvoYlXdhO/a9ZPZLk+PBam3ig3SmLVvJA6PPME3K3UECZwcN
JHU0IDfniM0Y3uTg/Ra4BT+y4U5K+h0tmCOeh4HZMeiowwkSN3yyN6UoVjLN
gjcft6Z0yctwNTlC+Tn54wSommFmlfIohl9iAEllkNU5P9s6LsUKKSwKYyEv
4ubztloYRkvPrB0i8Pj+od74vh4OzSkWHEpSa/yqbaZ6fsqIuuqOkJLopahB
ayxG7bffo1QrUCi5bVirGE2TB2eDv3H6cd0nvIPTBwuk0lGRf471yR3s0bVe
44cCF8D66EHC/MvlG+9wT6sxle0OGjlFVyhuqPiIUVCbZ8jfnsH2NipioyzR
+5mj7HxCbUr6L7I4E/rkmxULBro9gBy0O3i5Om5IGS9x85Yc8C55mmYVryUW
e61fJ189Nz8wtwl1luGa5QQx54dTZNybgR4XgrMurnrNm+f5p4tRUbzJEWyf
gqK+GamsYJj/pFzTKz1VIdyIgn9UAfjlf1Gv3ul6Cf2zl6ppj+1UMg950va2
taZiWQ9tV2y8uqPObj9Czkow4wH/g51gf5dIFAv0/JZsb24Y2Wm+35Ol6poI
9uyQ6Rpz12N2pOoEdMT+AM/FZ/ChYSN/dNzNIwMjzESrg/LLm+atFeTzcTT1
X8LXIrDrYhy71AqFwh6AZcMjXH0vEiKAcN5q5f5QkrLFs4acdkKbvaNoUD4P
vsSEGXgEwSkiZlHt8y2iU2vsi8qqXr+P3oPWEap9HT51U6vH4P43P1s0gjCF
m2zqpMj/M5Xfzpr/yGY1i7OF7YUNJpz5c3Vp74BrO9VzQed8RzhSVwFXm8LG
DgiZnOBzo7ABDHkmFHpO4RGq89sFJRPCyvknnHbRFVorLrtAiZMC4xEM1Sd1
NFjKzIbyiuCvHsjXTr0mm7gnQLeipdx/H7dVvDn9z+P604MomMEG+3XTYYZ5
TCBgz89b7TihSXRuHlpZrDIYP4htuB31334VZOO4+m+Ce9gQYo6tB57lbBn6
3QN1+y+mUsh4w8VPIrHw0o8GXJqQI726yHvI1HrUI5y54MWMzovYzd8CkyRR
mcbirbxtnDZce496LLQ3p4Q6ft71fW+XN0PKWOXTvk/KJNUKqDEnRr1anUGb
Wd+CCFo4v+QAg1gWUzg+PduxprUt854Oh+hUCUtLEilkX8eNAXWI2RMbISo0
c6yxxWpsC3KZ2dUbJdUkv1Q8QFdJRAjPK5NteWgZfN3Lt1AIN991DagqR+Ic
Y7zJxPJtJwKFCHvVvFEaGLkwYx4MT9Q5Sx3ZnCF5N01lvk63uEnPxC4wipnr
QwYqBpjlwKa5/BKzaLBJKjbborpEwCtiutBYrHcNz33EYwiwRriamVZCTYkY
8MsaH+t1pxp1gYhX3iqPGBF65uaeN9r38JmkLoDUMS6+MjNm2w+cTE/5kkwi
NWM7Dt5gjONUL7UJGOFc4Z4jciIJscb0GeuKxEEbgw5dSZPahuggub8RPvmf
NQtdaqmdr2xyHQbP6rveNlV6NjbHsriubtHtidur7O0MJgU4Zp2vSSPyTAEB
kYGHfBdInscUQqhv/57kxKiUapZHZjA8TiHe/I8vDIosslPHNpGj6ROPBM/O
meh2+ZnWJy2cRbxpeWEYmHHy2NTutQ+r3fjk7O6xKkZTL3yHSzfhW/OfXf5E
UmACyO4tYi+M63GyVfjGXbg9CC3IPY8BxJK6evFitn6LudeW2qph8EzNwjgB
/T0sQYPs87pHJfAiDpEJceK6itcKKYemnEbgYN/4ZbxfFn7HJofclRsGytRA
s/hEoj1jdyS/eL9x1ZJ5Q6VGEcXhWmk8Kt7clF0j4Wl9ZA3BuZDLiGh8skT8
PjPSTfPQ+wuvCIA2nYUphTaPiF2hzooPdiwbq9qzuJqq7HUVojYDpxjvJOpN
KdVL09xeg4orvXUMWPfsvKD8rUBXHKyKDF0/PNzeYbOMIEpkiVG0K5TXscjv
RstdUckVr75psjWTZ2A9uFULQdOkxpZmAcZ8lqhPD2L8Zr2gONtJ0T7AwGKW
jZbfbuGAhIfpwytnp/9TK1D7IgsKRAvq9t//+G52XQHXwy5q3YLtVINeIf2q
X2AOq2nb/tCG4RTu7A2xIpIEJx45UiiYHgbqLrS30ShZRmBhhwf2ocjTkw+S
zxEEYbNOFUvVGS4sfIK/WZQWDJum8bDbyfSWFb3Prl30mVhn8FP+M2qZFYVZ
6X9Lq/6nJ4uDtaiE/ZzGNTVHEZ4EcCC/OfLhfmo5lNX44yY1Em20xPrY+3gM
saD+joWecypOdROFmdtjIS8S7rRqdnS2WCYuAU3RsbM+L34mTA27cAX5tn1W
7kIM85gnl59R5ky8zw7pRpuPf3Wluyask+16F3wvecoCFziLGu+S+9GoZQG7
pss+k0zkM8ClnS+aX7EYJ7o8GpR5yIoxO3uHgryXYOILN/vx6sRcrbc9kVaD
awbB8J2NUySQ0VUw2JbRsDsjafdcZjTqoP72g3v9fCZH88z1onsXkbsCH3ZO
vaXze6QfIynrIPRFWe6ZDVxfQtXWPMuh15ff8Z6DWivMSdgeMr4c1ZuSkBw0
xxaJdbODoO2QqJl4jlcZF4u5b/BMhzYwkykRZyTqB64D7OkSm3C7EmH8otzc
ZtvtvBk4S0afMt+bNo5R44vyufzEApasBcPeJHCi4DJ8hSF4xH4LvDJF1aEB
3ONI2wUfRoWpbbn203mH9xhPIq+dJaV+/xUMvC7I8H8BfKa3mnFqMREQBt38
D6871AVLoF7HMKY92coiN7v6RaGZyO16KQmeWSFYe4MT+P9kIjQz63uGRqfI
tZGGZuTst/9t9gqAU6isoXEDNZgNTxX0QBa17QAkGF+ghCp9owT8Utw8snXP
G/hcoAfyJI2IXGIQd2CpsfuzMwTxVCR6lHdkk3C21+Y5blDWxxvpZx/TlzY/
S0aswrtb3dfYMP/YQwjZNfF0aYklC3vZHVUG/CY4qQE131NhQzJycPeFdv35
7VNi3H1lwngoJeGVNKHe/W6GGMc4K0zUzjID1QGv0Ke0vwY2Fm90rwtAil0W
UcGI6hhjylKlq+PdMFsDlf5OFVXu5UssTN/VEQQtzLyFoNYTazIPh4MjrKJh
95bq2C3AmsdzTgLfKomMnYJOXD6IWUUmX5Nno+Tz5+T3s/zDYzSAqXgvGV8z
+u20TH+Zjk8fify9WHuy7Bq6YymXbQoSI8KzjbqElNBoOzDNr+4DdjV7YTbp
gz2Dp3jqy+qhfik6JR4wcQuSFQjZf8BPmelhpEW3rFo3u9Lr+XF78dg5Zpgt
E/bh4j1IohOY2wtof33MsTp/y6n84t9eei/LjCTtXnGyObQFSud3jXEkn3c3
NnyWc00qX0hSsNO1rcjK0ALgYFFNNEcAxHDLlcsC6UHN0yDnhV67928bDYYq
ZW5IzU2J8G3TAoFuXBkrI8fSdaJJ7XHJd3AxibMAuKXXrR+0YcYVTbdu0+aq
ZkZtP7c7vQMYfAI8vH/r4247FVUjlkb8cdDA3Jqvs0bHJVHH9gaCekqgX9Oa
9Wo9pqGH6255KA13emM0sDQz8Xlk4sHKO/pi6sFmG30PaPiqvbUDHCV8IZoX
Qx/BHF3bkREaHixVDF3ZmS4rvX8I9JjxVKL1zbZtk2ygbrQCTp7XfukuByqD
orc+r8MmUSwPpmwSkg99wepaAoDyDFOfaCEbTMp1/DJXyeUl92JxdEIvzMWe
bGytv7swjdgw9J98dh8lrWkL4pClTXM7bT68NFrkhRoR2iVBBLC7e9EzFU4Y
w/LhQztmXvoC+WWqZ4axHzPC58qEMHGmjeRwzAiqKOBSfnv4989qglZfMZLt
mElRKPK7FVVgXf6991WwMtXWYeVKSHt2LtmGKkTgmTEkWN8YqYeGA9u5hQhI
+HUhwvKL9IqvXIBnPWdFhVP/aMGh6A1j6W+5lkX1rWJCZjogxQrl6iuRbkxm
LBkC+0LLSsvJPQ8rY4ZEZ5utrZAGUzpAb46PBsZnDznppVxH66/zR9L8ovcf
yOoGf8qpZYgO/yhRdEz+uRuDg2S/6RyZLCCeUJ55UorxfbmE6uartGdJz+I2
b7T81/EGHdWXucgAC+DZPZUNnscNqqQR7Tz3vKho3oPlZzfKpOmWjKh86k8n
seEH/BejKJN/hVRPVCMU3A/Sj4Ivo+T8isDsLnb0diEMB3T7BW0Igm0OXaGO
Wf9iSp8ekKBVE7zvcokjNSuY2u34St6wp8GKAKHZPwLsxOJqpG7JAeKDUq1E
s8QyPsAdZC9jojY6YyaeSexGHRqTWvdTO00ZWJNWdgIUH9BTjraWh1o7D2c0
JhDinhiDWRaDjjR77e2tQwrRMlIjuX3hmdJv2FI2RCPbN4HVrh4+lNtOU2+/
lAl3CUFvnjtntsstAnKjQ9LSl7DP4CQJ/FdCjrU3wUFyW3qMkPXRbARrtA0U
oVcuai8a2Av1ClX1l7A+1cEfZQWnbL2xPKdusIGLqufn7FJcp13Ko/ekylkf
OdOFG5e3N4qroBfM+esM0gO8Q9haaIIfb3fQ2766K5tonlvfH8vFfbRQIW86
n6en92wkbrRJwniFtRk81YPJ01Dpw13jfwdJ5+Co1VI1YtcZSgTSUlWj2Uus
knxhgPqDtY6AhRhV/TyPakipbewYzW23GyyJ2buCXU5+E6RGR4DL+uNA8twX
CdVBrFLqiPesBpVn+iOLUDvb+rCKGAuZ0WbS4q0uj0XDO+FGdlFXB60diOv4
LY1XqYnod/e4lbS5b+Zz21tIsRX4v4O8cUy9+e5c9wI0149j6lDQXc8ogFv2
514uiFHeGP19NYP/VuHuw+OrZd144m9xCqmIzrLNG7imbxogvM7fKaHkpM4U
qynvSV72CY22pgfioLAvntIi4yZQvgTmDQAnAZNGYaJu3kkFfI9HXXcYu0AP
k/gRNkKMMjuOFlobN6FNCAUAiluAnLW2p0yb4f0s4UfLkQsg6IJRE+G0AR6q
wqGqhI5QaZXlQQ+JPjJVhwxukMoDbmv5hGuNVhF1MQ2hWJW8C/ooHoTF7jYe
mtVr9FMQWF9Pgh26G42Hd9+C/nOPZY5AmanDyjrfrehxGoJ2sbWbMiIib/cY
2VUPh/4nwGTXbgW2g6YKiG1KsgCfPmk8jkl1EtnwPXl5Ctl15JErb6rzVYBB
mRgIG82thKKiYvlIkyyimrD9iE7pfsKkU0Mm99a1b3m80nq8B3MGm6TDwIKL
vmzy6tpXyhQppUAgqKPeSVVrO5gKD/5EGcFlsrr/KxHiIIHFqKWNL16u4Gya
DpRPXgY4SFyC7S2fVQ48Hk070/YoWnB8NwRTo6Ck+9rn4s2vD1LhwPp21tmL
CSOD34WCvj/UNjiWmYKU1CjaGrwWRxcY5qFwDYwmG3p+oTUWX7IuuegMQnPM
OlUH0ogdbti3r8G4jl7RKG8ERTqRhp9/bi6BXh/1z/kaNs5KRUxUNaE+1BUL
3Xqc8fDF/3g00ahNk+qVf28b0CvITEv6pUdGaWi8UL4K0NPppG2iWfF+0VT3
Jai0AjVxOcaE9pvxDFNChL5RF0guhViBX1psjMnlv0EP1Q22xAXxw6GhXALC
EqKT5VlN4ViTTqE79SsGb4Y2+kg/yml4Z+oMzccH+HREFiq+pzzXTk8HkL+U
LzIp9Xg1Vzv+NsCI2HP9luFEsbnKFJ+6dgyuy1n+oyDow6o4D9G/EUx1JD1F
XNbuzNH10OALv7AJ9UrrGJ/AzWk0Dy5/Opf/wnHt1xaaJx0R9ldH9nKK+Akf
ADcFcZYvxIb8nWT7F/zI4D1md6nju4kE/CAJiXnUabg6vuuBkmUoIs0SXOS2
+xM2X1qZnNNmbJZn341pQaabqXORbctHubRxz1QsrlL5PFvIvA0Gd614OLbv
6UxdgkdA6proMjqYT0o8gUMtKAA8SQ1zRYq/0TSh7Xt7KbMATCxyrJXJ+Cay
0eLIRWVR7dlCmnTPCvc1jVWxbjAgfEyD8HqzRJk1kWHtVuJK3y2TKycuBhsy
vjo5TFtEC3BtHU8yjBC6/QvAijLGAOMnsfMAl7tNwiNL0dAQjTfmiEZaojsL
Fxmnxb02yGN9JPAVBPVtJgcjKZf6lOvcveQeL5hogtrKN5I00xjtwTsQYvQN
DZjHHHNod2sDi14wuyAGIHivfaBGq8PkYaNPFZuSNFcPxQYdWoLjG1r/5WVO
PBzsRajDQhbhbQ6IoaEwCqp83G8vVVaEJIuDpuo0a3i7lOVWLT8ltmmmeyX+
6N9f5T2I16qXTP5aq7W7fQcwsuLSGrgh7PRxkOsFKzj41X0kOdR7ASY/AkWK
sz8CjtqZH2AGOrTxumm1kS+vAsCQr0MDRK/1UJxn4XOnZIyfdORSgX+5/6rX
6jtNUnKiM0n+MBY1cixa/GVm9TM4UYjEy4+h2NmHSP9+UuEOvBswdT8d2DPV
lHXas9OpzMlOcNfYXTOfTqtUHz8m1Ropro73DVUbga2NMsi6PL5ejAtyxbjb
x8/rGzfROGUZ+Qyxo3sChKqxK1zXnQ5DfKIYBV0bAeaKvxzRBoQVmebx50MY
nbjsjC6s3it9M7hyMkWD22SCeUMOv0GqA3LqFgZuGHN1b3DqX3nsMy1KlQNv
uSuBwAtOEqZ48VK/rgtmDHnVPJDCybJ/jGttlwhFYVOTJjBbo2RTB95J22UZ
plsDiOZqAb0EZB1RlGn5UniSmJ4GOIRPNwAJ/hBpb3gPql1Jgtu5gqU/r1Xd
XiOANjP6yQoZDUIpGmromRtdO/18txux8HEJP1ZecsT5GqYw6F+u3i02DcbA
OIXzKxCyFVPbMINqLVl14P7X20Mldm9X6vQCafa7ETTWDquP2+bBAFc92Jlh
FKlOpl0VyT2XLEL8Z5KvUTjATHBfGgFYiF7/fr0WEP8ZgDs0UjVHY5crbyLc
YM04admNrdKHQnHTgdHufob2rik/d940I6xDprkMvlJaK2O8bb4e5ReZkONY
on29Utk34uDZnO6uXF5NlGwQw335LotOkyR/S3LnDPYc71f+cyHyjOc0Wdms
Lwb8InRNrWTG+ygmPWw6fc/u2Off/w1egwDk786pCH8XuAyUtDWjwNVT8jGI
HJg9SwT1npyhGFAzccva7g4D+nGl5oiVdH0uETrxJJUUz5lo4AxH1FpOBdJA
VE9lWy+gdv6PxwUWxyIyG7+zrcl2Z9hlHWz1NjNYkzcAcjRChU1djPFWJr08
jitqGsOEQcfLEMlEbFLB7OyannimWgQwnU7b1Td9sj/g4H/Jt+O/daj7F6fL
WwBG4CIgTSId/RDUwxoex4V5U6DY2L3v/wMKZVlskimkEZ3WWzzb6HRmXdtI
x8yJrtLApmYvW/MUIGUEdm2Jwc8t+xuPYxNP1DSbKfCmzIErGYAvM75Bz6QO
QczAlxyt9aQu27OXoGVHGfN/MjpAMTqaeOc1Vuz9/ta1yHxRcUVaRWoqdt6+
0cktSrZAYlcivpS752f++0ntOv7xteO5WXCtW2heswVQMgZvQwxhhEnl2U3A
DWv3f0cQMwpjCDGY/krZ9PTfeshVauw32F9o0UP+huAAf99pC2UJ1k2ApfQM
4XKAoHA74XTSbYqzfypfiHjTho7087zjjD8KsU2q2/ArFd9dM4Ds4tRACb4u
0rR3wbReSSdItf2Nt0Q+K+aw+VVZl7gHrrW4e+K1hk2xgRwiEgUOstU6+Pco
WtrP7wn5oS8o0r7shIJS135BcrNu0VRxEg+tv5pqjfZ9U9nL3EDyWeYmUFDg
hVzcgUZozwHqd04bGo0WH2AMROs2QHk9NtIYZgnOeA2ehZmt9rvxBOMpqgDM
XjJC4AyQuNrveYbmyXFoWk7AXkbCh0ayfnCnsVMu4Tq/92cMhjBRfRBfNL5W
nq71xiXt0YtA1ri0HzK7qTmOY4Ek3uEEmiLOd5KKGuqtGAjrrv3O9i82ENS9
Z/UpkHq4I1Um269CZ+mV7rnlbuuuguKfm2V+IHHM3KpWXsclcb5I3rePtkaa
P7343/iPiIXbNo2I3J77Q7TYK72lUGof+fI2bmxu4heMYzCq2npkYi7w4qRB
JRF7QBPryGfH/gwp54bq+dRsSc/MZVnZ+2/1ikxSd4TuWHMxKVU4yua9ifzr
+AFJezDHOfmIk0IVZ9MY85CunbkEPHdKc1zMX13WL8twxUYnBdpdqjGKSCr3
vrac6bwoCqDsKpe2B/E8cZdfPm6D9W0Ut0sswkMMVdWsaHLrlFobDsZSvh9j
enp35BGdyJs0grDpeoeCHOtaKxo7kNIh1Oc8sf1EhU1z4I2v+1skuhCQXujv
0MhILFzU8GwPuTHFxzW4jwWIRBS6nSsqCQrQxvfHU35w21/npIMh8ixzYoy6
6/kTUYES5ayhHZ+hMFtveGk7uQNPl8bQ4p3b3pMBcW7jb71jv3ugLWtaG1CL
3+92gOF9eppDWwaMuZs7i8aO5YWqNtGYgm5jlLoDD0CX9wV5krovRJEq1JIg
q+IrxyCQweURdcZhiZhiQPqhj6XsNPu8BynDagMooPQfxdsPSiKxTxJKVDty
ngCUNLrIvik0K2HS1YGgyE2eBUBei5X8ns3K6WO0T+s95kIn8OXywOl6dgmm
n9xeSuUKhRZReEzhWmkxuHasAY/aLrPFJyLh0v75C+o2hl4F0NkAkuZBCXF6
47hnpmT5ZagA+ItgxZtGeuM6KeWDSGek2Ftg4GrVSTuLaDZwtfml9jrHTDkm
tfiAR0LWpSy0jOKWFMT3NpX3V+PM5wtCLoyXq/fXkq+Clt9hetMso7HQSDLL
lYSWbCk3WoDxP6JX1JR8hp/ptcvdKp5GNEqbbl63fryZtLFtAZxV2nyQDPh3
klUMx9Q/a4WMBn+Gj1EAjPHCMYGid8/aGmrPxVo7YCdxVdzOkSNmegnHqnAy
jsPAdMPL6yIQMbZj+7lqFBeUXzzPdPBSpGQSrmGo9TOlgn2SBJ+sovI5AozP
9FnL2zC5yUPQJdFfLHAMq+Xjet8iFURc1YPvxjepE2Ah2Eu/qbWe1h3Pa2sp
Cryb1MUeh6AcS7w9Td32MsmWU26uYIzHKjsuK4p1tvO+cacHXBpfZ5dPGsDR
JpS1aETAtCTtQgw4f/fJUb22GOgcRnxFEsdIYrMUYQLvgKVxpLXIXR5oD0vV
3bWQSaUFlac0IELp5Sj1X00BuIW9MCAVcq3S4agwqPLbUBLp58G4wtQNfbZn
ryZZGDAOksCGRAv3E5BOdgJnQ1X9vM23DfXVNmnA9XE1e8aoWe1OT5evOY07
y1lT+g70zD6Dt/JeGq7pTkKA2Dsp0xtvIfe3RWi8S98p2p0SnXE/P6qft6AM
vB+bqGZewuCT75MzxzPE5g2Y2E2Z1LIECqYx7/lMaeAif+vRTjxNMCoLnlZr
X9oeAl1Yum2Bbm4v8FZ9hDBDNZFoZeQLW4ev69oHYqnwm8ZZoLkvgSiwZkpk
bAVnIrf2MD6NuSep4MS/a/wx3H/sQ0VLcQYQ9ex+7M3yjxEm0W4WVR4AxHVA
/tk9fj2QepI0JuzAo0oDKOCd3ciVlHmlqbVZGPebbfbKd6i6XWRF/drZ2Zo3
0WEX5SCtHrKTqsRMFyjPJsrS9Hk5MADsi/AhjjcCW0wpIADy5lDc7Tu+u8gB
ccnPCj1Qm08jLutS4e+vMMBiVolvZMjoSrwfx8/YYMXNT3nErQnFvSudh/5s
q9JU+I4ZAMbOYElm2roQK4nuxe4HnqcS+BBdhjPIUppqW0yzALiUQlg/aXay
fRbDdy+38qL876ymYUhSIHyRigMVsAOU/agXmdtYtZU7h2DlHStJtTFq6nTD
JWaUOUSwi2R/+rGwSQZIjhj5xm/fa03fCCuz/on4kHef4Np6N9sxyRgs9+/p
hz5vJn5lygyTISSbRKTFeLjFm8bX5XWdFND/gvYfpv99WECdCY+KtGy3gOYl
OxbRhyLZb8W28vMgpHEGpZ7Iw8U0D+9ajY9LZ7DvNu6IyLxPhKPePBvtZioo
JGgZGndrbbSG2Bh2IQ6UW7n83UNnuteE0Ne00+9uIf/vlHQ0Mm5rQPZb8pWG
SEz6JtMaFd3EncGLVj78cqhX/H1/SVtVkUPkcJtBAwqdOgDo0vTltByIh7KT
gRW1TV69hCwnQqUS3QA9dwFXZ2FJtDXijpx2SLcE9+A3G2womQ2cjp5Cs2Xq
ojtg9lVk2r9Hd7P7OrgE70KRrqjD+IBIPklY8Ftq/14F50Pd0bt8f20PYvjb
y/thwELr76WNHnAWClIlL4NiGBxOB81wnVbO1Zsa7uPEaFIFr/b2FJM4L+Ky
E5dzHwJFWKMxBgrmpjWbVBNMfYS6NeeANUeDCVp1Lnptp7QC2g6vafuEt0K0
hKCVBJtyIJGzA33dIMQNBYEA3JBHZX8gz2Wmp4IST+myL6KJwPBdvyACFlaP
+gXNW2BP5UAZgrm3b+BEQiBbti4L3iACRnQ7pWsmEzio/04lCgU1vHOJwbWN
GiqNw8hVdUWyWBAcfz9m4TOZ4CiDeSN0//ePpiCVSX7ITrr47DPzIdI53MpA
PP7vJIu+9CCxyT6rOJoX9iDXyc4Z79OhJZNktY6t0xGwE2kRi5K0hQoFl6nS
HJlQDU69UWoez+34zlrWLqZjF+N4xSt6NoPTzy79m39to0CcotSiBjZSkYd8
3QNRUqcIO7yr4oQ4BYqW8EGqW0fRQtQphAscE35ZruOqJscEK5N6qgSanVpU
Q0UZOcqImPw8KsadtIsWv2z1eSTPVc6PvEM3ZEGrA3CQBr8b5xCWl3vUyNG5
AqwF/lSzFdCTyF7rtxDgSuiT9/Ew19sdtnz2NExGzBqhPft2hPk5mXxqO53J
VTeo5bXwgEAel743NGcTiya3nyz3p4ny5h4hthEAoX3XlxT7gKvIR6eFuM4x
PwofrqsqK2QXfctEeOnVH70WDglMUQ6LtSzjrGZimmcfP4Eail37tYD8U/Gm
o/H7JNIAKSkInEKH22PTwoezHkb2Lh259LyS1DDm+bDSZ1u5vHMxKFDQTYIM
/OA1ec2EU8jfXvZvlifGm1F+ea0uhb5gEOcf3h604eIbMkMyFK2CH/JD8nJG
Z9TyIgg8tgV5mQI85288L/O7JJ744ZJjt+jNehpC8QpZSoFGoGlzi2/rLjgO
BDDgNXdNLjs+WZU5eCLirS0wYTj6KXYx+calWSYl13d6BlJCrAjuF4/hXn8c
ITKOhWDa0joHDdGmpjkZrwLy2csDGKZahrHu+k3kuLh6HTLjpHRhRzRLsScN
X8iCf9OnNwtPhDkSvSjvf6en8uzeYq7l0ALOgAuGWUfXESB+jGmEzwEdI0Q5
NvVAVx1funMevpnPl0uCjSMVruPIfowczoQ1SCFCW7cPDcJtH0Ga3v2geiJp
+g78Bl7IPsYteQT/8sfwB0i6jhb/pxNwgFsCxn3Wpip7j4imgs6zRguTlrBZ
qF88XyIQ9GoesJTyIpar4Lj2LMCA2pjp+nAmNy87XEqEQpzw3+TkKTq1vgou
2uJoA6x/1I/hbO2dguKh8jm4pyKyKMmZqIpwqbKhWBCUGmJwBLuKDv3qfq6j
VufgjZVHuNVQrXk4qxFhP4YYA0hHjZJLSxX6xrIj5giiyU8D9GZWDNw786Qj
RjQyGUUuRSa3LEdm1Mrb32Ztue+VFFYELOKWH6zOz6BmFH+znD44p7jWvQRk
m5DX4mPXS4/fko67ZKehq7MhyFXjeVpxxfLpSkNVvNgN9DgVDrdUzu2lVv3C
cP6thZROklncNTNuzvTfuogdsks5sIlgiSGJNhyCSVH8s3gFNDP8lWmSvirN
1zuP49GCN9nwtAfTHB/Ku99OLWKYZsj5ZEb8328fh28emS9Zu8b0tyNvXzte
//+4XLU6gzh5dVVxaGv3lJMw9P8z8QKrXWyuiPNXk1jKh6LHm/CdZarGnh5T
84fnjeFRD2/I/w1Q7JRv+AP2BxhorL59HQpBu3ZnQwLRkGE6pybG3WcNpUqJ
/lv5iSuS1vriJu/8dpBQ7shkflsyTMgHzNEoq/e/ICkHKxSRPaSkxotaX7LG
ve7HfGM72jN3vxmlyHtD00JR46SckiuZlSsv/N2CKJqq+AFJK1j7jIv8MikV
2ing0XOGN1f/2jMD+76SK7UiqTEuHtaGFeAvWPWZA380GA3/zsrSH3MdBuTf
W3Y+7S78cfRSB4/V9776P1l1Q4dhgzIoxYcDWDIS3f/q/2UZpS8/GHBjw08z
lhWRn1QZJSjagxH9W2856CHCgwI9sMQNhwhPRo6YemTwwIRnLa80/B9ex2if
jYBOUozEcqnxyepAZ7IJZakBEIG7hsSHkdLa

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpejgwxE+Cxz2nPNk/Myqu9lmo6VEWW2v56+9Q4h5EMmloL+TGrFqsS0rzXK29+2wx3bOF3olqSVSY8JEw2/z2NFiMmFbRgC8pZdO3dvYvaYI0/biVCOsqtAroX+wdAniDUSoJIEbZpyVtwPbIEqXtoq4LZ0rK4w6uvrt9UAF+nWOEQ2d0OpC6w0vhLGUz8tm58XUPCV1R43P8LtukC90qZXxCxroOmRedXGuPTDAcxIGdd4lfLTdXMb1pZnJDpS6+5mRTsICwvrjwqvhOJ1VRoN1DiNi2B2t0K2u9vV1FFuuVfpSoa940gVU+XVuOx99qPvfyXV+u5EzNQAO+Oy0rkKSN+zZKthjtRP3c6FrsXKRYOeip7kgesA/2Um7qKAY7F14CeqVC+xGK9efElIFRGskp/XDDkbKTHda4GuFUPcYILyLOURRReXqjPe/B+jjaCFBm6E60R59A2x2rGPO6ruFLMNg59HM58AlfU+e7NAfCOENAEqmX03cdRRHO9eQ8vEm6XRhJZsPSyT52C8GevMihVbcPEOMFyoKo8v1Kvdt8voka1YEI4Azg21T1q8XKkIHVAgcD5BwM7eK7YOTaANBCOan0r62UVYO6mxzkZD6l1Qo0moYChu8u0oDoIMsxGscKDfMqMzIKkNqvKTQbpso538w92pWHOZbAQZ3pol0jBtTG7ygUh6mH3Se7dXZm3XnHSYR5INmsAy60RpUM2RqPRsShzPMTq2creHb8ZMN0gZDkeRVMH+QTqXCV/GwZiSe2oGF09uIBgcSuPA70pMA"
`endif