// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZJ0viKAhROBbLiRzAshGS0U7gn+iV2aZdr862kWDMwYtB99p3vIc1fTWzbMj
xFA1cAsXnhb95YF25+kx/VDeJmcdAgXda23wBOLfg+Ngpc4Ob6zy5VsBFHoP
HRocoZLoS2mkVFhR3Je/cHebDhXXx//li4In3tZvRSojXSfVTIpgK7uYStWZ
+EbHDmSsC/xGh0f1uaQ12OvC566CRWIMoDgcAMbmENZCOk1Me9aREH3wr2qz
oKBNjO+dtHBTDLCS4hmEeZcACCEiRGMgo2+kwaHs/7MV9YjWL0IJMrFetSuI
MPLvXOKsKT2jfMZYv0ijmM6sN7jPqXx8+zpRLo4uNg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aACbiAtzdfgwjjLmETG3XRg6I836JAYat+2eGLLcqhhF86LnfP8w5nT9yebZ
FDm/f1Mg5BZccdG1dqBD7JO+j7eiOR2uxXLw46Cqp6nY560j/UTlCY2o3A6/
ymNBoVowZj1X/HB0T+nZGh8T+rFPnrNYm2XYmOWR1YJz/UyFqKOkAQ83K1bK
Z5opy6YmVGwCFUBH0U8e0BUbryUyC7XptXJaa2bc30I/E7RuaXPPpdtLmt5c
Ao0CGUlPN3m/vuvxehcipshtpkjYYgjFqfFrjnbhWmqs74gdJvN1nIUU+Ju2
d3NF3xH+XvNcwFGKSAhbuFUXwkUdQtSzm/yccgm+0A==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jfA6jJ1y6KbPhWhKMulG0ofxLrOzSfFmgSsuohKJTdzAVHloyM1OX/NVNvaX
z3w23S0hEIYJohJ3FBwG93Ao67Br/Vl4CMZZlSDBlap4y/U3Qc613vyvTToV
L+RRjqavHPuSZFqCRmoXxuoYoUfQvh6U01TZXA0SR6Bqg6ZAsf5I5Oge702X
kaofBQIY0hoATZmqyrkuHev9vAOnTjLGIPNAEihtqufAwppLAqKUx3fBDPqO
AOjgoC0Pk4+4vjKO6AoOMc4MbzsarqWglYqO4D4zeZXpqWxbu+Zn80kr6ERU
hk2A8eg1uRYsGneohUEtN88l5m6JG1zGucF6g8LKnA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gVWPjh3XPEJBXDbRUdxvx+uoFEdlu9Cge+jh7bnm1R+Mj1wu7sr8Oxa+qg1f
YrS2UN5JH2Xj77C5JrflRqYaNLEAOlVjP1qQg6eARvLDMHPBYaS5MBSZ4qHc
9CbHNqNeaFp69/DqAyO5aUSTJOONcMK2Jc52jPE7OEs3k/kKy/Yg5nAPF6ko
rEwwXWP1xQt3insquG537ZeT4zK9dSADo0POCOeQS2+NepNCPbXb8LOK9Hvy
43hXvyTjSa19SM5WknNDQAs/pOEGiTFwnk0fa6une45gXmFT2V6aDgwhHpry
vux3UVaXIvQxFPoe3SS1nCFJRQreW+gvYvLJzkZqmA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JhuQcR1G9nELTfxf8Mg6zx7iakI8W6C1DgG3FsaAof71bXaa6tBAXl/50St2
vjuuVFBrgO5Qtj0jFVmIbiy92PJUtnFqIKiKGFCdBcD69sd5ykGOhkyA7FWP
vbHPjkOvhAdUhrtXOhJobMX9/rdJ6ptnPZmHNTAEj4Aa6cU8WjA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
QK161C/KcmHlJ2ByJ3BHJs9l/7APSoWLIK0Tm+ZWfPaPshdOFWUBDsI+FNBg
UD2gU/c5ArnNXSjyMhtSW1D+r+/aUz1PaWsny1n4r9TqvBpJfokqMSrN4qNi
zg2SA9N3sf8AD15U9iSG5TrptwV+rPDJcZfrfKWxSCFfvQA8p+W2XyaopUDY
iCdG/HW/gu0Y4kzMMWflRE7ixO1rVPhnjtlRVu643lwQx5kw0L2xwmxAGYQU
ImQSpn8bte4MaN+ICCMvDJ9nlEVm0teiNvDQ3x6BOjiS9WP9b/YvVXq08hOD
Ik5WZO5o8Ji5DD1GI+NBZp1W648SnJeFFrm3yzqTJsy6etf+oTAmuRjEGZf+
031lceTLnrBqCaT5ZA3J4CCBq9ib9Cuc4ovVfEsaIhdC8ahArH1fkHb8EcS2
6EaaXtY+iKPgbHb/rCztOs3RHqOSPvDVFcQgRkqQs93Mzj2UjpEU6hBw/rir
0rvaHQsmTG2i13VB7zgPBWISgGVscipK


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iSZF1ZYjqLrQPAfCAnQ8BEnfqqiiB158PgNMCvwHlv2uAhgUOxny1/rrrYXH
UVM9VzgftXAGcVZ5s1WZBQnpdTb4v17X0XPp+ItwW/TCn8LJEX4r6osUHtcq
arXKClVdftTr7FHoS6kDjampwKdYugD/KGp8lTmMxkf7YvtY3fw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
su+wTmECKCxJGL1jTbckJkwYGagYxE2/hSq610lXQFHUGVztxAiANp65RtfU
CchmudViEwIVNU3hFtLh09Jc/iPh7StduslmP1uVy+g4UU6uGNWuPjIg43ne
vpc4Ye4M42Z5wa9U8uxncGe3pPNT1HpIWjrqeHvpAvP6ajh7bkU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1152)
`pragma protect data_block
FCCWY/sgU3MEvReJ/A6BwmHvyVwwOQa6GmkWrOGPToaOmW7Q9v/wxnCkhLR6
oRo+K6n1i7dHu9rFzk2XXNfpLgeCJtKhM0tteZnBOZMH7llka/g02ExPVer7
eu1w8Sa4kczt2UwUlT1HdAQdiAUKR1WusTQ5oJvxH5/qyL/2W7yntvbmWa2b
9HPmgTcFrQGrZZnr97aGsYbY6aHs0kAwUzi2+II6qTIVeL8pfQ8XTLL9dJd7
xJ77euQu/6ebaESA6LrFyhpB0SKH3uiTUNlZQhXrV9vuuIta6i6Boq7rs7QA
n12nDHuPf/jP9KBmg95ExQ+sojKAKYE11boqL/JvhMb1mw+tnDNNYaYnGjKZ
wSHYq2v3ThkQE3ThOTPM9Te5FVbuVoA5C0AIhkqK8UCUcymizi0WYb27aBkZ
zAeascO9F3Y699bsoWyh5+BG2vbblA8ZRi/alK/An/3ZfBGGEkmWrbIUwcE4
87+AShEs1qCJcjg/x640NohTzylUX2PdcWGXzGDJ97nuJ0LcpzGq/nvncEmm
qQ6GImryR9EMxwaDWVWRKj1Zix+RUP9iqVoCBUGggNqiAIhP83Ek+qQzPSp3
y4Wug3OTUbc5gPHQ0xXEUvyIiON2RDsQOxqgaHsYLywLUAfTIC/hpb3iexba
qPyCt/XfNwdqzlkDCELwGdsJ5mxfhW96UbMK9IqHqJuL47+e+fhOApkzUjX1
ilSvXPyEus0NJV+8nU7zF1SzE/JNixFfKToM93i74SV3mhGVeEyjtpDR75WH
rHeTYoVmhfZq74ecUgX+DiF8DJigGb0P79FvI8m5YiUMdRR358soZVLrmMyr
ml9lI3/FcnccdRlCcRdEMKpXGsWb4PLFyX8jXUbATKkQuAqZ9MPtSTTOIwe0
BgLH2VumRzouFFHkS4pP9jeVtbCZIzAbMrdDUrwpSi+JFXYq6FBh8SAtcBy0
cWM0UVfgtC+czNzXANZeSYPZqIG4ASjn7PDqFQYJm2lRyaHlANsc0oFRPVtl
SasxvbOCnPldUpDlp9UtkHBQCkRLP2DNhwa3yxpC+7Hbd4CScWDkYWQQQEO9
CqzBp+F+db5/L/gvGsKzVd4fWSQidV0Yi5yHsNezoQZuxj2CUTOvcm/liZot
NcX1cIFABSUy9DWFyydGW3KDIAMWB2ymDirl01cgyeN++vX1lv3t5SR81Cse
aQc+O71DFH2Na+YuXEs7D5ont6Iw3Vju7UGdZiJ90ciw6R7n4CxsHvAI1+nd
UXXksgzpkgagLROEXgXT/Sx4r8KydI8ytmFagnWv56FdVSC0cSvYb9kulDet
uDPfOYN5V1OHgTa2oBpk2DljJHuIAaKpFnG8uyHIy1ZDiwOvAKKH2fq/yCIJ
8nrUrbBbsMhyG9HchBteXt/kCKR7I549RsFXNHM23acxHGYXYtjiZ9HxjDY5
ygX6q+p6HS2mmRT19xxCMUq+AFXunUnXuVcENRw17le0VpbRntRaRi8vikEO
A0bqkBFBjLpAmu2XFtyTpNw3EbcDMUxnUNou

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQoyoLEdPVMUQlxj8Yja2/nUqrpBH5zwxAMvTXke43erRdjqqhijsxxxV9u91eq7mA32MEREyBNJa8ZgkaOGcUzYNESlItPowwuq6Q8/kwCObQbiYOA7qIPnYuPJAdOOv15GwgBKHkxjd8VhAh/7y1MNntZXDXHBci6c1ekAPtzMkAB/7lz3E1CkVLdWucFHxX0yXwSzoU7LqfQ9K6tXQJOrVTFIdjHhiwDStiCW5gxORu8fbPCVAupoApAb38nxjnYczukyRJNcyqoL6Rl9DcFnbK/higrWXutm8xr74tlrr0Xsh9rtzrDN7NLTydR4WLgb4/rXSWa97wX9s6RPdOb459H3cSV9PHjFIo2ndiq+AHPUEmhUtuXkz1Bn0lavfPgWd2t5F04HqkzvRXQXbcAl/x0xnFITWBWHEE7qWEHWzCYzxpL66uWVpJAgl1zhULv4nmHO8WNe0GckoMWrQkXHexpcNUp9bcKIaUSR82WnvpI+tjADLF/mKwtiPeB2Gm2DIDyWop4HSbMInyB97jUuB0dTd0Lvj4N71U180CpayZrQk+DoWYoIpOHZZHwYdduV4wzI3g51SBMvFS6C8qNL3dScQou/GWKqNzIVluKA+rsHl6/Sgz99qXWtj6zOzJ2FOpxjqo/qlpq3RARsLDNw61JOtRs9U2Fc6x0QDRUyOexKt9II3KQ056cz/EbOaN2oUOvkOowsy4jWOPS4sz6HNh7PvlyXnXCddnpp6avf3b/elX18lKlSSxedoDCAWOfgqqC94Shs4nB17HOOQEtu3"
`endif