// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OsQBNqtdzGTgnIG0+NmLu6Ji4cC8YD5IHD6QPPC6V55Evx5BIUUd19d5OKTw
WVM9001czZEceCSIzYTAkW226Scn99RC5bfCg5GaMslwhsSXg8EZ5nJHomog
4RnNTn3s7Ai21g/3VqkkOVRb8nhFwIKeYaa8NRa/6z7xUitG5Bcf8S4ZuD57
7Erk4RUM+TXKExU9nQ2uKAUu/BNhuQcu3m58gpeobgMKTNneSVg0nQT7nZ3o
+7GFY3hymt9QTbUR4WBxuBiDslDpl6fYdZa9SsLseqYsJR+wIywHZ6HgS5XH
x8NECKxQtyrAr0MvtBic+DenpWuSCHWtbfe8O2DtSw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JpnpwqXOu7MVO09KTC20WawINeNON6RcwLR++hhehlHzkpdm9X7RWPqa95pG
UxKUsAE7x9uE0h6D/gLiwYrx3CQtjz/ICAuhexOfQL/+RG1gnN+dEX5Ka5z5
q0CLYbKSDsLG/9jRHJekduBRRmCd9AUPHjCA0yT4jLA+j/ugbgJtwdpnKq5Q
jvEMQoYT/0ZqzpC4YvtwybXWb6D3M//F8He99oPV8e3xWDoxRMuUorL8Lpoh
ZSN9HRB5T55iYgvZYnJnKpCRAyAQlssRXhQ+hWLkgGGK0nAPbDy19ES7w5FL
EYMcmaVJfTG/681cSvcjMLiR47ifigO0Z4XhA+gujg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XvjkIqOzvEtyGtMbMJsVj8o3xNINvY7dLfvpIRWcAEyY5vfiR0HmtKviJi1O
HR7v9WYp7noNVXx4XzFH22Ljrj7x++dm3LcgpzxbJQqZHlF0t8a8y6v2FsuP
llmTFEoZ5Lo+ztZhEIYl1lmxBAtYw+eJFP6hC8Ugtz3npkzKLNBJpEfYKccm
n1WmnmSdmBUKqIBd9Kv5MyqURugo4N+VMEkq8mZdB2234Mup3EzglvnmvWpf
s+84V4tENUAC+Zj9ihDIqT+zHdvD93H9RaKVImUvkJ89SUbolJRNK8eQ5KQr
hYyBeFq9YH2hHhj0RgbJFVx9Y3ZybuEwwQ28dvxnyQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fv+KxUGHEvqNooGO02tEl6fBXYCO+ygx73NQskcT66UL/eM2l7f3A/zf4y5o
FfDt1ZaOS7B0qNPAvkdQbq34xSdcO9qzM95NC3/dbfpcBtZknc6X/g3Cc/1P
L1cGiRkgeGTxKwvoDowGm+WEG75LQKUVPrUQjFAVGrvimF9vcnSFbCx5JJsR
qeTjkSK2mFxO0Ml2lqdNcDEuA860DRPeINvN5p2TnWbT6lBYqqUDl4lkcouM
u60mHE0bw5B2RMiSvnZxSmhEzQrfM4iRNzywNc9KWgR7Kac4XS2M1/411xZy
aL+53nfUWyOgks8VqE47PGxmIdDeztAQNDUjsH9WSA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hcA+AyK88ezw/s4xDDGZa9oUT+7vjsckp1mk3HJ7KyqusKxJANNA1MORZNH8
E0K8bm8NfPdHxS/jmpTCkzXga0/0645n9G6VFsDWWy01u4huHOfWaDXrMWIG
Dok4zk7KXPHWZNcZGTxv0XVDQv05OhXLiWmHOAIDpiNoRQGQCFU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
AvmWYObqnr4yjVIXVBuS1guX0yVea1wFN8Bo8OuVtkBOYPy9LxopFLRNYebi
h4L4L/uY9FgcKVSJJc9wAecTnjnK2wXvj5wnDDIQfrZPUy+D/BApvZj0pGW2
IOsHDCqnX7h2xdtmJtCGpBSl1sKvrqKRtIGz/ZG4bXdJ/0Z/u61d4A6Uoa5t
jgrCwDA58Xcj+JclMusYcNuRN0YyUeeesAUZ1XEDITsxNkViFywuWhjsmG1s
eF1cy7wQXMMO9eNVbUtQ/y3cmrTB6LD+F5iWh1NiQ0ctTv/5dRzZg4gd9fUp
OeTeXx+jl1027v6xQ0Q4iODaQBZkxUrTPWGwXHmEfnZmC6LKIYyswZzMbQQV
k/iVo/0QY1Iag58gJwBQofl0Fsum3nOU+T0s3nCyGNnSz4k/7VM9ErKUjypG
YenOJknRo9XXHlD880TufM5k8A5O9I25EPUweFHbZaDlq7K50uAaLJQMsp2f
ebtZAONyNYdOlKdAHcQpSjqoEwh93pvy


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JxBYW6fQjNJjsV6ROMXp3R/rwuOrmpD4OgDifKjPpvuN6BhX6B0K5Tw9BN3U
YTNtiZdwxHJax9HY6jvOmTuqefizsMvRA/jTHOqagMzh+wrptS69AZB/uxSB
o1P4ZmNw8YlKggvxQ1fNN5UgAd+jKSDaSOuuIadvlyNMel+XGAg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
F1is9vieX9c9nt/h1ZWlWgjckjMTeMVaC2MYwdQ53tZQOQBbZ05jDFUIkjzi
PH03WmZBz/GgrYeGmS5ZLYd96ZQsJpd/7Ljpq1UDro00LjTX19RjYZjvLwBB
JkFm04gEYvB06qjfsedhRQQodTirXUBfO45qR6O+oxjWlRhng7A=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 59792)
`pragma protect data_block
JfRQVNFcDJqgJr+cZ/t9s4cvJG4uLlKmzk3on/rUNZEd4aAS1gT1Id3/5Qy6
oPVDcQZClKg/XlCzaoxY8OI1FM+q1y0IYEoXE5FDdvYodLggcxd4yK+W4sv3
u+H17twJ6SGkK5KXWs9pA1cmaexmdN+024z9uWO8IilXHJnRmS5nKJ7Xkze7
O+9lCWs2skYKleib/47D6epulqwvNu2yDBIsxmYGVQDnu3kcwnlEis5y4sYU
GgKCqjlxlwFwb0H5rtPNS9DQ9jZVRGE1WI0xMKi+bjLjrygY5hk8QYALQXNj
etGtyPDJy3SKYcWYpYSWsvvhDCRa5AIS9MDZiVc3r6m6TNnY26RQeoNja/3V
Sy8EkaqN+VQKXbFwg/Dg130/zhyo8j1XgxwbFq9cH/3q77Xu4jfwDGxq6dQi
Jp593w3Yh8vMjV6O68ALN5GfQSoNPcI0TY+TwzsFoaFJ16HIux5M333UIPhj
fLdK2hxvzk+fcNMRkDAI5nKjpBu9yBDvp2Cn7R3bOJ3Z0qu4HDnUgPMTbLmO
w1AHmRJXaZmZd+t01ralGoQzslaVwrsB0EunPj4yDlqHXB//r0jR6T6dlUAF
ONHmHH0/NDvgDQrZHUAvLt9pp5QOx8zJcP1tRgO/AATi6VMSTvWkGXpOMD4S
T4xy7gdYgnQL2Z0pUynA7INtC8cteNYI3X2hYQpRlwSB5Zu39X5GnVM21RiP
OgdWll/Vw+8YRr1etOZZ6htPwGOI6tc0nee6LibvNdcq0+F5gD+Lgk7spzSh
yC+tcg7SHVr5vmtRyqq22S18uqx7TWc+Ip2HovzY6OtOMNnmzPdPzPRSip7C
jCPFMW+PiAXdD8ub8avJ+uoOWzdVxDsj05oe/69cNjMk/SRrPxI34PqkH7wT
h5iv+B8Wp9/Ytsw+Oa1oyirzaXOOhdfZzBR3o0t4zjwde297zk076fEBPv/m
RiSXA8gatH/VdajVpsJvv1JGP43FP/FtQmCPLrZeWvCq+HpVKCqWw8fb22Sx
DkKbL0kHLjxEr7sP3f1XfCQYOlF+Czq5LudFA+baBLU2ad1dMjTjNaf40802
m09r41yeGIdJTn4A5FNgzk3yY8ruTr20AGuUe2y7pEeZ0dXkzUHkhPCAL8aH
NegVaVMT0b+sc64bVj2C71wiYoNjTpYv9APGtei8nv3WBCSF8H2KnenAEEQc
kWU9qMbV46sos/+fRKGmRUXuCnX1C2rjcuNBwCuvfBMnndin71di3mLxKbjq
jQB/lBDcF+ZBa81W0S3zlt17lPsO5/OoIxu/nsuF9VouJfaaATYS93xX1Pzl
kZIvnFWN4DxddqL11tPnqdcICbndG6duQIp5ujDLAhKII8aXGF9yfbGHG+2s
Y7G4OGKQp1vLHOi4/9mz4Kk+nYnbDeLDduDRnQ1Zm4Jsaw1RXVymgQSSxz6D
IQ2hLKcvx+LFEhwR+GhDLwF2D7dzNg2DuJODrUgYZJQZJFqCK1wwYbkD1An3
7Qb4PdYf/MowZ1NISGIaj83QtHPfhN38KpgLSNR7mYD/TVZlZXpI1o7P8KGG
x6ibT9PsrkM2+YkDkGd5T6QfCu4tFAcxaNkj6QB9GIfI8JrTdSPgxwuZ0TJt
Kocla5dQYWYlLUq7Ycm+jFrCQCvFeM5+6u0efBMM+KyajL5JC27oyMF5luzj
l04VmIAbSSksgi/apOjJ9hZEALNF2iWVOJ4ivZSZMkGr51RhUBNewBrt4uNM
4mZCKmXCv7NlVZm+IGNZWM+e2d+xC/MJA44u4kwY99m6WmNQeqUk6dKo850L
nVfrabk/63xyBDHvek2f1cda8cMAzKo24rdr37jOxRibX8PJN+5TFEmbdB3R
S4QSAOsgQ6gBRzoYDaKboRjFSPf7EjJ+9XzqUOsH9Vwa8vC7SgIRYNXO1Kvt
ONnk2araXpAwonicNkOIh+Ge3XYhU7yEuCGu8kR1oxs8lONm6y9axqR8ySTx
Mrr7riXJSBtj627m1Kj/S3mR/gFZNNTS4iSPTIMiSZvYBPYey/ksSfzOLYuw
2zskT/+xKdUYZiSBs+0XeLkJBWhywnrvN5QcxJjj/FtuhLPPK+Z66HbK67xy
swhEQM5zKeQU1BkAUgWjiM0rTdqJVjFJ8ldvQTogIkXWfZXfRsPVYvI8pf3Q
Mhg98WLxqQ8nihB0pFEUbU+PCx6QvMzQ0gkC4bhMbzqefyFX/70oAn8M7Fw+
KTPgSukVqFkZevcATZG4vIxCJVACLRCprcjjv9rLiYH9iX+ZwjgOkFSdm+U5
aGsTsXH7ZLAZdHAVmdqcfUz8oXHqqAvIROgH73pSELiQ+c2ZsBG90YncTpGl
4/PeeWINy9ZlpeGvJweb7YQ/8ye/dk52IFpBndFheneiCI4d2gZaAcjPr5x7
ZwQFOPudu81LZKukUylAgQby/SOTAVfe6wPFSKYrMWXZ2JlERi1nRWsSo28l
PZuRFoboziSGPTgPGZ0CCth4WoX/g80nOfEwR0RyOa3BJJBdSMmKuby0c6OM
Z1YCmvWjaO5IifT9ngNoeCmC48gEG8O9EgN69m2FJi9/SdZWR0/+yL/j7S5m
GKrzi762qxdvfPP3WdcT2XyxwmzCMuVrc+KeWyyx/sUy2p1A181ELFi/VZgb
vS5DNk1JcJGN/uj2+mdJaZXkXIQwJuG6zHMSmU7kfKfCJUA22gzL0mTvUGcW
ZbYwISq+v8tsgjiDlhj4DrmoUAptqYD6CmV1yXf84zAQtJAADCfm6Xz4+KMQ
h7RpbTgY1uFql2c5JBe/qYlRT3/Q8HhJqEs7dGSIk2nCFNlmjw8zJoBS+EKE
1j20q46157ivVZzKKtHS3Vd+ibk6VhoPdc4PgG8dwEzYVaS007OIYRXS+Qbo
pZb2XXrJBBunVjqK20d+LLgoHexIvTqIle7z2I6kfGwMusNkJNUDHCq0REZp
G1KtfcusWmVWhpjPhVBu3r2ES9pSiR6y8bJp+5usuikaYugFCc74uWp4Z4B1
5ifKDcNc8li4o25lUlsVNLubwz+WLxHuxndV/ed7cDnezGgdJb6IJuYtMR+C
ukh5iIZbQe9YWZpjKNNd8bQEUkE0shV4VOKIqS3UUAt+euDMx3sEk0L6rxAD
PtuonD+xqI2P+Dg1qoaBIc6KxLypHx6MBwfa/C4OARDVlrBT2XqbCXsqEGuj
NnV2ZVwqmGJGmDNTCMB8c8dxWuTFyhkxbI1VGlJ4X50+MFXNKuXtpiRohxpx
j0z8cxZbA67jr9b0HcAHdUC6wS8P9wZeEU9g2VFy8tgT4rBIR8L34V1ST4tV
+DanU5i4paZSlUvJRiVuMw7sJDEIyQMiYZQs5rV/i5G1NoLV0hj1R7YRjTOD
DQlSNNoW8p0yyat58zRqhxJ5pmunWjZwbpFeJ2p22RG18WsRWgTdKIX0hkE4
tJrzEMNm3zgMVvb9/ntRbYoWpXXdNu22IcUrhPIcwlH629mQFdqTdsVbhi3h
RR/ZdfpBGYsCiFbVXPxbAtaY/2dOhZ+zCpZW9f9LP57kD/6W9kgOX7RTbtjr
Xyc/N/3zrjbfoRFWHg1nzEpXB2QnQNQpJgtoZQbx0qWRRz+XGptBO11Pi5EK
LXpYMxIxUqSnBUUehAE7kfbZAXRCLi4tOhbl0/uDC+guKYqtsB8NrbgCInJQ
iwTMTvqEgKEREIC90r9K/BSh6UI95pNPoQXrRZKEJQsxqbLxCLC1H3EoTO1P
931NZirtEFRsgaqTeJ4SfyqJ1QrZ6NSHLJU3Wq/LUwX4cbrR5IkQRo4uE8xK
ZNLwvXz+YCZoIw9FhpU7iNahVGVtW+jIfNDyeqb3X+XfclE1SOB4fu/WZqHg
u81g5r/daxK+mnB86BUQibLZbHz6sfnoiVCFIHwBpdoQQurr1AAI6cEARmOf
Hy/E7TgYQ9zvd4i17fzvDvjVUxQwWmhIbNk/nVipD9U9Zoe6qXOfKLB9HRFk
vqAkVWZlbXz856HgZ7tSx88c9dGWAKfnoAKlucjgL1V8biIPzpCg7MH7uIx9
KedJ/7fELXt5Gix5ClWsBqA4qPTdY4IbcMT2nCz8UrPPV3CAErZiywf3Vs7+
8aqXeEijL6vV02f3jKZ4g6XmxnJabcGAj/095p2HR70Pm/xVLxfpuZXtsx79
dc0WQjdcIEd0c0E6EuDegij5y/2BrWveUwtUP1SmVIGgR/NTnHrYy2rvmMzl
xMYD5xf1MtgLIfJjzFeQvI0z93sl1wZjkq6sBksHeHDhykv/UDGwdZMYwHBI
1IVTCFkVTYdgY/FDACYUqu1/Qf9lrBNjdMZ6m0zKncSu/o8tL5VnAK5MIyy3
0OZu90+67Cgj0zWqMYCxfNQr03f0CRnLO+HK6gz+lpEyYAGjRC4NxdJrWwgy
/keiqPbcTwlkhi10bOlOSyr2yTsdbzn/UEfDF7HcRDMPC6ZJEKH7BmszwgSA
1b0xc8vTC/PTBqtzazlU5gRlvCM9jbUTMccyFRkGFLToXkMjs8E/EVSlTgQj
QtIK5HZLxVOaB3CnJxntKlFyDkE5kWiBZjFC0C/noKlBjIcUPaqCSouuX7t3
UITwEuQFIzZRO5e6x+KKM8PstYez1ovZxy+zhAvKCo2xEKZr/i+9BM1XYEu9
YxvHPouO7/YIyMoRdDrpsmbwaHpt6sHSzXYZFfy/NudCBMqN4j/ok0rUUjei
phkJUhvIqXOLWrMI/YZNtth55wW7IN3b81i1bdV7VMvJDFPqsR0MhC8kRdC5
fDdLzsDWOXbeZJNUbFUZq882u0S+jRttZt0eZ5RX2eCNeh/RkhTr2ck2kLRM
FQ5DZ3i2gNE46umOYaQ1NdyZRxve8KO54uQDL4Q0y4B0iG2Uo11xCwsvGJGR
9X9OAaZhfom/w0FU8SUKp1BGpMEcpTKJbmRdOV5lUIgKyLbMvjNA9MoUrOb3
BsAZIz5krmHmOucLwGMqtubrhRKvXm4ZRERdKD9hUH9aK1yG7c8sODHkp8jO
OgSQGNJUjb/UmBHxb+wfeqlIi28AbSnSUUdg78C5py2HN3SMQMpi5LA+P9/n
Xq6LDqLmdWq+nwfWST3FZg3KOM85oM4ihWazU4OS4bOG1AL+qSNJdNf/ed6f
kDi06+UAHXMuz8d/XSnHFNdNe08GBDRHZ1rQvPIWS2u6Knbvman20uzDpXCk
SPrDmXIFX/qAJKU8bVX2uv6ORKZF28dCEa215na9gCMOGC58Rm61pqq7iDQk
bKTv7uMbuqXtLKqvk35hQuawQA+zAE7zc+j/2rJGR6lhT30HuSeTTEDHAqyP
j1tIE/c7cWi0RnHdbuUDauJSyhWK6qWUCuovsOMepGbqF8xIhAgKuC04ajL3
XkjPRQs6Qd0ZoNE/5kUVMbrh9Mdg2Ys5/0k0oOSu0XGL+c13X+M5aCPqd5Pu
TlNmHEmlfIXPY+xWF6cuOajXP2lK6VYktTndkVkMhN7ZKOqr8nzt1VjIf5Mi
CFeFO5STMEzuzjKk2R4RRYPSbMEn1dy9NicPhVxNepSCkSD/AotUCkKJr7Ob
HxggfSD6PVvOWWWRXb81jEBT7JiAOqs0tdwj5g+QXD5PoSKFiji459FlKjle
RDO1h/tQZMXbpOkOtWhklPps2noZ3T8Bm+xdQhH+Xai4awitjt60uGS2RgKT
BCoICSBrWJ1sopDDgo7n4K3cdcmmakplzxMZ4HKPT/udYVBNAqpKdZE/lEaJ
pbKpzGke+bOkts6s1Y/zIkKy8G8rnkWTiGAxR25ccj2qUvHLLhGO23YtRhte
1NCD/Zywpf+uOSCaC7gE3wqhPnmD0X4VwqEcDu/ooxwhhjDdpSC/UZ8IdKZ1
cOSOAWpEeZAa8wRhnPaVZDn+3xcIWGUwJPl0anhNyExnUyIIZDkQzB2ZOEHO
lQLExRvkLhkPQWFqDXmwvemEed1ja5XOVhm4ZZNVpl2EBl0hQLFDymLIPo3r
7FeAmF4tWqcQqEwSUHIQj94aF2Knpn4eRg8szwsPIoWwL5LsSN8B8M2VHB4K
tV5ut1BnJGA0Fq7qzyLDLempew2FlUoE3cVxMXqqTmJzi/tWmjHXXDAf1XYA
RSXQ0U1hpbrUbWe0C9f4+pkCE13OQdVuRVCzTTxX5xIT3/u7JmrKPm/9Pokd
GDzdE2IQ/FykFs8n/LnOHsVrYwMTKxJmDB2lEVa5uvlm639yOyVrkJH19ypE
9cORXsBhutBBsYXoiIVfmCr3E1QjfzdWnc7CNqdp5+hm8I8dGizrUkPdeQKG
eH4JKN/mDTQReaKUJj/tDzBBhLPVIqDO+6NOqlKKLHP8x3WM1KANHgHPH7up
pMDMSbA7et86HmwK/0rYpOPgVGx0a5pof5teWfzaVm98rBJEpB6Hom3zXM0W
7Qen7b1x4Fy8OwUlWbTKfTevOij4qZ8sH3XuEh1FMIEblUASt7i643zRKbm8
YfGXZ1FKMk1Okql3kU/6P5O5brW9ibzblcQIjBOyBD4Yohf8j7HN75MMZMJi
OSxspiLoIoOwSIcGuINmgc1CXd8g4/UDttWbEmr8f7cz7K/vvEJ+Wmh7UpdW
L5Rxms0JlnEV2KalMkCejEZRSuiaQW6dpCs8KtxhIDPIO1MDc1WLNfhlZpYV
whdOuULZRknvltmlperOBf1drZcutJQI01Vxqb2Q5Nk/vjXhi6LwmB3zzJKp
KrHJMgDCCEoZe3V7oVba0N4LdQQ6//Tvw7jqb/7MXSEaESux3tjEqB0ixjst
jJOiXNU4aj/x0onZ2iZ/eSjI2tiBq6pCsZ1Rus7gYGl2XGRHeJp5gQJCfk0v
k+1n9xt6YdAKC8mQCbsdBuPZB8uLpxez/dyzbV20hX/xwG9k7M2OeB6tchgx
3PpI+Z0YnAit4TheAJwAtmDaaoM1G142ntdaDinHJjsG1w3LR8vpi0M9muxa
nDgueygVHnuT8J9pWrP/1pKh0TygFKJ+4pOFzOsrk0KSNPPxRnuI458MV8gt
IjNSYzgf8QC5MgtXPmlyNL98rx/DZlYt8WPH4AoynrJCzTPEmZ4/kxEYzv+3
jioSfczM4ns7693OYXrzNwZTgUWAxsDfrveUYgmDP025JkEinKq1aNdvemEB
iZMHMnNKDINP5bB1jPboCkE3TSJPpywfUdInIahwlEgE6s96yCl+uclX+4nk
K/EvxNCYviaotm+OMDjg0WP80XygWncUtmoB4EJwhGm2WGlQOwzFJA6iVas3
P9jTlm+zPPiCgoZiztBGepHFBR13hA0Yyh34z55I1h1KLYIvkzsy8Usty6SD
Z2heRQ94nzvxZDOOTbpiiNa3Pnybhhx+fHfq1/DLFGnw0wCctAFKW7xTr+dF
6ITsqpzfdVuZkS/f2nMIJXvutRyb9fenoraVuSZrbwP2NhydHBI08wOWGvQI
G7wgsHC8ja3FnQqtiH7fjOTC2OcE0IqZq1GpUZDIyZmV7+dur7XPoF3zUnH4
tdezFP3bco8xpbhHioeHsK06xQ4TyMwtxsbgl7jaZWum20PnB2UptKmfXdzL
p5OltBdXcW6lVZNH8bLnH20lyfwKrrL2NJGMMMNI2n4gxbqK8tIynrPwAR1Y
/EvN3T1UsbFc6ZOLGKT4NY1TjrlOQfm+sW3Wq/GEMDS+wq6A0Ld8+uQHTe9v
CoG3EkyWLwSRbFzFZJlbSnO9Ve3oqGA2qoyhBeYjLVrUNelYz7Pxn15V8xqe
R0/YYkfUy/La7XNuJ/wYtibvkHLWEJGaw/stbz7189sHrIJIAGw9sR3wjq4N
OkSoJz6dnR1XfbuTheExXYJsjZide4sb1x+1etRp+x9uCHVGHKCaJZJ1uMeD
6bN56U+qJUpWeLE05zoxYjQMeuWZiMEeebxEbEWdfDTFxBV7MQnnOhumxdzA
bsA7+f9IRdY37NlW13PVOTaWW6BI+knO/K3lG4uR66fudkW/TgOcXgZyQVTL
aBnmMtO1NB0oWML65FVQcbzf3lgfqJQsEHS8YNEl/wyZzspP+lNLgkY8DDGW
tmofaHpv2GofRsJeJUlY1ooXP76wIgkOt9bNlqq5G8rCJ7dci1RIMop//iI/
B9tdp1cjOKyV65qIk1ct1zN5X4FkVigxacItXRkFsDZO7+8CnixMee1UPhWZ
MI5VktzomAwtgzqq21x10jPIF3WLH2IxapUDwKokilr8RX0eWqXMSeQmCWnp
ts4erHGRdoN1hi9l/TJ4sMpnM1EMZSIIlZaG7lodNILsN7ZSEkjJNqTE6b59
0HrCYWSX3NewPt/YF99zL8l/5nHXO73XuO/VFWnbaeB1viGNCDt5gW1P6MSm
w0eDtP3NlRATublntFrpgXxLxfH2nd+xQHllex2YRJMw7VAyUUpwh+8JfRL6
kfknO0tcJZqrC81VqvAwwuY1akFCYB765I/+WrnJOjd/RuewEV/Y9vfjbClh
C7NQjM2M7dWyHRUf9wWye33lBjqc7hB0OUvZ2wXw4QLvOf2ntZ8WVC8qs/vc
nbk0NIHUhmcfdWderQSyt2XcQG+9nGq1r7mC/RO6iiIsp64HD9/Ec99Z+YgZ
P0bGZ5rBaPHRGEo7ftB5vmMPFWkTGod3Q2l+xZ3QTJ/ZU3f+6b8BQXoFBUoc
0sduwt9tc2oH3YqEPSbFKaZPjWqcyBskRj+FHt6B6VlQ/TLenahhke3Fmuzs
HA6I2KKeN42zDFuT3FMUlI7aeEWMENUDGxaRqP9caMucRywqDR466dkR26bw
lIZGsAklHAC1/rYsE82ZQh8pbGDuQvvGkqA+WyYDp7DfkzjsNwE2TD1e10q4
TfqqUNCYR64kuJP3TkdXADlsDy6ckIBnGkGZr2TW3gA8W7WrfKxZb8OfsRaN
PgH6ogLJsO3slMt0qqd3r3dYcAZHZRoViZM1aqituhAS7SzUrmYi7AQMWXWm
dB1A83fsDiJtNm0JkX7Ghl0FlN/ORmmfirhGg3FRx3TQa978MaLi1a4Jemg/
xmaZ/j6JQKFNsXLjKyD3v48qdudEcuTUT8M4za4Jbdz98HC7R170ydxDVaoH
4q8UzFjxdtVHUm0E0XJCo9VGBtQhQyadYNAL9bdzXFJNsixna7c4PlV+dXOf
pPOJqwgrVxNzl5sQxcVcH3a6UwnTC+70q3VTmTFoFEyau4EZobgVfh+Exw1t
IGzHeQfZRI8cguQXI8G0y67lQMCnnd/aut5NoDpWouAfg1woqTzjjVK+DC3G
R/47InUfkcyCY4zTNovds7PaURNBRY1nc+fLV6L6oAUmcUQQE7Q5HaQiY4CZ
sR4hpieLcp9VSL8o1XeSJ5ABjUzt+YvSK7CszgjrOtcM8VZp/trM3aTbAJ1K
Np3sqeoq6bsi9p+2z4EQixCp9eVDyipEV6GRefZyTmexfGwuMIsKBub9rjgJ
3/v+wtuycuVyKlP/9bChEPoRc3XCgxjLhci2V35wsK97XKssON8zg6Q14uJW
zNmc3gKcnvFyfC00LGZWQKG75h1Iv5Gpg/Qq+9pqbPVDofw//Ex6LtuYVlPo
1650fqp/GONtq/XOz0jR7lZ7IQ27nvgW029ARcDQ5W3IasNjUBCVDpWuNKhU
5Jg579h6FNN41o/p/R5ykfR7LMfv7oZYeZ2NqnMqgeNWpA4I/h+ygUn/BRZk
QyxKZxS4s0fQwwDa3KU1sOEXm5YqzpgdExRZnnkj5XTByvPAzsiIX9tCQREI
tJHwkZfGh76u2dc1uYrB31bD0+Irlqfyf3tDexQLB3UP4t7vDdoM/VEvM7VR
lwUrRwojd2F37gMn7HLjbXxUtG+vgz7MKDP3+hhgAuLBEfOFHzvFFAIs95qd
GHBNVcDn3JxrEZ00GheXbvC+Ky7A9/z2AwQcZpdZVKSn08KGeJvs3Xd2uYdq
SeHHA49PKKUSoEVr109E0wVTg6q53VK0zNUoGMqurmZ+Nh5jMBZapLM38eZ8
5O6yWczbqZg7pgUUycPWkY9t1czMgYhzWSLUneTvjlNeqGcIPRk2e9uxEBga
0WBDkVATQk3ahTE3+BhLXveFqBxxJ7UPG3d96x9PpP5xebU95bSpB0mgu9a+
QfRb43y4p/4/uWB/HxrwawgXtZsVNEq3Zr8l1goRjZeZIgiCnso5f/+7Yzh9
Rc4tJLMgdIntl6tB5EFyCXabxOkRSNTwt+IXWbA1g+NYHb42DhTluezGbGqY
vaO2aUVYCDnVeltM2zf6CX4/QzH+uz7a6GIe1pNRl9yhebddSUvR50sZmYr8
Bg+FM3QrcVDnfUBZNLNFKFdVO1pvECMz4d4+Hw6YCC/oVt4lA7/3fptZpKY5
kaBM5eOuiAcqTzM7bsbt9jf2jL+7SQVG22cGyko4CRxSjplpKj4eoJrdIvUA
N+1+n9N2ROpJjF8BpDV73UqBKl+OKICWCAvjHFBFuJYPES+5tJMtLHz1IOwN
PA+posII7nffWyphRLHrpan/ZbSxPymDJ9K5sKGdfuv1HW06GN6rVPrw/b/L
E9kWCKGUQSav05aK8tskt2xxTAGs/uHKeGGdL2VA55YRuAH3vRgPwG12rDCo
c5fLOZkKvHYsvvc2jn4TQaleKkG4JdQ7nVQG/UdXCObJHElp5BfmEanWeWkL
ac8zDXRrYitCnYH84ncBsnoAur6f8MEpwg9lhb7uGE/Q7eXODkOObdJx4zhk
/nxUbs+HSt4eiwcDIF1odYJx5I00Ma3+LlJVSuL56C0R0z3RebJyv1WLgKcA
A+RA9Ys+u4GdlxRqX8Qdv+YJsN373EW9BGhL5tMx7SILjJQLUdAFKxyMWDGr
JAVNdZ2NKHs2jg8o9fJHI+nCNgjF/ZuNOK8CQrq0lwSagH6RBqCogyvoELM8
T2C4aHFJ+W0buiydDyeZG7QQygle9zBqN8YElu4Cm1/331hdIdfct1qb5TiD
noQCxBIvvpjSEQ41Gj6Epu7EGIn1cePyGjtesGxbeSqP7gvUV99DHeMIl71c
yghVIUIc1N7arA33QJxnM0e4MAxNsC9KwAq3bz/A4RWvVqjbHuJ0w6+9SAul
0Sp1jn5DjIvID9vKzM7OY/CNu6NpDeOzTAVlLe+PB254Ca3JH7eqefgJizX+
khY+LoCgjXzOEMBnubGYWZAan4Ac32JcwwFAYA6Z64Uo3p1+GVDbcP8XIVmC
zWtkIJxeFEuqWoIKDgpTyRoLHl2U2NhOlHdzbf9D1wHVHXraVLZySnZbaB5n
2hBm2Fi9wL5Pi/QaEeSZNjNCak6jvRD2d2CwIaiAG7JiJ5g8SxyYw9O5TdJk
7XNrIRYgXhrLyrCnTkqdscQvLgscFbHSwWU81tX9glpGTfPYkqd+8jQyfWst
D2Ni3W/30DWujTbyQM4wAsTYI6koZ0+jz9tjTt2xROqq5o27SfW2jezEWS34
UfMN18A9P04Z+AdvgOvA9GB9cQjgG5cgOJK9fyviReaJHbBrzbIJ44T7TYc5
uDZSYGxY65H7/26XZl6f+XLwWLSZyQ2RnRyE2GAlr6IwhAA8e7NiGJzaHroU
uf3WjYn8eeReUujPgu+cTs8E+gdbXlTdiG3569RsDZ8LbwlEOHGOU7C2e+0I
Q0I5WcKBZL7WSVbuXHCT0t0g9hzhEvq8CWdC+V9bPy6R9uPhz9Q5dY9/aZYD
vqyxrf2nSlGdkOXxjY13K/1wmV7ROZpLI+jUAGh1sh0Gx2W0hKYVoMtRFSdb
mVL2zCRVdmHtUUH4VRplFy8Z9dxv/eK0NYObmE3lYJg4/mdtN+BhilhOAt9q
Fo7T0U4ovJ4ptVvLU2nGMN5TKdN97kzehnaPo19lrYZI/VgyK1+CeMykOWPn
hCxsNZvhAyZvznOYPXn85SlUr0mq0hylf0rpONvivzdtUQENpRtx0yEVnf1H
Ha3RJ0oKVyzCfg0QvWAlp1Crfj/c04ZNtztdk7dehtrRhUhGzDtz36HMkzIG
+KZKzD3gxHg8rGop0nt/T3Yj43cqtd4Yw8i0Mw19lQnLErqGbj6yPnzTmFDn
e15laWgBtojemxr0fRXKajSoaRnzovdKqHgOP4m4SBdx3qp3Sa5erqYvWeXW
+yAAOiCX9i/wlMiUw3dBy9f+CrWIlTaxERHN0HPTUEyp1mIJRUFjfVz92O3D
fTykKgHV3kheIbK6VvCEAoC+q/lew0OQJf2aGja/AfhPvplBTH3zxNg151na
MHxoTlmBdrZeb226thKTROc8ltCqdWmPdIKfSRbajE15PWS9ElaVDDGbSIIf
X1irEnaL0IHObSMvwVf8nDDKZH6y9LJbz8t1CANqe5WgjjW77eVU3mPPbHMf
5nrI7m6IiK4a002ElgDEd5jyFB+QFnusAa3BPYerNeH1GY7pZn9RVAfSunau
VCDcGkuoa37liP0E5TMuVtiBzs4AQXPubkGNagUYx9Dz+er5n3sMSN6KP81e
3MlmAJMnn0DYpHiUp7Td8t7n43G9UAMp8nLrDZt5MAfeYIGxw7gyZSQx4SO5
M/Fgl80Eb6mja3hZtynNhc7O5WFNXYMWdrqQOj5O1yNLXwTydDGPgmkCUPpG
yBE1FQme5hHmR3EPNeV8LUOeFvQW5GEeWf/mLxyQxn6Q4FIpRGzjL58sOE1C
dAb+4UrA+xaV/exJ5HmO091sFFJd4INoTUKlYCAOZd2Pojbobeukkq6vjo56
uJw2Pv/sa8sDWlXtAR7DBMLsZI7x3M/YfFI9BGWLf4VIOlMtQQJC68xMRYZH
VNkLXtzwS0hiBeg5g1tnmCTt8ZANDTcgBzIBuYhz3f20PTw7xElQaauo8QAM
nRZOIHofVDZz4dpWZ/OzRJ9rEYj7IGa/zlQr7QJhtfavP/TCiR7v2iZeUM1H
fl+30XlUrT4vzQgTipMRLxiNuMYPxOmsQrEvtIl7U0CqYautR3TTw8DuYNE1
iCHLeHYV8DH56st4cBIWpQJzZVD/s7Ys92pHtvYdLl/XGEyfj0FMuc8h5A2r
ttQ3fkn5ctjjKC7/6+xIT6Hu9pZl8f3BY4j6V6X+gvsuzfqCb0ahL+p+kpXF
N6ptgohzQL29XppEZlQk9N8J9/z3L0IFM7iTQFNSmqTgW/2u8hqLE8y0OKFR
Fs/DyT7HFQg8sKdOqF77Z3SK6lSlBFwFmvp2ed/o7yDoyhmXUaPo+ojIM0hu
5GjJVoPozl53hzD47mquiBQDd2mL5cq6ej31bLV9c0p1k3XmmfzmYegGChMf
NBVAd/HvrN2xoOg4BJtYkPnPH5ffr9rKKVW9GWrxlk2+QHT3Bd+8RlbQKKo1
ur9q1Jc6o/fnpsKH0aqtHTQNG1bi+OoNrut6eoC8UYpnjqD8EIDaJ9xfJ21M
Vj7bAK3s+R1lRRGLui8WL1Dj7I6l51Y3KKYauav01Wpq/haEhL1IacmLUops
wdjPmj0pgt/GgOsX/zIlhenVjEZzW0238VMTxEdmI/3OJFjkY0iN3LvLAlN8
jAziypLYTNzyNvkq3Yr5X5JhSqM1Iam8Fv0p79RKO4I6lUO8xHVcKRnkgF6p
0vTi8BUaYXIBVhOL6TP58io/L6Cim/LvDVnOEyg6YgvI0E2R6zCAyrJa675s
6EFb2Y+PnVl2tYDRaNUOQLv+LHd+DaVF/CYA7UBiEHUxgLfHLmud+mM7+P1u
kd1NF/d9kq7exFkGIYQqq5omWjhpsjUuMdj8YgER0WIeKqy9rgq0L3bCfgfL
/kItfwmvaMOkgcX1edMkOEy0R1hI239Svr5pSX2D2PB0uQgCEW1E64ktry65
WK63/t9vhm+E2Zy2/0v9l1kjli2XezWu0eImGiT9cQuAcQeGffGuhgLxQtAP
SED61FwlwmLMETTKQAY2djZCtLkD5iurTAgVCRBNr08r0Ymkf3GssmCW6VhT
JvYpnw/2A/tYukIU6eWUimMudVJBtEBCtqV+5AF2M8axc47/YxxS4y4ss8hw
jjDmkHJp36UyWUf1f3wDXWsvzpliDBWQAdjKOTgOBskQ+xvfFpeekcm0I4ND
rDW7/WeJOSw/CjhuqDNbYHuEaLMzW9NkhdG8y1AJDLkb+tjVsWy9+KJAU50Z
3Q/T2cGPfWuxsojo79g4hOhbJAeMXxl4JlgDEe/Ivg/PGqBSuSmORfA2fxt2
O0UVC0mJS+GdrD1SqbcBPEtW8futiKLn2a+SftG+3vRxk2kWzfxM8Ge7UpQr
RAH4v0eW5AeKS8j5lWlEvVNPCRdKXuK4y1t3dQeUhQ4XZiNSqLbvKiOw1fNc
fXq8SbDOcG5NHV+u0cWID9rZihhpwJdLfupODPoa6LwNZZ35Vfyu8Smyb3zX
Z22uvXgB1cahB1bq/RK3FmJc/F4FBKxhn6FOAs80aAk3T0VGpGTold2Mydqy
o/bupZPsIqO+sCoYcvXprGW2nZOseyeRH0ALvxNHBjwAeigscagI4p7+H5vz
3OU2ZUKpdw+AtTDbrmGef/mzvdvOS8SzDoOsbnRajt/d7t8r1TzQw/HuS1uw
uNxjNdUGeIC3aXEQU6awnWswxx2abE3ZGi8+qG9QvcpKtKKv/yVs1L+KjlX6
oOdjn30Ymsf+P3oV0ZnXBgK7Mxm3fbA3MKYKpQqVGPySU6srdGW7A8ViSJbt
1fOB8aP/cTKitiOAp4Yma5w8fiacPKibtkvv6ASUrVcUaCXHqsgOviLYJdT9
ScXZKablV+SIgu8zh4rw1+oeZodDFw0I+2jj/L+uumDnNTEBc6Prl0YH2HFB
BxUTI+jUugOEgKdugIXXox8OpP6E772VaSBCfCinXPWeyZEwkg1BzCzQGIpA
8FFMjLKWFG/QMnK0voUMGMNPzwTub8SMdUjfEDDhPVefqtyFjgv0v8n0DTdS
s9U0DaVYvcKyHe/ATcrwLC2VS9y9nlB81YQjzTZTBEapZ0WYXcEhV4SsrnDp
6t2p3Oi7rQl5D7THrWCZPDR2IlqCDElTHdkIdY7bpUT+eXiojl8w17eKRoli
Ci8K83E5k3nGm7ifckK7ICGuYGeQiP3hNSF0SWXVkA2Wn/Svq/vyeqQ5ocow
lguF04todY16vBKMNfIWsm4GHPWokzy9hxZE1RvV7dzUneQ+a7N2lTFP78JW
iCPzcgiHMFo/FDa/Rmj0l4HppK7IO+4uXkXoa3dd1Zn1Ud5erFBwi63J/VK6
p/0k9lh9zR/bHhEpbhx/jtk7L6Ezr+IDHYVjSV8r+2Ccjk92zPgCzaLBRQgU
ckJ3eLFc9+3MWmv4BpEvmDF0+eCpMOuK9kZX3Z1h7wGiqQwO7upEgYL4rE9h
qH33EO3PYvryEEw3DHCXCKzepzOCctzBuVvMrZ2nOERsDb7uZaoC/8OEV7Fj
8sLDBAZfmnMpfHzDwGxZk3u39x9IMMy+cnf8GgDdxUmgrdJ0Sx0Bz/sBwxFo
j/e2/P8IPuTv9TG2QJFzmFgb7GS0RU0G8Ily8Kjq5iU16rgpegbvkQGwzMDD
HRaafA3wFp4ctXJ24W4jpk+ITcyc0JzpxTLLwDaWyDcwKZiLRcytHWf/zvn2
aYfrf0Fmi6ZaoUMxcPwG4DzEsjIUZG+gV0v8GhZE6Cre2jE0ehZpOinLv2OU
8o3pSIgYUmhNkOKlM9TtOwHHok6GqceIer9FpZIfsLtBdcePc6Dv5QkTLHby
5MKWF4A9Q8zhYBM2eQdYsGtrV9ipKGcPVNj8ziQrPHbw2N+gWQnS65HCZQbG
LoG5JlWvovCMaoBVSoElOaCTw79XpuNBi2FmufNKBDnv+86tmcTU1ifu8Tvk
BiOIhV0lQiI004/RyH0EUf6sObZzos72He4TjSXN9PAwOgUAdi3WNe3R7eQc
xPBKHAwsXGrSSM5TrQd52kIUx0ja/5EzMe+ZMW1pTyBYV84zouBnLS6TEsIy
EQ1RNWq9RcrNKUhaheQO12eMsCzoifZp8OICjcIhA0ly0wIT/bykj3mfYpQR
MJLyq2pvWT2KqwY99XEbM1QfuP/w0zok5GZvsM6VFeATKbZyi9dnvtTUAl5D
dxY9Lr4XAHgAZYMo2ofb73Pck2NKXzIc/OwyxcwE22SJGBhv56Pf5TVAaK1H
Iv82bEGSfSzHNtMblxzjmyOW1WnCf2BU6secGF8Xg6dU8qpMc21MmiX1XY7f
0RHYWCU+0tgLExUrm6aRtvg36zYMLrvU8Rc4Ms0VItuhqbc74ljhU56Le4XU
5dCkIRuLSmp+E3hwWSTU1vl2gZY8YEcemJxqFLNJ2vRVLDE1t/7xpO9SQ6ct
dk7BYVMwAuQgue9IX0qCmBoAA4viouZbPbySjLxbaH/7BIv/31tE0vktC0li
PGJSOQSYJjpIbPwt8+7XtejscHEQj1yJ/S5iXPDcCw2eG8Ro+OLfPWvfjyyV
dJ1a0LxMhIVXVLoAAGj1UeNz3oMyVboIG++G2+YiU7Wo+q0tdasXdm02SoRG
WaiJrVmnPJsidHovjQmf1lyZZsTNpDnAAdo6spjQL1nVRx8oJRodZs90Co9E
iYgDWGxXyl6w+bUvvhaWCjpr5vlWX2rjPnoOBpvAQwdTC+Pv1pZnW04Qz56N
NZjKRpPhVLCsmWXdW1pKM7IcnUp0bw8r3DLH4lj+EBy1HsLjTMip51EQzDGx
3AM3aKVEFpkcdx1OgU9q7+VVdvE/f6SAzoVPNcExbA5ueenYo/CYGIs0/55V
z7NhcjM1PVX5fsLkYAQ7GOHyYWwAnPJ+iKyCCWmkUqp6ZK+pNjge6SqYoPSf
X+v0qBTcqwHb5yVv5vexZA1Mp2s0UpgTi/b58rujsmgVcuWQen6312VciXad
6gf6NYXbn51vUhg2sP7jV+eyCBNsTqFcVeQtQQsai4sQaAy5IlNI9mkGZNwI
F4YPsf0vYhKyZ9ZxuHfTqwQeKiuu5hGu7lkeCl7H5rhQTUnhRPC4T7LVHKAG
xGtE+FhShGi57cSZeGPYI7tfRjO0m3S9TUOmMbE81OJz3vo9ucUdX4U5WWp7
m2Tx+FTMxWuaw1C8m2HQrwU8Kk5uZCzySFxXhjeZapcil94l9+Ea0TFUZB+b
uKv5Zk7LneQ7gJMpEoDwI23cnXpBzAmo+9J8yf4fNbJPhuxgk4VRDW9rUTjZ
/kmG4cPEymiyfU6Wc7sN4seND1y/I8ehHJ+RuPBIxbZg8zj25tDy/s/VnQsC
PcDvtCk82gbfTtrAOKx7IxL5n99Nh2TM7tQ0ZyJ/gumvNRJ1/dniIf9GRRdu
0n8pWW1La9tvFIJq4OpwmVbEWw6Qla4iG5WlM5BhoG1ypCcOS1UbS2DZD4m5
gIucMb/mfbeXTOPQ23+4CdxEE69/K/cZsHhwCSnJBKhSKrgQ82a6SWyHHVq0
LCdichulju8nc7wLFfi5rnaUXt1NDPwXw6/iSL6KMa0EdKUDoG/7bI57im29
Cb361C1Yn1Bn34gLbrjCyJu89VPRNS/dZ4TvEtHJeXrlq8akwSKJSr2ZYRZ2
zFd+JLVKp3nMFDVyF3hMXhVl1sC1SZ/T12+tUqCl8yB2iXCuGQxK8VCU6yd1
B40E7nmtpNFHQWyUmNshDE/vbrJDPdnm/xzMhDlfPIHS+f6ESjrUnTmTOLQH
yZXg8xNVt5REl9qvJslJ521rF0uTiSE6EUZITa5LW9uV/+aUz+ajc4aqQzAl
Dlqyhy7kBnctavmKgvRv3jn+1mFtcGyMJ7z2vsOJcJhWKFsi7mSQJxkhuDqn
WOhQ1agVZXX0xXQOr1QihtB/3ISznWw/W494xNYxdjiX4+4DiLtypy8WTgRE
RKQJGxK0cVLdFotsYF0HPq0v3mbcIhfARIZcFx4tkV3l9Ed9BFQtwcUZ5MSm
vSArShOOsSnal7kMKpDlw6c5ECTVzXKb5gXEE7Khq6y/GX5tIFK8WMUL5dn4
4fbkFYXTUSQ8ngtcS5HPtb85eAGJRpw0Cl3wu2n774LTBBIr0xrv1Futpp+p
QW0yfduHup2ndBprqz3dXAppUbrm1FUliiH3TbHRIUr0Xq4kPrWNHk0BqvCD
6FS4A5RgGz6m6jMcwq+tUQ05jthsaSk7eSvze8ueiiq8i2g+mokTC9Ji+Ake
RE2OVNptzq65XKyTgtSiT/TuM+7C0Rp7GO03Leml9GI8y3m1906XUuV+V/hu
mnsu+Q6Vl3mAvkNjQWW3ZCoMNBx5TfvEXlBV587dXrEzuATl6p8BmKfDFv2y
4ekhZL23qtRHeMq67eXTQJop85n+G4R62kje4LjvbUqvmw0sRBdwg3+G+MmD
ryqgeMdA36wnlqo/I+gWyjLFywip04IHbYnjE58iLDGQupumt2bwOKXMdzh+
3Ulo46MtEWtgsuBykH5T48iRm0BGU2HyGNcrQWLd2/JMqyy4c+xOn2v/Qqr9
paDRTNEmYIyaGSaRJ9OnEuH4ETT9cixi+JnJzos2pzb3ap4ND6dKvpfStzDk
qLBY1wyX9HawhkMMEX4gN4M5SI7xqqVmUeG2fBBXkvpMGdnRZx7sNfh7O1HP
j2hqaNL9FnG/xoVA6XMeX6ao9Yci0IHXWLW0k1dkgl3peET9C+r3rw3xb8n3
kn/joEIIPxiBxOzFjKE8fTdY/XoZhL5BIZZU9PAXXmWH0JtLSfBxnjwiHD8T
Y51REnz/UH4SVeqUQ/RPp/aQltZrY8Ws+yWisyfujDnr40Qq2e1xoITpxXA7
ro8rirp/J8FHrLfPaKfHG6Iz0gO3TviYzZa7JtwQZLFD+4s6YH+55eAAXBpf
iYLZFRX9J1hqYGJQAn/iHpewVPkVNP44nczRG/Q2ykyGrLQQ2s5pIje8PSwm
pjYODDLMVMGssQH+30rXgevbv0o3SL2JWFk4HcRWyaHP66V3znNcRMOKs1A/
huEM0bASj3YtNyz95p36IsA17WfjVJuos/NiIAx26Vq9Ko9KeCTyu2gVsAog
mFdWZ7JPrhLM+xkqM7wcJIz23JMM2UGlzEkclTC4FGTKzZxxC15QjH+Y3bqe
B319atMOFOX94R9XLkTsS/duV74AWox6B4KXfUj1unF/2aZhKCCrb5KZp7yF
XNM/pIKRW076h81L3uVLIDb485Nqfe+HiDSTWdAbgbk46MDYDMhWpBh602kQ
ASrOYhnvuIPO18E75RQaNkPHiBT7cRas6XErEUh+W1crB/sPLU/zXZWPkXKG
AMp7L4WkfxH24gGlqFmAmUlRZWizIsukw6apA91s5+0+pBWFV7D8WGeJNBxQ
YRLH6b87fk0Gp3QzTzldnSg+i/QGYeUO32Tur1VnH2kNCFMry/x1jotMOEjJ
5MG8VD/4pjfZG5RPaqeD/STuUxW/YYkpKf9G4ZzpPmUMXluTPvT7XPkmLFOg
0EnptBqFiE1lNhljLMZFXS3n6I3cdL/u0Bt4vxvv9ae6IE+CFEb3+jhSc8Wz
BxbdMcZ5eyTexnW/xPH8TE3S4KwrvdSBjjIbj0auJGasIiMxDjcsehK0qIxq
0eJ/pHUmT6gndP1D0wR6JEh017lv0oPNtF/LTm9F0U4I+BQYGjaWZyCfrIcn
vaN4Y21bKU9WDpjuYfWLAk7zsJaRwxIp3pt8/v3aI7649Qj0jIhqBgGyTTNm
8jTBKUKslJ1lz28GEGD/OvgWD3BU7Dii152rO0IHfI9gx7zja2Z2/5+U0aTC
a8TjcW66OjLoe6z8sCqX66in8rx4nQ2e8ZIv7PmqVQXc4r6PyPVOD2jJ5X/u
rXVwqQJHRdnXzrMABoRGjAAVE0o4j/Wy09pu/Tvlp6UcraUAZg5LDQQvirAc
MrGJqXftX0g8/HZH2as/kdtmzthnHd+WJzss1JpJ4QuVhVT4pXA3Z0+hCvhv
z0wSY+IjDB8NNB9tF9doeThE43jNYoBFoStRQzev2bOw9MB9AWpRXGWWn6ho
hZeJiyFFAAsDtL7j+8xlxuOHF6psghv5A3bsFx2FMmuvXMB9T06fOFfsANt+
FDlwlyH+ZSsBfybaDTVTT3GECNSwq6td0T0d4uFSTtcQ/LsW5T/Jabq54If8
glAsNsJg0d3OSBoWqzKKIROL+07uNogIGkIDlODMRaxCADy8eQikR2cGaodb
JCXvqf0Z57cp7xAlDx1MJ6GCo5YSSHdWoY/rRPaPxk2c8z0ZnnLxt2vyRPv/
AGXI2BwXXyqk2Rzgwx+sT+dM0furPPUeCFSzuDLXYgTAHOyV/DkNnjHYAHpa
dAaIH6m4PAxLa6iwhWoR0aiVYTRRzfrPGpfWZAWzIz2KdeSLIh82rYSQqDDk
t6oCyDFWzDu3xFMJtnTtYo5ZtLC923b6Scc9b+60ckNdmkztQ94oeq9M2nnQ
KmuSNcVVfo/uGBn4F6YwzLSohW2ijp7erE2l9cN4ed7S+CShJHOgHK7FjTjk
xf9ogv7ys8qwwrMTAethdsoi6n6p2b0GfPbJQIxuHxGPaI522fcJXi0Chtyn
UfQHH0Wvw191+S8eGyrtJezrQz1hw1VED+2eVb6I31R4luNym4/sBRjZzxMC
jQzFu1LMw0WbeK9a5jQgtx9GzIKP5nG7ACTH64EnhuKWfKEOKD9J5LYQAT6P
FJOiizALSQJrQYzHEI2/A1B/tpIRyIYBqQdqCau3NhGQ6kB4aGIne4/xiBYh
fhfvVbqWz/7eJ/+hKPNTKfSQQjNLrFqh5XeKJJRySz0/O3ilDiT+ap5tqZwW
3oGYb61cKmj9BEFtVV263hryH/XBh/kU4qKVdT5jAnWehB0o4q7Xo1gkoFVx
nGdILqqoTFLA4rubFJ0QpKxMnZNA0ab3HpEZ81w+F58BXalYk0+t+neulM7E
uMrSps0VNPS40ncoDa3uiFfUptDdpmzpOaF9A3berpGDUbQVUT/5paWMagAz
ZXN+jtmZ5IEm5/RZxeAJkkSUcgld5rnknFNuRUXq7JVYOzjppPEHjV0K4DQq
Jx0z9o4bPtuhpAP1ppDRh2xdhP21Pvv2v9gns4exWEu4vGQlow555M09br1v
GkIf9jXtknj5fH4DffD2IS83yRGzBPakkVbPebznoMRrUAnlNYRq5ikFt/R5
7iI1Dq0oVGiNoYGEDxT5Hk5UM9S6OAzT70Wc09FkEuuG999vVKBdnmitG2w2
sw/gPOuCUQwGYpAtMgTpcdnDmKBMDRkfG9bWxI11zAadENfhP1GOCsiOj1N7
R9WusHVoS5roUsSnUx2NXbTg2+QQ7fwRiRWp1nNhlG2jOcfkITBxpKv8LsG4
+NnIZ8W8fhroUtPw8eOCTQqaZ5rPgEqffL8rHz65eAOMoWgXVrNopXUYIguM
6h/h0fwZZ7jCd/xEQy20IkatrwaSYFA2Ah3bY2Q5oD71yW4DXb2uRRTSCNQt
j76wkLCqmCgPENaahwtRl3wZ241yv0MiMExBMwIMRQCEjOav77wL3L22ApMH
JTFLJwQ2TaoYBe6utQheepbD0gR3wQcu5KDYz20rSTNJzOg+jEbccC0GQnpB
fR1M8PIKyFo/5HreMPOLXJmVnn8YmBRoU5JlYxekqeXzPkvKZ4UPX/vI7OAc
ZCdbRPejsYqoUgWnsO7jhJAfVyPVf87RWrLQ3vLU1lDyc2sywtHGBB6P44ql
OMlJ/mhNhEnSrbYymTrvHSpF1Zj1n8SFL8kvO6Gjbh5/kZhk0NrsPi8nXHZs
Yd2l5CxCkpSNgEZK67BumvHePibFAvk6HSYmp1x6OAErtzSZ4PSVhT0MiIN1
qak81AGiZufv9aJNU64qT+Ou+lUEjAh0Wj8VNSExr5SI0nuT8Gs9guWnewQy
3syiJ8h4jxFeGoJbUD8xL3n3vzkjVMDfeySxeodxC+F02qdED0rm/xqHPBQ4
EmD9Wshbu2zWmgForYd9N6f2PJVlfP6pNiSM8Sb7B5ez7N505zQy0H3Sx6rB
wOWzbpNlV6I3eRnuA7fVZuAFj8AiS+UmPbkb9MYCu9Gx582sN2DtM65sOBqK
t7C+FUd4LIbJbMM0psKcEoCpnzSqEZs0NTbui3flGqYxxf4MHJQLlIZNVrkl
aju1klp1wNXRYFqzTNSaUNat5y5ijTvj72cV9mGVwn9LFub8RVrEa08ERuev
MEwsrqLrk2YNQE8SQAm0Vpc8tFugG8f0moqFmTbUVLcDQhDS29ZMDSoT1/g9
0mtxIBj2yAlYN7gC5Om+iMwpO0WH6q5V/WSKCd8XsWv5VEjaO/iD7yoLgJ9y
AFV9lRxfXppdYWb5CMA7vut9OHguSIs7NRz7VgmJz42KQ3afcPFo1JT8bgEq
iacnMa9yrYmozObWIW2rnuumoPfBFA7P3MRxQ+f2NR+Bywjk0oX8wjYPkAlE
RL5O/dk3RS7/NprjB8lXnLK/6JvGfD4kOcSaXM8xdpWVlrXygCoubsmj80ej
Z7aFQbfxJHXv6NqW2EO8pDEEht2HDTvABcBL2fkhGh3lsJuUvShSXPRGxAZ6
/6H2ZWUX5hNkec0iask1Q+mWS1vapr8186sxDv3doNo+1HKaI7tV6k17pHVG
nUHGRBOwSjW38U9IdPjKUI65s2VKGM5i9zW6N4ubkmxhBdol5e1MyeoMnM8r
lFr6yJOfjfXr/h8TtksRYmppigcFZEltAy9zxspVPkz/RJn1QyIAgXHE0evA
PFLwCriIOBoxZJT2njcPW3Auy8gtxzbkbUyrO/F3TndoF5eLuOpTqhUb4HEb
xoOTSblysdy4jGZljB8b8zlFJWQSPOSmSV5iJXJCDJL3/n26OKZJaiUmYqrf
f6Ch+Q5fIlTCduZSqj8Y2oIvFjP27aCZnHaKfP7GKVzytlPocXpUrqzm3TOT
NGYa/rUMCMHb5mZ9iYJukkfFRoTGJLcR3or/0maHC4JDVa5eimjKRC5/0/eJ
mEWvcZjGKOtiwcrVBS+jMxOZsT5KxieZjkKacbQs4WZsSErituKlIQdAIjV+
5qOpi9i/WSEiVyIm1NjFi4MIC61n6tBB5g57Jol54ZMMwQU08kTPo3gVCtPK
8IYsGuPZkF3cRAPUxCKrGuUEg8kSsPa9l80dNq50nst9+o+IzbNnoIaNavjn
UQRi1CyUaog1vv7jGntQONxT45RCDh5l/GUVpKTXUwRQ2WwLTK2o7TAYbZlI
PP+1X24iOSmdAsb2pY2B5rH8UV+EVcOFwpDU1p6nDaAKKpVwZ1bvO964B24s
x4uxw7kkzAkkT7fZ+BQVDC7NDNygF9gTphXizwIFEIAr3U7Syh774ZYeSvBN
Nnz6pJG72VrXJCPxq1SHUiLvDsrCWkVY3jhxQf61gDZudfNvBpyRuKsIj8dy
H6/ySqNzi8ryMZ3oblr4UKqYpOCf6VhveXJoe+nKliIivcP1QgEUbGYVzpfm
9odSgaPNnYS4t52+vpAoo/CwC6GUSx9SHwmtPcMNw3HOcnOQfpVxHpmfZ86P
5Zw1Mnu/3gJUtyoMHllgWJtxCJP8N8OQSfIq7G9zQvT5CZltcMD0jRmBHFGE
p4SQ8gKCeMDY5M62Of/ECzIDAnef8pRfDUjE48GqlZOo08ykRKpvFFCjiSPk
i4ioerA0093qwT3HbMjv7vpfIXxOGRLCRtAV0CXFRn40gxpSYHLhAPDxXI7D
CpRLzUSVf8bDgxvBK6GUN6iQUfhQpcS+myGDPgp4qUP2GRrHaFMlKua82Zi3
K7VkAHWlhxtRzHlvzOJcjzsJJQo1hgqFmhjnfGp7fbfW4pqnAlV36WaiZrV0
lz1NE2YL/YLTXs64R9AP7SBgucWm9fxBsx9UxC64z1uBVIrtNVCv5TW6LFqB
jPbBIsDwKH3nIILtkCP88jePepiMx2WoYuK2VGMhlXQB0YmKieBTxRejeqra
f0rdWevswadysbhhdpDIKeEKAxdSA/2v5rWPw7Ry45V4mO+r/M5nuZmmNpmX
lZY/2h2tc0XsXBzAzMS+fgPzqCn91cP6Hzl+m0nmZbRK9jwJsK+vkiV8SUYH
kkEsAcgEuujaCUXUcdpzpzM1vjkGUp4Z2WIO5HuuWDmw/0E1FsQzbVCHYzn8
cl+MMZc2ka68uPlwK9XLfKs81w/VujWUIydzCe4Vw0H/wi60BSW5M43ZjPhk
WntSWuUpQYmhXlEupkX+TeBRUiD7KG51kPPUzEOnfIM6QG13Byrv7qGneUjP
41sttIDYYOHE8y7l6vKaMjYXNj0zveWbeVwRZRdyX+609lDn8eDZl0MHhvD6
OL+XqXHowvgsU31X+9/c0NPk64rp12S/81vhinMcUTUTD09caestUqRtRKMh
7tDmgUruxIaoXeRVUgZNtWI2J8bcotym4IHd2pvxmWOnLnLWpIUNp6w5+Hx+
vZ3LuIo7bYSfX4AL0Ik+5YD/FvPVfzwiTJQNlyFlm3hcyhOqBx0ufOO/p9We
LYh8g0ZOLacFjKN0544+ugHtaJOmf41jgu4Ppmob3DdGvXid4g5PZHkWqMRL
0YY5zj62HbinivlSNQ7guF7Yol8Rpkhddiankpz7NcMy2hmob/zTHtmT8Ftu
iwo29c5xHayuzu+ak5alrgqb3PG8/oatnyKXpYh6dHWol++10skrvfDkMPRy
K/SrDvjxNd/9rDTguA3uoZ/yAqD5o9WcrtBdzpKnG//aL5Wbv+//c0CDCELN
zX6CtgLNpa9C5V/LyolLsu7YtPabPKT8W3AXJ78gMvkfZ67WRZzLpivQ9kSV
CgRcTjl/vKOxAUKmmM5CJeQi/UuNntq8PtiL7zPuVP6k5mp8eKC0wSTPFO+R
F7qQbROMBSSFfLGO0bBBcTc/OBEXAASvypZxBxGmbxB8fUEqYlUmbntRIfAf
Cj1TqkYu/VbfoLQWjAeMKABCTDnuu9B4ob9EAcOSXIk/gO6zObcQ5W2fpZOQ
X4yhh8cVhGJTNSm9Ox2hQaYdb5QIf657Y24fRQhpBEgspMGFlbwrm9UiIVp9
ok7JW3ZR3o0+1J5whmfIKtd2GPs82RHDjSUm2H2HmxSFXS7Wue8fJAruySE5
YLuWV+U7IiMsR6XeQe3CrsKKuERBDILEVLcdMr/4NIoyGElcRDMTiXVD1Qz0
Z4uKb+De+8Njw9TuuJfwAhT30hPugFsj4/+W+xN0uyS6kUhisGGwXuM1S54D
3ovxLBHXzNPFy0SKWIvLEKxq7c30NtN5v4uEHXk0zfvWGNVX5hoY9A6UCs+h
6rBEGo8PazyKypLajY4BJzLIMPp8k+qK9ioYxvE8EmKT8jPWqFeNa2FHvl13
jDwkglal1G3GeMKv/5BD3DV1SPUysOH+51Fp+qca4tEfe8QEkwMqrBRW9DOj
iUccvu3vrA7vxndpV05v54RaZGKTM0Ls88ChtuF2MzIZ17K1XoBDi/Ui7VQ1
qI6tb7AQojcCC+6I8KMNptVOyJCr0KCFXt+sDuHbQko3AiMIPbgUnoVnVMEz
R+/zGA4D1xRB57AETYyvlM+9qKZGHZXPlYohutUzr3tbh7/8AgXhnmpMuWeE
/HsbfoophGfKEcmT9j9pgR/AUZ+p7v0zdZwCYR2TgNP5FIxJ0tbfuUcp5PsA
KsqA9IfZxUMEtYBEshyFRJ7iiWZRbaC52jRUX46b/sK/UOHvnpPETVkuFuDf
Ha65aVPQS8Dse23LgmwTfCZ8SloovzJhPD5/04Lb2dH9oAV+lTQ/fsuzFrQ/
n223aolYK+dq+6ZztsxWZUrELtAOwZOktjkLewNKV84fwKj+SLy+8o+8ILWJ
e/6BtXUNNr67r9dk8qZ/bKs4v4YseV+5v8evq1LXbvJiGlQwC3DvgiDs9k+i
6gPTY9116/Tcpd2Ig773DkEr03M1lAdy2iWeTFUWwtmLYX07a6qV2nmllbjz
5SBaLxlzJPtDWMKmRlVLdFfVJ65GPgoUv/Ty5/AWcOokz5ULyRieeAYZceLJ
ozjwEgdRWnYlZHF7Rlkq1gCRPjOHcFNoLpbxYQrs1AH0lqybGBU+cun+u7d9
rG7u+grL50WT9CyfHGl5X6Dj8DQeODkQ/WaYcJdGClJuIN55CsETzbNyVEhV
AqCYyH75LAdoxUihTdH2ZGd+/sL5mW2yVXrkqpSVgC7Z9OrnJh4yOPp7Dvmw
trKQdw5pAkg8qb1jvGx2AQzou1WqaL9QAMxc+mbn1DiySEGOiRL+ceP4/Vq4
A/J6oRDbJ2D9sp/EiMCM0A4NVkuX2+gaGq1gzEQXglvRXhIA90MCzHChKl6U
FGuJTL78EBzJMpQ24k6hk1f22vc+snWQdgjhdzPFKWyUzY3/SA0RjXZUUmdx
fbCEWBGlVm/VsVz3t55GSdYZ8+Jej+J+5Kr0TUsufONvuG4trspCGMUUq5XS
uFDNemJhpmFGWjMU0bXeU1OfCFG990mSe+oMwcZDcNzLzzjx2VEKET1vzthn
rRsTSNw2fYSiq4XYwumJYBlADHJef6daO6k5djbWOyjkpNC305EvmLTuWxJY
eVpWxFAMyYZTC7pAJXuB2KEnH/Ogw5a25WKcl9ztxa0ZaZOEsImvj4hi3eNh
p1S4hdCOr2zVokaE8dpSY8tUe9n5yTAqj2rwCsYP1Wvmd86vKSKoN9TsUizf
15SnmHCTH941hymHH9VhHwX7PutJnFLZUSY/zH4AlzYZgbfdr2bqy7RJGRl/
U5UQQXPsT50BQ6Sz071T4qtzd5MqgjejtZ2hdvgAHd8h0z1DHIKjii/mbyRR
29DQ++Z/Tq4aCcadCuQPo44/fqnqLDYU1cs4v51QAtllZfAwEHo5NKbfyLvY
ysHrl/wvkvkb6LD3EevSXyVWbzkEWJIXfenSm6ynGPIQXopq8n8TpRWFPdhk
ZC0E0Qj0GRMk29bOQOUNzz5cMPHXHvF8nbnWnoG9Xzn7OcnakZ7BEwD07XXh
Gd1hbRU18GUXemp/FbBF9qXO5Q7C54Nc/w9P2DwhZq/0jYm5CEJ9AAoOjJND
PfX/TFIOdPQ2RDlZiXR9nC1dvE40+uQZJVQn07rBNAGDBYaBU3hmiiIEP7Dn
3dFPrZV7YWA6sPdU/CrVA+FPAg4Jk1FIWIjXVL3kyQzhAgT9hK/HKfJ79r2r
bS4vkRDuJLU1c7JaVQ2WwI/O5v05gEhPqjHjabGkUp2qUBtgo/D1jBnS/ggy
mfD5DR1wy4fZhY4fZmrUfJWdjB0O2L/IzRPkMe/067miskIHKRontyP1NI7X
HtX7bXBefVWDfnwHrygp7mCZvRy9KW22Eo7MRPyyq2JgEF6g+R9gu1jD/ZX9
lNSzbuPC9VVegA+Aw1oDgzLogh/SPNg7kjWsUFG4ZnDooy50wW4t4z1mOF7v
vmStTQLIqyc6UyxQAEvbbjJFvlV0s8apzkwFMJ72xKtHMlq5Z/N+AgYSkdEI
8bPW5ywvgBS7sLnDdx/wsii8e6YNOYbTs2O+ok3MKr0xMA8itJHB52wGL+Uk
xSkwOlDzDuUbb6gcyjlN2A/GRw4mEz553Z0AYDXq1Vd1f5CZ7yihDyTyqI/F
zaA5RzadSb3BqeMoeJ77qEP4IvHLuSSAVJUWisqPkPDkgSOQmQWd2yoGDWTx
A5QOBp9h3RGLErIDR7UslgNA7xtyyZvIfTRfYFjyfr5E7zKjOe9GVAtXzIaO
AZkVaHHc3sIHi/1WPUpKgPCfUdczEy55s4Gl+4+StoM+7Mk8l/oINgaiFdlm
QYQJZ9nsd4kpf+WVOHUzMeBn2IwsqlcjIVctwBjyJmfewN0bTnuzcZCwWXDz
7nQUYbC5GnxWi/YcuqfYULLYvZ1h52ZMyIc1Zz+LrZYbIXMKmALzPjhnGjr6
VGxj2Z8ou6dEhou2doPUSRHCwRUNEkUPhhrAZJVho/9hDAxlLqipdT/LV4uo
fMBIHxczRxtwN3OIGhuMYXca1jWlS60aohNhoF97yuEl0z7Kp1xEV4WQyvUq
5IenNP1cqkasgwuMGl0L3hFFNv58h7yjXp2V9u7Lc8uyKxO3P55mkaR8HHo4
I+PoHUknLkLfxVDdI6j8Yl7e0s2IfNDfE438xUfLCj3hNaSlWQBpTXu6QHCV
zDOBuaQwkbUs16WwVHnl/H2r66421zJQYGB0Kb0a1tD/4Iwr+Pe8KvJkarkM
eUdqnMCIvGGfqRkv4PbTn0nHSEcpxFp46DNbneuA98v/0kidmnh741O8Du4k
QmPmDKO579QvDLYmHNxV075RL90BMrR6bG9PxFdPCzU7iZwwKPZoQM1HrVDv
iN3ts1VZ/VKn0BMR65U39GDVqGejmhRvrTzDYRMsfwVxeZJE3zge/TzYW1Hl
Vq8ckXl8Lh06MCKZEJ+1OxF/K8qZPyDpzF7jFyHjvxqProTjjn/CEowUWl4w
cwc//LWBC4u/HlG4hh6BN5Mb1b6OXACc7c47bHmViZ2kyMjA0jXwMILjN4CA
ZUtdgOL9Wln19QLbM5Jp/5zNqbLimAA7m7pS3ee3Q8P7d1nd9IJgRYbcxpgR
/LcO8sv1FPHIN69IBtwVX9MuwXfyywBQt4F/q03IKMi2v/T2oYhFR5uQQDNc
BI14Zi3L5OGj+ps0p4a4NK20VUQvqIHoJN+xGEISn2guyV+Z6jcpML7YMEdX
vkvw5h26tJlUjmR4E9OYp6OIAUSfkzw0noFPux3xdLA/wf7U6BNm48qyC2mz
p9HZ7QLg3wHWWJju7bX3TFlllaFYpaV3M2zDfikjlBtW/3T1qLbRDeqcGTIg
yR8a8UU5FmYOM+TIfkDzlQ+BI0reiJI2nMZICZmDTIMvLadfDluuR9/3oABr
SZXlmvJVNU4+Fe2fmQREMF6O28VHx2DLudElf4l2Yi/bK/UNJRZxB85lwvZ2
zPrAihnqERzBmqm2qkT0ss6wgza+8Rf3AC+HfE8G5Vkn8bmL8rQSFhI5cyfg
rhvFS22d00csGFoui8q9mDN4ODJhdbSrj2PaemFIrSqsPsHXqXFiiceGD7D8
5Ki92W0XWNmqJhLMbmYVx0cj4ZDh2Nk2qBzIX8avg8WPW4AsgaF+O/brfjd+
VxC00yOBgskOQ8SQJISWVT54G/xJmGwXqR7c13A8+1XLa3gMCSXa8ONopUOn
6Zo+FerrvNLi8F2aMna4C/7dLI/20D2Z8h1TbtcBCoHtX1l6rGt8cU1cPJHc
z8tGkp8yBXMLDEX/ugUDowrrJWrsbm6s55bkIhjt8s6ofJvagh04tGO0ADTV
xrZasRqjd3/iLJ7VIN0FUzazGaX4NMJyOEgxyrWuQi00Jdcs0iXUovXZdRC+
Sux2gDQPPAgsCYbI7Acl0df9+BMKQFvBWum4zJ9ZplBPyKgfLQq4rHOhVu9o
Wr+JIlD4GW1lH3xA8f+wcjgsEmfaVKU/eb1IAYBSlcDQrf7pKm5c2UhtMNpk
oPoGfh0T2jsbeGMRXgEBVoMXkClfT91UWNYdbDuZUZ7Mx6v4gikwg1aa3UTh
d29VmByCeulDReiGM90Kl0RD92/rr8C4knDVkCMb+e1cUgvppZcSwz8F8NMN
8qjqZhzlL6Q2+i1/wK2ztRGNgIOoVMhFruPzIWOrg9WLC5Qivfql46ztCZr8
Mmu5A2siGGvOKiggUvB45NXm+SKstGoa7o4VtF9Q7MqHqqKuUJgv1l67BL56
lmS5cx9icxedepwMQn8W0ANNbdCDwrKkc3pOUzTXCnBNgoDDsIuUqX48UsFQ
QBhncsEJQes0z2JN4Pf2GHht/JvqObnfJVWfkR3y18uwzRl43bpTlx+j1GUO
TgwHMYpCgQvmFueJ2tsjOgEn53OLLk6LjdA/x4Tj6hA9IBVXYkPHoU2uuRmE
UNd/W729pm0x41ikEKHP6ydY22K8tfQDGKmhAWCky/+jMMUeI/Bm5eFHGMtf
0RR0wpKmhDu/ifcBL5fu8gwULn1+2varhMw2Y7xlQYLvvN/MUnNzhijQdzda
Pqi+y3+8IyWA67WfGdQZuGMHlV6n3E+1QbyqCLMmVPLp5ghxh2EhUbpdVGuf
OlrwttPnxep2k7eMPiGz8CanpfECOsF7tH1qohay1woRkb3Dh7pWUhUP4vq4
cWcUzvINNWdhid6tVlUWIYnrIu8EubLvzl9vYU7cy8rLVDTXVKOeSxG4emxx
jucxuyZa3yjVF5s6/UTZYQJXZI9UjrtwCmOODr3JtGxUdBgTOTxf+BOGJCGv
XeLpZ8vXcWyJxvn1F2KPIuKTPMphlJWAzihwIxVAwlkiWvNJ/T3OqDY6jR6m
MkFAaGQ++w3yPzlHLNYtuuMroeeEnkZE0s+Ieh1JMKumvIbG4V1wzEuJ404/
j2LKm8k2v5hMCJpl/rKZ6KkWo32egTQ72fGp8K4HytoumXJM0MtT7V7dbd4Z
ykUyGi3dEHqly1Y6opBeV0c9gxMKpRySa3U8PLMVl8CvW3KdZ98Q7UVatq7c
u9P8mWNrjM7veiugR02sAWfy7SwFoMX6SYc9mEZ1y1W8PEAHJNKEOdU9uQTU
mkeRP/2prHfUI6+/RIwTOM1VMXndGFW2u8dOVnyHOyYhOwZhUSUlPMRzROKk
+6gYEjWAhNonF5ZBJEHY3ZIvBeHVNE+NNbe3NLg9qA1yvV7TBfbQK3fTNriE
6HfYcpeElHywqpq1tzHD3n+E0n0voRXn+PtxYZv9U+OFU0Nk0+iyCxC5iyi0
T8avE8cpeVnncPXLPMCLIFwUJw7aPfkEPkSo5ocvr9sTLSE4EjyOwKNLcdJ/
mqjHyyAFfBZzjuHzqvwgeQjlqAT4FFIHi31bgWghHgEceRcjxIpEqvjh+950
SkQjeefmhCj6cQs8o/rf/YSnkn4BGx9hcDXtry6yqj6R7S5KEXhQq7l3HKw/
E9enNe9hLs1c8CdS0TU30M7wCurpuDxx4eMyCBXCzNRbzzOjqwvaIUzNOQdO
h6CJKU/2e8RXf/lZRh9tf+AqDkak7STmS6K/kKFlc4bopp2aXtRXvtZcvT0K
wizyDQ+2SVItFhASnrly0BMTQQfSy7OsyaivqADMBOHbzXQnX4WDY65dkpL+
2cUVpABQX+0fBAgu8REM2ddOCq2VqXMX9tNQJQ0hC0IQoJu0Ak8bmgVs6w+t
Z1KybINsjAeil4bDTyS1L8JL8KJFcgXX+1KdpDnAxIsSWc8xvdYMAC7z6a9Y
qHYaAStHjT2wAiewsQ4+m8NCbeh5PZMp867wK3iGe8qW4dPotTYSbCd67wfs
tKaZO1uijUujwc+n172ivO0NoctO/L3bTAYManRKJbuCom91ZN9MAqPFcDSN
weBRGYW/Lso/5vdqFRoDiRw/L0LdqhRG6n8LorKI/Q2mSNkWCEvExExey/ht
bXFGy2LJJbPHjrEy7V8MG0uANfZ1yEfBDXV6zbMp0ic6VIvBGDOIFqAAunXi
QzYwuqebX607zXGcvBFIGIPByblBUEDMUmVA2Pf7FiDWY3DKDZpvWSe7mj6y
fHnxymBc0WulUlgH2PudGhoRCLHWXz7fIW13W5CofOuhf0IhiEEt5q1HbYKF
P7eUp5xASeULVuclE8hdvXCjm7T+kjY1pjAdfZD9mU4Vp96Y0usoXkXg+R9A
Lk8iDNzCZS8hMuQpcf90ma4Kus1fAN41SEB4PVlYWbzQcbKdFSNb62nfs2HM
nGM8LOaOQjbJcBlVWErws5pNY7/BEKwqlqm6bZ7Jrcut8jo+689I9AOVYwGa
snvCMcjyPD1wJTreT2jDtFW/wfWpQI9ArTVoNosgzKnR8uivwJ1ZPA2FMUHE
Rz9iXQ/ZBfVX3CiFrseLzhQAHDViTXmwFdYWE2eUltesB7E4xDgFGqHKi9nF
Smo4EjaTq++GUI/bSsUeS52vJ6tF83ucUe8q8Lihkb4nYlvRExeUk9+lVOza
M75cEbkG7OipHiww5S/qm1AFEcdOac3Ec429hltyR+r/CK/6Rp7o+sV+bnRp
QZP8p/FzRcIML4VafzzXzoZxHHT7Z5MjFFtB6Om9JHDftXJ7wmVpEv6YQzKQ
vFEhdNSOqcO6XJy9GD0jaL9jPzRHJlKJx9VAzXUXbb4os2JbrPpuva8iHqPW
ZzkG0zBrXzLOpWrA0N4l+xdJayXTJIjTtywm6BGGRsHk1hXkqB2yTAaZe28D
TmteSpG0x3DCN5hBFrsdap0XdQB5gLRnScjMTMYWJHEtaxzDccAcyeUSaszK
d9VTb9nSTGAZIegDETUhKtT07ucd17dNjmjO+6GKl7muiN5+5kn9kEb8iUW8
fRj60jQTTSAczGCvBCqvRqO/nI6+3/9xLLOJ2Ozu0AKy/v8VR67u4yvo64Al
RAumJlNS7bLKoRqUc8QTMw8f2h9fvstiUQcd+K5EKoHAzBFIL1l9oPI8N2fa
5Jy/5wabIcwOKFzVlLWb/mwxotQP/C9HuLsYDCnQFgEQmC9d7C8d7YWo5aHs
D6miZ6mZmTIwbFVyqoJ2pYHskP8G4rmO3Ew/KLUXynpCZupUyrWBeAG2OlTk
PmQ7n3Eg/wLNZYy452M+Oi/0Y+8qxxZA0aKinV1M950BCmAP9dne0KJeAN6Z
f8gAnHtoxD94k0Yj9+R3QjywGAQHMPtsviisIH/OHEqfngsYZy9sonXV1WE9
LW3pXZZ5ketHCTD15O5Tlnqo4XMaBCJLbMAuF/3wXMhwGtmMDXHOI3UJ94JK
Uct5xSwtYPQGJ5JL9qBLxrJvOIYGRmSoUgwIawVx929oWjWHdYOI3srZPaJH
wc/+h3FLp8GVY5GHacJ9I1m829m3h0hEOTezXgBBtmieiX/tXHUUVyAGP0eQ
l6cnEzIZw45tcwV2CQw47i4mljDzXl86quouL95yNmMMBsD4KjIPT2QxlwsY
vhwEhcU+o2gQMmia4ZGrd7hBZbNBvpFvyErbh9pRgMpZ4ORa1vFlus8EY1Ri
pbjicsF2FbezkHCMiPbQ3x606i7ApXxtwzDxhmiDcmzNnihddXPMoP980Fjx
uo17jt6V1VoFzldbtSZSHuNKQNmj64FlSa8/Hio+p8mZDQscp5b+XoYE26dz
14mJcbRYb2zVVnuArk6UivJoHS6oVhd7WX2txCQ4OrI7uJ1d2udwXrrsYCNu
kt4QbIACyIkGBGw0PIh9beh+AuhEs0LzJJxQz8Xu930hqmfT4J3OvGPlGjdL
j+rmo7nimVR5Wru83z3WSKdXn2M/W8DHhtoXiQt6HwCoBRb7L+ibVypR8RGw
MmPhE2Icsx1NVHsHZCULNmMsbaK7XDRUog6EsvYI+phV261pjUk833eGHlXf
QUm4LefwHH4plYJPFnHyz6lQ7H4E13280/mZNypQvVDs9TxUL5xqxzx8CIRn
cKhRdWXQFaJb2hagWdRt8RtF6uLqj/n6b/YvXXS7L6qWc21rT8fay3JXXu8Z
ZCC2LKaqvnBkHN3OpJ61BMU7cJ03tcQ0cZQPmKMVj6d2X2KUmwhZ5KyqTDwO
jlHxYGH+lI430G+Kvzw04uwpmHvAQIKNU2KLvvE1QXNXyCzMEOpthoMI8GVW
hsp7GZifVO3UJdn2BoPqX1HBus8gsA58uUl3BCfE2gPIaCBvtSs2nLsf7ePO
CSarQs6AR3b6NNXWIeP2AvQ5GrhuK0QA29T92kID1qRzH/Zog//JdNBwnBVg
+YAb2DiQBkE08skUk/uTX3+hB0kRtEFwkt2aVWh4DXSX7kFxzOUUysx481bJ
XLCcl+/JVMp10pYNj73vriK786wV/TdPwqHmOi9FNaFO7wlxaDkD8dJoKRn6
chMgUzNs6J2BY535eDIQxLv8s8208WGTIOuwvNsyeUN2fMf0K6ah/T6fBq/3
0lc71mXWSfnuJQh6Ng3SFFQl+8Br/DJ+BIE234m6q2TrcK5pyXvEwzxA/aZK
21XudqwB34Jelk/xPypmxiiVtzt/EOU0jc/2K4eUhtulp7jLGYoM1mSorISv
sxh+HZxxUuHSne2vO04iiiIEgk/Gu0eoIb8mvSAmU6eqqRqGXpH7FS25MBEO
cVzvMDF/P2/XKq9Lrb5WDlWQzcu5QKSqQje8cG8hKJ+GSbqgyYHwY1DVGD6m
RMTPRD+n45NwrnpjVq/z6ff4ZZFKYk03ajGRo60Fh99y3Arrq4GQPTg18oBn
Slq4dLOSoeuqxq4GWUDbmfDHhHyizi9EH5gHN9uzGChc0e8FvgxsFx2Po0Ga
uUMdLKXfkxLACMezjy9KqCTW8Rk7Q+yATUzdlCQsDzQS4ydY8QOcBV0gA61k
Tv6cn+5tF1xdm0sTsbg6eu7TvU4XGoDnSHdZ/5OJxgVL8Zh3m+WsiCV/M9tT
zmIcgr6YxrSQMwtunsHwxeRq4QPUQoDrjc9dUurrlQ5aeiD0ByxCRmUz3yiX
cXoR7XU6kxvcV3sWi6cCgZqm6RX47AMvxAkOjWKzqiTClJHPq3x+Pb/Rex9d
9K5/jq9po9nEzFF+94VwwxEeNq0mGWHr2P8rI1Kn1iYPWQK9t5qVS0reZ6v5
6UuxSBAucrt07FHpwrPqPE9IOMSJekSm5qP2ilcUPBxgj0pXdvMZUSsSlqaB
eDSemyWjqkaygqMubW1EJpV6uOh1ut288ajfuROkge0jfiQYotypQsJpZNnX
O3r6xFgimaWCtMJd5v81DcZSwevPPf+PtTw561c9Ydv+xKm+LWWb5Ytam+wJ
zb4kC77bJO5Q053s63sG5Q/1OuLDvu63V4N17WO+FX9+6KalY6vPLQyGjSf5
CN4LSu4JrMzCgt+2L70tKXENhwzZufB02VYKKre8US/tTjYfZ3xHxslMlv/i
SBtzbv66LRcxdZBQKWkoS8kxwIzsgpfDRtcV8i3GNYzEyie/O69qYrbbYRmE
sKd5QT98a1zogfyGto7nS6VG9Y7VT5sStaJXZJ6ly73ZW1x0rkDFMlJKtReD
PLfhff1tdd/x03HwaWqVZ4Hl4OLM54EO8O7JtajHJNEl9f1kIRAwkOmuVqMP
heENkuaO0QbJa2KuNDpMkjQ5S4Ae+61ObHFRtbTjt56/aq34zsfvGLTp0Mba
lCTDucLcH/Yp0ZCIQWKSb25gpMUvv26KjPp56PESvjDrh88EChEkG1EWCex2
IRHlN1l6+JTpXS3lK4ZJAO2vANZZcTSlRWTMtjsYB3Zf9nuuDhECq4Zdp2Co
EAD2XIdk4EeILXrAZPajULzLfvwoBNrgO4i7r8Kd9vNq/SSzHzcJO2yw6z6z
MSv1VTgRbIyWVpbkIZt47nabdrmA2a76KkedJmKxbpoCrCdVrjmKetE6PLnx
MBQPXfaWTHk6q2a8cU/B3j/a1C6nQwiB2G9qXwLwSZtWuDAzx7blNhhy+Tfv
P7vKTPfvVRdxo1LD+iowWXykn9BXkz3o7eKpRCxiXPXQiSddcJqUCEkB3XRI
tA6nxQcPIL2Caq/+r/FShaL2BOhJVIS86/1w92iqL8adw+Yi1UWyQUljS+CO
PmCNFpZsPKtaNybdbrueJYj7V6+emM9Pb8ozAaz6IBjnITK6rOzpmDd0d8B7
026KDRq/t70ZDpwH/7/0LCRyBxzrWcMC7IQAQgYmOXh4a9tmJUbdbrTwDRXj
xc2+PrdlunRsDVSUMuDqAX56D46Z9QwuyqzQlT09+LPmN4JESXg6ZWGupVva
PdhYmlSDUSyBUVqH2+SWsmW54CXSPlsCsrjdz08NhM+sJZHTqq8tQJGTQbyK
dQJThmFYDUx2MIn1o3W0ZsCHSbaV7m50dVuhzTuK2ZYTLNIPOWRSEWxkcG37
VHQW8xI1eXNh9BivkUGMVRyYp9xs0nFo2dqe4OLwHxqoZVB7gF4PtaK5T9PM
FfInhVgXhAc9Rf2oFfOF8Y9libk7ZDrBS+1j7vJHJ8S/KH9sr0xOIZ+RT5gy
vkG+/TYw/EH84wW1kQsDNQbuJU0P6ZVC42dFIM3CMOMV29PMfoZtihyAJZT8
dKuX2+wjpyymNXWZneF2YvJ3x21bk/HIuCP5T0+lVVSf+G2epDmY/GEPeaal
JquOrDoprPjYx0WMyaQ35sB2iJx8CLM7RFcjj3Fd3PlXpq9aGyADIQh/Z3iM
MnQtfvUsvcEb7vDckiUIDbupxTdj4hCj97NORs/XWNV3YiATPtGZY724snZb
gYnaT2TnCBuJX0tANkyKWnDLbrhfR2sijNo2lftRSoJigkMLQVpyQCiOTUW3
M7sse+92wsXIJzx7yNIe5ZeRhD3ro5etjZrI1axFImXvpkQEZ15M5eeqSFPe
SgYNZk4eR4NgBpyOVJEHgIUMC0mg0rS/YbgkEIRqZOuUo6sVoZXi8n+lVza+
d20WsokR1mJPTjae9WX1WGbagsqbEJMowL766EpwjRJgZi3iU+ublpDqSczj
fQ7xx5/QNZVXWw2b8tGtvJqW2nBZCKz7wl4kGudKDI3z4lLV0nzmjbWVndcI
VXETQuJAtpwTNZIo0WuRTlQTleq6586Hm0muHmmgFc2RiYMYNGUai63bE5de
yyU2ha8BWEdt1U68sm6+HP+FyftUEvaI+sJqOkj0zu61J26sarkgb1VeM4qE
TMfqOdV42EQbNgxv8BMSF8BMk77t+Sgq85dqMGmKqy0qgqPEpYeg/6+nYSkL
jzpm6RwBnE2jhwoNfa8fVTc1yOvIo0g76QBFGM7Em0IHyTvEOgCYQdveSuFm
aImjNQ5asOVhn14ohxBmWsEGMC/Uus8rr3bUCJOZlKb/Upu82invVt1n8QZ7
7XfJFxncwsLZTMrHhf6w3BedILxgryGbJO/rChk8OwMaBO/B1AUQMIdRGeWj
fl5wWDGGncMpgviK9zt6RTzYJcMpsOOUho9QAbwYN6aHx23HMYFrO+yRmTxX
qBDxeZX9/FJ4wk73cTwZquhM9/6GWGiAJv8DduW6YUHvabn1z6IhP/MQdd1W
FMgDY5yMj24rUMNm+11YlJDkg8MScz16BcwCkZ2b/mYOhbzWPL5elbIZyuoE
6do+D0ku95x5hM8SrmRGMp59opouRWmWFxpyIfYUCvcYVc+hvmEB9N6kI0j8
jSfq2gyzpN6uVZEnw/OUMAJJPoN8qtSoeGBltyd1zu9Osq6vzfs/jQJYVxbT
xg4QhHtZdzB8QnwsqiEp98J1lkIftcHuejM5HwykWSAZvgzpZk1+gSzcr/4T
rLOpr75Om4GYGkm/WlxeyjD1A9e7HM+Xk6hu8mit9Mn2zVBgvB+1ilKTOjKE
aKiunnkW+g/HZZrI2RtBIa/ThqYeqUFbn2NieGBfY6bmEZWtTy0qCGuMW42M
GnH61DBCTkJ2oCEUttcIIEZP3Gnvz2N6fH0GwFSvZuLAEIPpSq90P8OHEseN
fubyisqwYwzbL5iQ0EwX02SF8EsIEGRd93fmAGAbmWIjy2/QAtKr6eJnoPol
okWnFXyTGpHUvxRxWxTxWOOLQvNxML0BYGRbFTEb+ZE/HK/YkedBiEfc+o8j
0VXSRhbQhguQAg5NipZtbrg9daCV061nHRRf6FX6WKJr6UhJnxs1mzG38EHI
jKaRgPxM3J2+rSF8cu/a18F1E5rWbyO0rbnXHwXJMEiONYCIQ32ca5HFvUfr
s7XP7zagXESs6PDNaCGLZUrHNWamaH5fKEihWmad0s+3sPdqgy34FY2I4Qn1
UQ/tMydRJZZKDFL0ZJGe/iV1azOYpBs2T+BqemcPlkcAU14Y487Hupf0EyHn
jNkjTWXv59I0Aom2rd9RTWs/lrgxlQGz5agOQiVNeVUZbfIXIJJfPnNaCWtc
mzpXiMAnyGXHoqpD7fx8fwtOOucytTjTG9y0ll1kzplNAT8Ak/D3PnRQwSku
9thW5Y+Zqi/PAXKMLp0lN0SuGwENNgU97Si18iMzYSRhmpS5KlCTgJTXYRee
VcXA4hFEANdmJcuqs8ybXqOc7k3aVxwwE5dg3YCuUUIxD6MiQMZi4EEuBOyI
gYwxpzYsORrGBpSEleZcWCHdWuD6eu7c+ogdGxxFB6qgoAvUrqvs2BPRPArg
nrGBTZt1YMTJxpEtzxR/64Tyf0RaX6MYMt7H5N31Hhqk40DBUPEwJMfeLvBG
uRSeRKkHVxLGkMfVdnyvNH58Z9LJt82d2v4m1uIDPB9XyrbaaYuIqRtqMAKK
uQ43w8oQwU0fb02k0Gkr4wAyIbR0SWcVoavD30NBaRTnusn+JJiryUblxBF3
Pz5L8NLTipaBFP1ccT8bei5KlyAOBIdBTRjh+rraBv0wDsvHFfC/s83uBaHP
DWswn4IAPKmzoexIzDOBFE9sbQvFEkyRfZyAvYhlmRcofqXLmjOGlhROnKTE
MMmVrNY8dY0q5ns8FppFJthJ1nQ5vcl9vj8P7VeM+lom+41uE5lxHL0UnJGu
xCX6WtgUgLqTpUO1OPCWfx2i2JEezVQwboxbyg+mP9F8Vr62++5thY8RFMzb
Er6tL4dA41t40bUGtBkK81XUVgjHqjihM+U94+Tq7FqTEWM1jKT+9rtxHp5b
3Upjfud5UiIykNx76UtWqY8riPgheGpyncrtBF8HND3RdYDT/48a+LfI6LX/
kziTNbd/kJQLpCq0bw8KMvO8ZovSsy/iJEgFPoPUSKe7nHZZ7sNLxIqbJM7J
qfsw/EKh53PTgHaMj6cDD2qgSpL7gRHeuaEEvJJ1eZBVVIrZU0MZohfcp6dm
MRRXGjIQXZtIrqSMQHuYSludPT/mYXrz22Ct9i6t4jPzzf3PBlVJsWFzcPI+
QfjVaf+8r0IWRuHmtxmxA9g7h4P75Rdw/lCqKPtos6/f9f0f2K8cBWhqIk7n
iWr/7gkvu6KkKihCmboH1ncnfQqYfhcHPn06gph+VRWOlRf9SX6RvIIjL9Ww
6DCN3cgPpShUnxxVPBMqyEchSCS5pdfGT/0bLBMfybmo8CVjpYqKegNp/R9s
JNJ7jPo2QyVUl1dZ64oWCFiyO9StRCEy82yRN8CHOHqwAHwyMUzig7IUJY6K
b5hnjkH/PVPxjNk1Yk6nTw6PNu/hH+IbD2NlGBXZknjxip48pKvinmMsXNGA
MS0sGbC/LSnsEbmqh2F6+MFNBsSi3Mw1IqJ+YfnWeZdJmlzn5Y/uMJfJa9Ze
i9y9izQV9qEqDBmSyZycoMCv1WvnB9FQwR7I4UbpN3uqiSnZP2PXyGD0znwi
qJ/jWe1fiun7NGYVB0f5sObZQAHIG5cjwameZPdWQum9an00IRu1X17hPrK5
SlTmzg4Ykptd3AjM7ujR6KfuvbI/ky/9HNc75T0ufJ9aqJtwDhJqjQuMkboy
z0TXPk7syj9Hh/lj+k4bFQY5+eALIFSS55id8D8M4ryfJHAZfD3AG/6cLarP
KHoH7uU/nV47aOQwgtTRasTkHLfcSR76J0y8febd6gV+EbmjcR/pN0oacDaJ
1M77DBsC+6+iHtW3VeMaLA34cSN6ERop/bGRG49w68nyw6Om6dLfpDRD5Ql3
nvo7BBKSjcf7Si10V/8AGKS45h7kACbnmhPPOGEWlObQD0+O80LZusIQtnBc
6D8o2GAnldJKUz4zsRxFOigmJfRGAlDXfBaDJbsS35IaokYzPpqQHgB6QGHk
RdexMXbNhoFnPVbLlcqc+QpU7hthiVBlJBa2X//X0ZBWBY/7zsQiMAK/fkI7
STEoKpXTSJ56sFXVzZNKnZbxtnWuvWm36jh1npUn3u0i5cQruOFI6eKukrPf
QccCmXnhuhMw7Zqe7ROK/OgSj9XIsXTVBB3EHf6fifaEj6USx69GkGaJHLcB
PYouo3h8rWoInvy1QZZXxs+FV4midVouWAOSU+2dCJMoCZo1e/bVX9Y8iczM
5iIUJOckwgjkvb/Eaa7aTy2bHDqCCSoTWqHzfhOp7UVf43AVnATwu1u0Sz85
DTD6li8JLCO14eshgSb7aIXawwa5HYst3wOL9jNw//hzS7bOXbWkijCT5QFj
z5rZC0v+66n3dRie2cP/s9DDVB038PjUfiH4CjcLR9W7rbmTUb0KAHuyOjf/
jbWyWqtKHNSVsmlxKkXruhjLrArV1leCk4jZh5BmapP0142Y7vLbpAPZCJbr
hZ6YOc4n6XglsrWHkuTQ39WHqj95f2uV3s0SOoiJnWCH1A51TlIhyk+IRzUF
KACeAqDzPv5mHznnc8kxFmfrQ5KQyUlBuJWU2649m0qZC2JUDk3xZf2Azy71
JSu0zrl6bUnZbK96kFHbp10CU2YnA/a68mFESF5TEgQmsUEqjhVucFN6XD50
uPYdIAUZ2EiUSRR6sqIY9Ljn7vywbJ5NRzJHavYUQltvhDS1ajLZs4pXZ+jh
hbh4VTlrAOmApYWhlDCEYZfJtOVS4JxUwHV32XZ6NEZUl3xkXScz+O6qK3ZR
ogcLg2MbBT0qAt7SZifu6BP2xSqqrhfQN4Nsu8cSpgPIsRUIGMzxaskx//UF
pkKjf6eD6sTg65Iji9D8bJIUYEm49uQR/oW3m1HM4uJ1w5Ilhx7sxHicoqjI
Pjvxe/QDs/LBTfndGS2gbdwOUq8GxoAMXTvACI8X/cOgjcufkYHs18z56Sa5
dUckdII618yGMHN7SHkCPO/xmaRBvYyPTrDyJKExoAx1KQfgdoEs4G5n7gcA
TUbGLvnbSpdG1tGh+IxbnNSfHjhliGWL+qUBfuG6s7MrXa7qk92LsO6Kcw0d
L5XkVmWQcZ45JAskuBfcxNMAcBcTUdB7zo8ALTCV38I789U9PCXtv4mYkDPf
ytNOfKtBncIBZVpF0V4hOU2Z3rVqC6LJnYeUlSSRUsB9UXDZiYpCx/YmJRD0
PF58axA7n/jBH3ZoyjqtvdhnXzYQiyhAq7/dPQaNskiz9qFdzitgdXLBkN4u
0atfmRxCTa3Dg6Vydob+Yxghzd4kzfqaeZVqtn2J+QjTgGNXHtQnGUkoESkF
VFHscIhyvtNBSVLdhwLZPyO2UnV8Lp20qxGDlReXtZbM5ZuS6z7bcR+cerll
sRS774jLscbrEead/cyE/fJkN0f4IJw4SO+6zjj6H9OVvGBFWY7A/Ss83t/H
IOW0ywSGPVcVUYpv4/poER97UcJHwrcfPwN+jGidyCp9jU5mxnEyljNIibhP
Nt0r5MMFzCYeofVB9MqBOTYsL2vJ8lMiCBHLg+Due3+TklrWirGCqN21GTQm
D74ejOSr57QXDSyW9mSSB2Owxg68Wyd3BV/IIOol1kChK0Q1ykWXQ7Bi/j4v
IEC0Y0NF1pd4HWSc0qyYT+0Gg9LfTFSOv8ZW8eIvb1GVo3/JnobNWa65holp
NGJWgp0iU6TYsYaLmM8fTvytE4e/aly5+cObHQq2XynIflYaZB5r4u82hLPb
qJhyZJQts+LacArWAH6yKKiM5fLtzQwB8u3TLpM8jr+9RDO4dxc/Be6ZwZUz
k89FR6g8mLeLFOVTd3612EKZZ4EtPxdyq3cIgYCShu+9xTqSYkoBLnKMZ8Ci
DGgvsjR1QRhqoBAJgxeNCaxZrUkRuUZ19GKQSvy13jC6z7IULLMtJe43tNWy
w5xTJl9f+6p0PUONbpXIouuuJlQ5Zgf+7k8BFoDM40bUy4kCnztbh9h2rKNf
00H17gwTq2UxSaZ42MUHGJOwzYF3KBqbdOHosw2eiGVhFro3TAI6N473BNIG
RkuKOtuPPYZkRS2aUC4sOGYviA3mu1fmCaFDH2f9tRQX17zhhp+fsDyrzoD5
47e6cVitxVvqspmhhBUk0D1s3t7chc9eUNMzLqyZryErQya61a/YO9W7f6JS
3aWwRkNKctbsYRObmZQUgPBI5okBvaeyola4MR+IiGRdqH5AHPQk72+eH3SQ
Uz7ZcQhS62obKGkHE7NhjmienWf9f7Xal8CwUC/KchmQ8/fK+Jjh7qO88yQF
YKmZd3VyqFeFz5ESagTFe2r7h870bYLj7VIHV8Pe8pTtvuhknG2pjW+uyuUZ
yJiW8GkabEIuqpK4W6QFvFCVe8zo7VFxQd84LQTSWS9IWS5z/NXvFMpayhDe
AcxC11zoF39vYPGZQ2HMw/n1g7tt+s4PQGvKJeawsbRW4p5w7nD1oG9gVnY7
pomR6x7OSJsBaSRXqeI2/mtM0HLX3c5znoetNQWVkl1lndMUXMlHyjz02r2Z
mCXHzkwrnr0BuYXpi1lGNFP0EGc6m417j9NYcl9+jP1mDZNEnvEiWipEd3Av
27zeCNkxLXeuAPkk29/0RKsQavZK3rAz3IrmfLB12u2R66ru1TcNTiqay0hP
rE7ST5IIXEtMESQFjnAHLPTEXbupPbvhofId2apJ42HsBlu9yU26fGUDJanD
yVaAXJlQzH7K6CjqMXua0h0bFhULAEh3SGKdDieCkGx2bW27PkT6qvaD3IK0
/dOlKC+ukYjgql3ZnZlh4pwJgHbIGgJ9oCUT1vfYDdo0Da9hNj+U3vc6dvcH
E9HTSgNdAuBmm2gixQ4vOHxd+2O+XINxo4ELY3eL33ojRX79VBMzjtdVdTdl
egbuEq4lZTO3pmZC/Pf+5RpNylIhVNjhs/prr2Cxy1z6mm/RvlrXXuTwaMrs
VrI0XjVQLz7qSZ3Cj5Zza/csp0jhKyfGVoFcaAvQfKZMKzQ2CEa5Fu8GetEd
yl2JuQmh/eJxLPOsvKzOMKVPuH5sliCMdzs5HeuKRJAn5z4TEzjJF4b/Wa5D
jijfAy9mUucyMtyofx74WolFjoig8VIew+3hjqxQAqCOOUGrC+GRbwI02b6Q
7OtVz2L/5NzjOaPFedS1j+2pt2mxXdzOzAq5sckr7gynN6P467mTLGSfBCCT
+qWN1wN8swFg/A/Jgmzzmi12gWo1t5vNYu9vTPn91esXiC3wtBD7iIsvrcJ8
I7lGp0/7Y9lspuv0aqx3nWkydxGo9GnCBHMVi74SMYzgpavIf6lXe7ZguCHo
k+1IYgnnla/YOqbO+joj20qJir7luNYQyCgtoIY3kd9tTCrAg7OPVdefvMrZ
5L6If4qaW+zzgO5E9wp2uBKAKPJte3ax6xElEqk2j7XzJDSqGHB+bdf3NSXy
K9PjivzWBhhNo6bI6ljzoIfUexcjD2OoEwPULuuqJXo4bQwSufuMgUZT851x
dRMO7YxGEbXeesnrrZHvHPIF/8M7htg+0pidTrsk45Ik9tmd71Wvs5vTAFov
VW74we+vyxNeGC0uWNcAOmhap35LS26t81C0aBp/oMFqRF7bfUhXanj3RTW5
uVUcN3CWemmOkDzznyeEim0FbalD8ZB5fihj7vqIwLVTeBNJn/1h/CCFmRds
fT+0yIZHO0Uzn5HzSgSc6MeGHK91dazNTZ2te1zzL8xbW1Cd+dcDWUC5+HBP
ag2MJbcu7WuPi87hWglcucicMYwCJzmrmLji2NlQlNfSCEWvtHXlc22tBhHs
Wcixo5WBQVAr0p9RldIrC5tAkB74iBPSHVCoRpOMxCqxlDhFbL1wm+Ns8ge8
WiO4E0YDP1hrE+Fu2O/TjQyL07o6IUbxv6pa2kfJ+m65n0+V1x2vBtkfJknc
QSFx1NziT4xSKWRybmy8+xK+NxxuIt7YSJxnTideo6nSNWGFowhYYgEn6EPL
Ggzptjbc1eUGvTm2cUTO8LGsmlPBhc+bThCRiUH1Cx4wNN94izKgxL4wePrY
KPa4Pqu++N3ZJJ2hNdVnFep7+546bGojM5eQ9HYnQsuvP7KhY1QRlxeXR1ep
YpZ8ea9GMbt9TTiSXvkQr5e9/savVWeWUlXUEPVexQsKbEG79BxuxnmUCXsa
0i7AOq8nyfd8VPSS2oJCmes7JSsfuusg710G9wfPm4XCAg9VS9AuYUTLtKoX
6x+pUhc+V4rUaVYaoYVMRnmRbfa0KUBIpPx3NK25c3G74wmndg47HqxuIfJE
JTRpH4krkAdBK5R7G1lGgrgA21/uTprUHVXVCJYIbLhsppBPDpLKhmAb+q6M
rXhtfZscF4isyEt2+t3o2t7onEk+uo/ghVauF5tQIHkgY70qxf3PJfTd2r0W
GRmLV7XXHTNoF2fcPjkVdKlTkwGDlWfuuFtfqF7+QkPqFQNhVS0oV/8xbJpR
tOPBXEYo3pqnPt6HklEjGZN5d1RmVdX+plrDsopWKX5HtvrbnZhB2LuQHb/U
s9Sm63/7QMAQN9XoVIamgRKV90yVPswflLLAX5ijnv3Q6NTMAwqYXmxe9M1/
cShMgfuBbdDdXaceCNumhw62r94/nzqmQ/w3fx1PaZpjZyJqS+IMH8z1AJ+I
WwVL96/WrYbLy9XAoTxwEVX8vFZVsyjDc3HLWiBMqVTsklGggswAq374LwCW
QZTKZB5SvB0JIHeFVFaRcufrYtBNxPvt/BeW8lyFjosoSDdwmst08Veh0Pzm
nGDBqrpGUHqaIFzlrUVZbFEcdhz2I8hLdQPtXW9/MfZFGTES2H2Iy7LWv2rm
bvcIJlyaJcAC09iI/6M4eFdotdFRzlOKNqCMNVE+tDcXldQQfQzSw7oOwLd4
F09+zrHgvaqnT+Sl5mmVhpDUkJpuEZSXSJ5MlcSjWzZB3inuEd02p6EGO2+M
C0JwJwFNVgl2zOw0PbiiqvFSMcqUtkn2cy0AhzdH7Dv++1jcTOdfbDmSLVX7
46YpQb7C0k4ISue4L9DR4tTot36p7wh0cdmyFkjkqaZGKJcU2R4hdSznT1op
OO+Yw6obl8Xs6vrtuw9NN0frO3OAjrjc8E1b1hRbJmCZ7I+6x0Snp/AmE+Si
N+aeJnGXYemh2rGiYq/HzIRcqEKwatdGljKu8/yRt/nrlFwr06Hc2LY7A4HE
5zsiWLkbqXMb3uQ0iuHUtYcvWPtVithisXhq9THIUo/a422Fx5hEQhr8kZ1m
Q3TLV5KZ7WX2W9p3+O2KYvLeWroOQKcflyuRoDpWGU4OhXXtGonkDEzdFcl2
cRYvg/3WdqsPH7wa2TuKJONmryBwPcX0+2lx825AfLfo049Btu+KJ3ilM4hA
2ntn/CVyCWjyWE9elZG6Rz4yP40fN1Ux99N8tQcdICJ2OCd8lvG2heHvj1Gf
GUItAVhXII40XdWLJgr7K1TDlxKbvOuAutHyu9QMloI4M51ZmuuxP16xDrbx
PJqs5/jFDF1TjibBTHZ8OZ0K3Ds3MRSVTHMYBzyG8/LnB4vBYW83VJltij5k
SuqIQp5FaQwiXlgoM7m26rme78wdfV4+Kq4lMxI/yfUaTyp7wqQvTZrlnMYc
/na+beftFi6odKLhdiy8QmcTBQE80s3fZuMO5p7JmW8uAp1+oDjMEguFvNPm
hhx+6l6sx8euY5p8gVYEhCScD3DNg0NpF2cYpck5LOp4t7M2wkm9QyAc7A7r
kf8nPYMjQ8g5QX/Uqttzk+dT5QQAHhhOnurEv8KeKybR4cjsN9cS6+T3njCO
w5EzwMzy9ppDbFjFir8q22h9mQZ1wjsY5MZtzxuByITTfVZoQQABZH2KzS3+
4wcuvwneDgNxaeGAjKpX3xeY+/3jiaaUj2j11Y2ztfQ+cZ+hPR2q29ggMjkU
xqSo9f38iX+pKwFFnf2nXG0Q6Ob+zWMuC9onmPCFgP5ofRubyGX0uwFgYERJ
wzVJyBtpf9AT4kR1OE2Dxx6oSKobogHzNgN/XGZm37cSomYWO11s+uFQqNfR
un0u60b44HaRheIcJl3Hd8gTZAdlxrU2ZF2zGwcAJZI4jNRhcjCVygm363Ng
7rsBtWGSlcj3JYdQfLsKrbXsxthdfNtFbIu2MiJCWPQ8tQd/fZh7WgdafCWB
f8IOeQdGvbY9a+ejGbsuVhE00/LDEBh2pn2YVdjBQLxeaFmCFByt6TQ9W0sn
qAhUr2lqdN9Y3vFUvynotHWAVUagCnpWSJkbXa6P6H4T6lYD/Er22g1x7r3T
uZ9VWHeSwHb4VOCKnwCoM53fprMipgNqtJjgY/f7EW6YtLkaloNHKI/raR0X
qTFi8w/sIQ5I6qz3QlIx4sIWH0EiQy+fN7uPW1ECLRgQLXPOc2TvSCbgVDMj
DlFVyhfTs6Q8Bv5RuqjhDdnnsSN0a448670Pyc2zGMiHqNInMngrK7cjzm39
jvyaNhmMHZg6nmnlWGF5F1DbPy9Mbha9apLtL/D16r9czxf4PAcEHSg9+VDW
4rGU2FtJl9b8rf2VJkH+52UHelapHXksDOdu4eEYG9H8xc2DQnDi/qhRH/hK
yVAJrkKm09J1YxtGEY/2NA9k/8n0+yxQe9merqyYZ6QToGIPnvb5gbFsx3BW
iQcfqc2wmkVWYAHsOFy65Xh+7KK66B8/62ydftcHUK6Ivjtli30FGMQlROVI
Q/MuR0XRTdqmF7vc+TUneWhKMzhnPk7VIJ7XQwKLxqzbPlr8REqbVp+quLAg
bLM7ijb0eux5pYOLId/Py2I4msf0RHUfYv6xH5zm3zQbMfVTSqjSyIDiVZHY
5w4HIp1StT7FRhJy2MMSb9tKNMHLGIw1LPZAA7gmBPZaEDQQW0YoE8/sr1M5
hWkTn9oAZZMGlEnZooZo5x+6rkCnP4hAvFXeI2mIJafUTe4dlg8v2tNwbmZF
lUWSmcaZ7JgfwXobdq9zYA/z8/8jVPUNd5ZRQuADSmZ0zU+ivP0ebjZ0bDkM
e9/eWbILExIf+E2fELI1IPUh3dwwQCRJE6C4QyivGq/wZAX1fmKc38KotGFd
9oLC2hzfwrGPbcXDkEhjsnJhyFN0rvKWKdPevSn7u3swFXBwlig3umVimMe/
WCM0FwVOnW2cm+Hy8bXMgNhBk1ZagcNC8plOlVjEdaIrmMscrhPBpMFi1FaS
xO+tD+hffRko0+CRhNgqSroQFGxXKNEBdEoz8vmxqenXwRHjsmVbESVsu65x
QCy76edRmsM+oakTxGZLksDBED1b6KNxk2QxZ0KhZi+YGD0158qQ0vNuS6mg
6giyIfzIJek47Hs1F2fn7jJkzj0ahG1oFoSPhz++Ffjoxv4e/1j4Z1xLqaBV
JArQfxmTD92AUC6GFBAglBUgExLGlK0u/XZVxq7nYhVz80jSx/mh454GlJhr
1Syxt+dd9uU/kKmYOxQYw4pyw729mj8gBQsVv53daQITWD1264kduXhc3c4S
sbSW+Cxuxp3dRW9FppFlWgsTNejDRgcR3GLWgZ30d3KV1KDYRv5MnFWB4Te/
3Yg5FkmGnWI6YImbezZzL66ubo4/OvoGdw59aS1t8MC3UqjpYkGQgDWYUKh8
8XdeoUhcaXn6az6fMW8ZxsuFMRj3sabic04BcE5BlKCivKfCHjDt8fchQje1
csLR4PWpTHaWgpHykn6r+hsGsbg/K6vjNv5kS7m0TGWXOAm1XWFPwKPYEOC1
ZjNXTJJfQkotxZcw+tEQBjtSitw/r7hYpWBZVsOfylm3pqqYq/GoF4h21Yx9
FDSjS6UehFJAz+0OQIZJEs1qxK7qcgv1KonQSNCkEofjofRonvC/Vl91F643
rcoCDldp6KE1kZ5UfUyzLeYkRBjMQLeMyM+HLx5cU/g3GKbBoU1jW6bq0MYL
hSRzLyFBWD745gvyccH2ZVTel4EyOMIl6f2FIDEwcay2lZXMc+udFFrUXHlb
EL63z0LkyOuOfO1woPKIM7fwUNjZU0RKEmQkHEfluPBBu7BsuE4mezkQ08gz
kIbt6EEPtK4cht8E/QV9DCzBbKWRARMfbFeF9I+UnOhCLbpUXTYH9AQHvA06
IIHkqyfWqrtJ/aNpFcdt7D7Ut9bgn34m8XlBqjT5rJAkBKZBzr4NtckNwqgC
h6X7OD1URTESbkVS+0XPkiVZvH+mtE9v0NiJkUqiVCi8GG1tO/KbEC2pJkTd
ElGA18q2w3UNyZtVLAyDjbhayFE7WkaTENE2IKBvihwEOWneII8/UKuih2hf
TIcfx3hxNhrKhpvb6wKMGwaK8YiwC4bsPQI2Wbu+s4+vgAyn1lhQKu41Mrh/
8FdIsZ8D5sjNjcHcqMfD34wGUw9iVQSCqqa2dbU1vxxgxUDH9IsgVSu9fpCl
VftUAKQuOQc2rJiZ9gmLDmz6RHa42ATvISCkXqVucqXLBeVtzSg8B0+pLHmE
MP9lZpdpiD7gYIlcGVVUMeU/2yE3GDsqHhHQ9+tqs71HDA4FD0CzRIRgcJL5
Lqf2CnZqzOcUw2tBDtqFujefQCfL2QaI1q8ablvilKawXkoSHbJ7sIUjbx20
oSv6M6Svz3ldvZ/48qRldUbj/RdPTdZ7F7n9C532nbr8nB8i+d+OkwOJrmLf
WMWLy0g+wU9ClRdrwOZat/THYEsGq36BK0VCBJxGMMrc09c0fl6huXCF2w4W
Sfx6e2RgpNYKdHaashd/ebOO0DMhj5a7sCLoly27MEt9ps35CNb66oqE5MHd
AjOI3q8S/CM93Xq5tdPdU9BHuMRvWb5rmn+oXojg0rokoJk1ibcuqUE45ZD0
2h2QnN04KN9XbIrueq8VqBevKX9pRB1ZeJDRiXAXgNa2yihTXHXIVSUNZX1L
Nayv9pYS1j0SWP5ExEQ9Tnpi1USYtJJt8fXesDNIIpvJm3Z8bGQiAjWggnyc
hX8z6m5CONoYnbyYKJj5NMplhM5MtFANPjqRQ2rFAWs+2gB9EWpT7chQ+JnP
+D84g5nVEzx4KG4nnbDjZs//IPAf0obLs/yQPwiUAhdlR0CSB73/BQ7sRNOS
SbBDLO544FFtMZ5FCdBBP2muvFTC9LQBFN1gTZmNgvJleEqE8axDg9EFuOGh
LntpDcc42z1dCs1gvcY8UYVhgYdjdHauTT/1MKdS3boHEzvxL9FhgzSMEH89
RL+MJzsdfPy8a3552G3hMmlCsv4UiveLNVjywxlDh3hcH9e9i1joWK/tqy5h
Ekwj2fEQGC0GFO7O51MNXefvpM6AhyWofLhCQAQI7CW75kU9c0g9Uzsn0sed
1PmoQObvNQk4ObVkQb4m44eheUgYco2K9yUwRpgyAJzTHZbN2V23ZnRsQfXG
Y8rqL+6oRUK92KSf5E35JZXuLLpGTLku8WXCk8oK3xeuB3zo1iMhQlCrjgP3
JkQkS6+q8J7KZQ1XfxOFJg3B+phaLMbB+NHfwxoCnUnZANzBnBek1YD90Mte
mxwS1ZWdr1UBvIpsZFAfuZz29moOaRgO3w1xTarCuXlqDy7M0wajHF2C2jqP
fTvMIRrSVaUWYb29B3quoyI0q3Lew01dpiNOvdllEKQMXQvloBLWg6fauy3X
KqAxu7qF89tVqdDIKLV1oRj5I7LfMmgWKmIfRKtrUMbMswQiPBWQjqLZO04M
YcN5hlxzGlmfRrwx5eTDycXMYK5jljKHxDpiYcHu14zMjEpZP9UBas5Hwn6R
KgU+DDQMjnTHN8QXnyD/h/ZXbrBB5ld+Nss9xvPBYnO1gzeTp/gnkAlXLBdg
913/V1gW8x/R5wlNo+/bqEv+XJYfCrqXNYw3PJrjR9Yq516NDTrWIwVBeBLL
VLz07g/iUETDNWsdef3RRKxezqv9i2Nhs8aJQu5kV0+e5tf5tAAPkl96c9GT
qRlq3oKX5f+bZoRzEWfSzVB2cACIuT6ETEvCR7AuhwglcOXsOhy8ojrT+O9u
m/bua8QXRMf7vxhRFkKNHRPif8hGKUfoVU0JM7pAAJRRiYFhmwhcjgvNhMOV
MpuYrYzx/OheevCt7zMEC0bR6/HCwG3NYt4VopftvSF46en7FKc+mLvSl9OC
9h8CdK9r+uhVHxiLnaCOZbQE96eWRoWYn4gHb7ibd7VXB7lJZX3bCOoQK6h1
PPd0wco/dMW/pdlqVXKOJlyfpCKwshNlqP0hfW1wNp0QtuziGjwJiiumclqh
epR5wHSrMa1dAbCHk0/DnmNv0sAvQnxQc+oaXdLkyebyEGOQKLKiI7KL6lN0
es3B3+lSwgnCazZbiBmGzGE3uIq9Y8qArZbow6qoS+ZPSRgS+vJA8SQ3dHOE
7dSC9FUkLY5+JmI5ZBlSOxQbEFEH7hFoxlN1OiVxC0JU0xGTmXFkGe1fnO9X
LdT4DUvFcLqV/jVlJ2c2i31Y7w8t5uAIBo45s5Mp1Iyw1AAWO4AARapJmXpW
deUpB1EymbsM+Cv7QI/Y+cKQ7cplVlIAY3xw01Evs/QYJOj2c5FvUTD3auU/
3PS15Lu+/FQharPj/76Ok1WaM6lChJxX/l330i9kxTroNBe1aVGoFtYUZSNV
L4Ets0XwDcdAWAsvk4JzLU/JJS5ifokXpBoga84X5RrkWofEIAD+VDSxVCux
aDN+Pcl1t9fZ6wGblY9rGZKA+jF/MbY/+PEE2CCpEp99pEm78lLKTC7en/ig
sk+a5M6CEtbWKf2VWkzcpTPs/GoyhUax9NZ6DQG4bNE7k7AY5v14PMffpEYq
wPdfSRCiMJS++jFGCs3Uf4SPpPFRRvbm5Vq7M2zCFbRenMY2608c1yvi5exW
Q7sNaodeFKBpTBi8gykm065cwKdslCWvAM5F6kcn0xbtoB2Ud5RRH/5deMiC
U1EiPGkspAEcI3LTHoQOiIfardsvg1GnYpfzXZKlAgxEY7drS2bpCUo8ERmM
wRVEkH+CWoIGtDkbud0qWa8ONOQ2+X3PLcR36gag1VBScBNQp/7qnRUdBERS
Zijp4kjdkuhlZ6dIzviOi0lD3QzPZOn0yRfu5pvBMdkX8FFMVMimGwcmG4uJ
8BDXHwXmMJ08g4gzUkeVVsRTyWPCBqc+WA49Dq+za1zmNJBasBOXuQdMe7N1
CqsctAOH9o/Fcqjsdfm90jPeaPBojUMs4NOQXNL/EvEkXTb1oxeQxQKwuQUB
zgGBWDf4hBVNRk3x8kNxvnIzcMp69BBGXNXI6evZXGqcrZ/Byp+F5Nbn8xwS
8qL5wScM62QGCVKECwc6OcNWb5oyWsKZjP9IGNVVwYS/KbQ6pO4I3+G6Jxei
QJPGUXb/wQFCTpCwdSwVrmK4lswsaxYLtzL5RP4b1TmNXiv8sgLEb1C+Naby
1FnslxNfcKttnkXZdk38zZLcGK/9OyAGjnTWeZYFxfqoF7RiwnfLnkHLq5VQ
pfrMXUpoFRDGyAPc9xNmZs90K4xCQIsdkBs5nINrRmqH4iFmxGaLgJsqXbsE
jrIcIP9gpLbv41Q5fnBAm5f4EFSHbxUoElPQ5DWikpM2VABaXp9qq5/V9ARH
/UxG7r0nIjHuhdbhtwCannJm7uhbtk029FBtfsXYlXNQjinvQc9dKF9Bi4Z8
greV/nZFORVn2NQL/NwPWz1B7yELQKmRySQqdwAtMDPKdn6Pfi+T4dGWIQGP
5YDDLNnhCvil2PmKgt/8p1M3JjSF6e7dZe0F4eHr+hkis9z1G3P7N1szJJ0c
OoJNvD2TxgMZ8WZz3e8Kt9rDtzIk6sZ9vIIj9OJ35t5ZnEhel/k6iRQulu30
4OvJ+hM3BOfPgMS2a05VCFA6Ml/nHCazjz2j299XbT0ditZRJAy2wAoxEZWr
ExNyJS6Jv9rMB07czUdH5oVRptzbt2o+aGS3nXW5F/6HJSB2dF8ISVIp94eo
Gjc+uOIP0CmnPMh5apaK4/pJLzeh2/mN+mrwXD9ZQMVG90WGhsH2ra1YktXH
5ZkyfmlrxtNFkplmQsa1GBJZpK+o5i6sSP+0WfaFNhdjzAx1p3PowrWzzINM
0hEmDTK7oH/yWLQ3ZucMm4pCK0YJV0DtuPLyEZABkgn8f7RGUU6JXAXt/lZY
iq4Og30tP6QoVaQx91x+yUsz48V5TH4+hbzxHN53Au3hVOpic+o33w2yx0aZ
R9941eLibxHnOswv+ZGYDnMHfZRT6iPwlAxrcdvVtn2xiB/1ALAXS5uub6x8
lI/PFA7ii+VG/K3YkPawZwi1WzYWNNPvzOi+pkZVq7u/cfv1qMr/YZheSXWi
n9eObdU978J3uHg0PTtRO+SBySQYroPWQrUSfVvZ8e8xdgoCST/hrhzxjTMd
VsRnYxubIDtMr3la9e2TvQOeUqTrjPHPAJKtgI6Rm68MXCatoBxW1ToSnjli
vQYGCfbOZysHjQw314gZqpzWzeoxCGxM3ZeV7fC5HUN9dJiVB8KaziGSTMvv
kaGvdOeklb3cas5a1ThK3t4+qfF034madqYo/yPUYzqp3ILxmWIYztcBXoGV
F4IxCbizG52V41fLtHBMtGpG62doYqtKPmQBm0xA2PU3WvJ+juJOcFmClt/j
GWcelhFs0zijh5zBmYvqLn4kFLDvBQ3ZtlQZ0aVrMGRXyU27B32y6nGZVV1G
rIFdeWrllt/yvFdZoKsF/pF9GRM6kqY3OGdHZ/5ST8AXmQ8eCYAiQ2PTntR1
aVL5xO31j23mXj/hmwLa3BYwdWCviKhNjBIw6KCgE3mRDKYPL2S9xNPK02Hg
Jb6WkfFd68ICW8Lq6oVSQqlUU8pzuGjkDU0SFiJy5AtUjz+Hqtv/Ryw5+ym8
6i7bN90yY7L4Yx72O/n4bwR7zgIbG7QFGSrusQ31UncVUSyly4m4lZFaqgeb
nxhxKGKZwBEw8AcwH0Fv/2jcnFoue/L2Xr+BEyUaFe0NVuYrrulF/dbzbg5O
NzYWNMEzQWRtGdf0ARV8UYWbEjVs35r1euSN10Xl6Ehw0/kk2ai+NE1pW5LE
/YBtUKpdulKmx2CkbWAdqsKx7APYWIKMyGJjdSyE6c3c8HqdgEEXNW+3UT1s
wr31aSOmmAbsZITZGb+mQloqVy0AVofMuY+tdsgehX0nmIAeWjAHhgjGupoK
FKYIhx0VQOWYGXiJ6CM1oQihZW4xatgeWG5OdykAOxbI/H5wvXQZNX3+XzOd
dPVNSJx1dNghd8Ah6ffbKrZPUyvhLgDT6fAhqkUGXFKdKJRC2/tLGij1oBUp
D9HBjzLN9YwiD6X/mpAN1sUe4wNSZKrbJoLDdPPOSv3eyg+M8EPo4Rbz1ATY
lUU4wo6bLji9KeGJxh+NwD50taWxn7/6K19u5SNgRJhMbdi40N8UKw9r2m1U
m40pBMeo3uCVaGbK93/mngy6bgML00fsT8p1XRcHwUAR5s0jHmHwdryJLprr
YYRtEYmIycTMcQEVJPAgG5Cu00XyYahAiPk8tbwiiCkCvgVMTJEIZecg5NmK
DyuU9MClyz6/Xa2JyaJsyivU7WqgvxjrybBlMsuoCbH3rS40bxF3MMvrsKsD
QRqcBtRXctD9B3/dVCrS5x/uUmya/4iroeU1D0OL5VN5y3LJ/Y8hnRpFom/M
okhBiqg72OjAJTUS7Nx9qhq1VOdFyW5zcUR3omFx2gW7Fr/qJUJ0AsBefg1U
udP1sKYUSTzx/AQsxkB2GgxvhIVqSNXiMEcaQHPb4O54K+8WMyBCRPtFsFxv
efhBPmfIwjosBXhSDpYw5kICfiF+tAxn0Ej3Ia1ScOaD0AFml7sWPx0VWwp+
S/AylKNB/vWHycd1cZJ85AhndMvdqzBCETwJxZ5XjyhIZumIwr25be9WoUDP
T6TJTR7bxtOf9fzL9kgW9XCoR9HjcB/lpwjca+21RnH1p1FQKyhNqjSFRNzV
AvqZ22mmaCy9mumvzw88/jso/tZAWCFW/F0eP7QhPKduZfbzX4WDJHKEMGD9
xzgtpNvEXZ7MVcZRG2nCfFoR5ldi6+qVL9DvE1UM5PUSpfLKE5mBtwyj33EE
CphUywmZsuVIZGrsS8koxvLBHBFfcf+/t1ui06F9fi0sQ0M13yH80/fx/40Y
j5OBYHQLVdQtfb8DvgN+e7BxFQyVh1u/ttuZCE/N7LUh7secXGeg8FTROTY1
PK0iwqHj43a72Q4zukBkOwx3RWIY4Di4Z+MZKqprcZ1OJrf8kh9ILig64rTI
i4TCQAtHET6KXGnpvUnA82GGjS7MqRu7s4Zn+Sx6WrcMFyzNI4tbTO4nJ15k
MWGSelWofN7MRcdagofiwEI2Berbi5ezfqi+r9qpb0xSa7Wv1cnCajgQeJVb
CBnT0PEgZ7IzbBvO+S7HFnR6PGb2EXrJ9FnVbcf+i4whhh14ph2fA4B0BB/p
M/3RuUnPwSftnxrbHWZ2mQofborljEgWYVzsziIT0zERVzz8bc2wBS8SFRg+
qpDZRI9WuAL6R6XcoPqgWuDRJ5hoayKp7LLal++R0nHwMFqGDde2Kwj+70sf
krn/xiRlhZPS+WpVLiqV3P7/g3M4vHVhLeST/SOrc5s8x1h02ShyNCVWnczH
az5osK0lkcQttREPFj3Dz0e8pK5nzzNFLekYvqOzJ2su6At/O3du9zPZiInl
4aQaJM+9z6dOtz9Tn3sQxG6PjiEoWaJE74t1RQT3lypqXWzm6qHWd9yI2RRH
cT2577kzoNXXpk8NWKYATxR+oK717q2Qdeku0l28npf3Trfrorn4v+Mm5Bzs
5Xbz45SnzZ3W7I5Nhn7X3gKEqvxTc+tz0HfImTNdOoeVScofJ8NAba1UAmBu
vrHftuG31hzyiQ9/oJaVUe9y7Km9IoE08tj8B+Nz6VneC4UifbpAmLZ+Kuvf
vF0sc91dfEu9wSba83dknErx+mmWMp/NCfVRP29DDX8LYjDtyMdS4oM7M9wr
QDFoS9T9FhmVJtwo55bzCXExC0lzNvjslkA3E9G8PeB20KruzTiGHmYLudqP
fraf2V6P+D8R63G+HZ+hqyln5oWI5O2rny+oqPsxsytwC3MCFoqgb2uOm8Ag
Vzf+2D5KMP9oiGtbZlCTyNTXvf+J7M6IbLTBpwSC9zW6JI/uSX0CLFj+EDa7
uSi6HOcX0PZGPZAE59JiXt9ddmBQ11jL4CKRJbIU20TyPkPC2akW8lcBAFkj
xl2N+HJOAtU3IdlXLxw8UmR4dq0fBbRvRMk9RFuWuZAI0Z5PeCeWSu2hdTRx
YU1Y7K0+tcg/EzdqnpJKTiMLelm0zzTDepBsF9+iZoNB/QgQQ+bnAWLeZY0z
baMUqOp2KArnUUIBjVEVRqFwFL/E0tlfRunCfHA1M2fwap2QeImj23vCuSjq
SaEgYB3Q1cgEASpbTAWvAHeMfdOLvFKzlekJFGvNExU/zStLyvtFLguorXoT
Lu5YZRU+cBJdRu636gdURRM7e2OIOI5cYRyH49Or13sUQyiAR4pyoQoNqHAA
ggUaCjPvjLQjp4i0hbZKYj5xyenHlUOuIhXf8xAuglfQCkDXZ46Fpyeu6Y+c
f+doSEr3cKn+EXnultue/wzzoqFSkG3AhyP27B5kCAa895oo0uUYubnII3Hg
owvBNOQzIFcZMkflfHHqWuKrNiy2KFV7gQi9+o+siLWCmHGLyW3IQFrhKg1u
eyMYTEHi5BEIUVaZPFpJhgfoW+tIYQL+plKdJN8OqqAAnadd/h/NJg72QMDm
1caG2mJvG7g/fsntZg3mziLF7DOwUnIPEg0XmUXOsSTFGQcF8ARxVRELxmY9
zUZduKu1jnODDLaqmb09PqOLrEe6W8Zt8Pgres+5Ufs6dVJaCCzcMsuO7XMy
RuRcK8RMHpXw3YFuEh68CyTe3N50d6P9BCxnzXK4qs3ddXqv7H7+EGvEZ5Sz
aZwtZaQ7IYEgwLgFZ6hRTcmlQiemABFKZ+1n5wBnoKlDUYa+5+C/XvXs2kFV
shUuhg5hKPEhzDPMDThS/D6vhXPw7MIcwRj9+e4vEF4/RV2nEHK0bGcdGKy4
Vw9U2AKxZp3mVwZ9s+sOagzseQ/0vdFUimPwC3Jo1xeJU9SxxVseemf4UI6B
mFeYW2HMdu0xNcVAhgN/Vf+ovWk/7saeBKHejGM/T5xVxU69igwa6KryEaA6
l6rg0l+WzuOfFjTNPEnGRq8oNPLV3IkV/F9518WVwbi/s1qwvLJN9JsYngLM
2wT6i8XTNiINW53s5ewmPG8Ai+4B9vaojR1fPJOqpeWvk9u4Q7igX2yrql+x
iHJC0nyzWC3Dgnhf8+uF6MNX93M8U5ioJ6AV9alDztYKo0Xq+InfD4FypoFU
a1XYLMpPoJs5WAd5EDlp1HoBld8K8B1rID7Huya6Wv+SWIfYKQTDmTwxSfSj
sN68k5WY1bGRi82dwoVXttDaT0fA6wWiYeDzLBpToA1NzJ3Yy2k2hQzVNRx7
wc9AMRPYpEC5zH+kDaqzITD3gN88ZLBth8ODneqifWssLKRP/Akwe/iUPets
DfC4QRISfFCbMyBDYOKoemkZ4o/05sXH+mGDBZh7LJbGdIzjtphV1GM8rQti
+Rx5qWjHju4+eUcSsI6a/8P7Zrlew5duRo7pk2OQ1IZjpCM1Qit7O87DjspX
AeFBLI0ZhTPlumEmvkU9xHt2Aofu30ocNuQx9QC2Bfci6/2vZhIa5VYpUFnC
gGuuY06Lg1bOdFZdJsV8KYP6jNGIJchyJtkr3HoH9WqgDkD+5dOerRgkm2q1
aGV4GPVOHjvDCLW0azMpqN7Zuwl8ekhSlEZTUuUyPLCn8uEVIQdHfRp5WQgF
EhZ9wjCC0nWo27YO9tgW2msO0DHByfqcPqAPCRLUC/4NKiA1/WTBtK2kFld0
cuapKTfOBsoAO7et5XeNo22TrEs9uaeVMWYP6/3IkjP5IFKs5ENWDC2fW0dT
6wo/PMUtgyjQatnSMyZ729xW/ZHWbuZbFZyXw4vqn8MMyKGpIVa4ru2Fvu1T
234B/nYOxDpTt2PMIjldq/Tk7QOM3D+2b2pWlfsbFct5IWMPgC3sHMx5NJhc
suteG3JFpcJuUxkUEqMtxXUPo10nyE5CXx9Q1Uu5qYHnAnwrgqqDtsRWi8s0
n2VmjJPufZQC24k6KsujvK7WPLkPrgosctMPm7/nqN+aKAQSLIbVIqjvSUJr
p06sGKtAT5OPsXwtARRfT2udZcDk3aKf5h3/7wzadKz5dDxa+xH8W1kLyhrE
usAqbuFp/AHGpqe0qLyi6uP4f8CzNaqkiDHYRgw/VNln5DhB0DWP3P8vsmqg
xH7ieFU3NUO3w7IB43T+2+wwDJTgWjJJDIzi7IhxJyK251KTaRREJXX2hhDs
SVKWHL+53Qy7zCxj9hQIchDsz40/2j4RXyoQguqzGMVG9EwiF3W1KNqKxhOc
O8gNt2FX/+yYLbeXtewh08PD+C/tTu4ZXzeZAIRkbsZcyjIOxL0dabWN/HPz
VUrfXNBvWULpddNXpihsjrKL2VfFWpQjjupNOikrVl/S+scrBdvVONlpEbbP
Ram5dr69obkzYJsAZQPX1iHUNuWvLMJkNmI0lchak2OaHlhCDrdYxo2vpjgi
0RITXpryP1Qg9upQJdbzafmX6g7c3gkVFarwaMwOAJafRJAUWXdW4l50RnPe
1gQ84IEGWxB5Q1+vzHbrrVzu/adwzqsUr8DSJ4XSIzWgQLHozAFAsbbxL4Tc
aPuX81KcnnJBbPijr9KhYB4Vi531nv0R0T6DVjzvJcxhM4pW6oUdCz9PTKaF
8gPvaAePlaQlcV9VddNx87PDq5kXptCOg0TDwn2AuRM3kgTYSSFEnZmfws0t
gNYtotCiI8GnqOx4COa5shgbJi0XrNMDAdWdYmNCuGoX7ra85qo/1Z3E4K6p
KgdwOm8Zj+SsfTZpUBwgNne9IRw3AWkxYYCU6Zuds63k0J86i+Ipr8nqY+at
grCNiTYGSh+WKwwTYjPGomPxzDU0nUdEmjy1uAGYsqqCU8MrkbFzRFM8rxyN
x55AhHT6Gw9minbGvRm3sktNIbhzSgMTb3G0DrT3gQNBflBnoZQPl8kULRcT
/VXdxv6CVk+SqbYKed3+5GJreXHq7AOt4JaOZOzoSOfcEt0CqeaHABGc7aSI
RGj924a+Rc7lnndywlBMkaLIOm0YsCHIhk6lzoh3/aVT4n4EWAgKOzUEi14e
/aUmx3bv7Fnyk5qnaP+8R5Eqim6DrWdGPvo2VpwlMIX71atrsh9oMhJqDfzC
y3Yft4GcC6+HshhoD4f7KnUzA/TaaqyOXQZf7lz8FRN82ROxPATUTyugL9Nl
3BGfr9DwuPSGPCcEYufaLproumPx/WoGMBKZ11RsIPMQmyVxH1tTwGp1B7lX
gVcGzT9dJYifsO/g/ESFulGiooHyyIA3eaw/HdQ4q5zjn3i9/s+WUlOUUA2t
xM2qGqLrIVAtdz9bR1tH8b+Ei2wz4vgDmHY1222M3lPsLGJfUbm+MU9Ha2GD
HtPAUs6PBq4zAypsV1G5WR5EwrrCOQ8eYxm8MFhhWHdov0TpmWepeEm49o5v
sDP0vWjOqvKcXCvbmFCxHbZT16C0Gnc/GV79cbENhI+3DxKMdNOeKNx+7wkj
FcOIZfP0HYOHkeL+huCOSS8glxpSA1ilQLKrW5l+M+8IrHOoO85nfS6FNrwf
OUlPA34+Ro6c5JYVca6vFX1jeFXEczKKe9AqipA9s++XG0n+y1dFuu2wuwiS
U2O1w/x2Yxs1JWCacj5ImSHM1vHaQxg090XvZ2V6FlfpuFtFQURFyqe5uJGM
nwkj9im0f6JuEmlnWFIh2pll8auBz4o+1koLDAnkDRha1qFNzYq0M8YrXX90
AGfWuYIEqDgN6swPP6NfyLTaaivHg4TzduwpKAfgO4c+DpgrPUVn1VJ01UUf
Ba9NwkxYqamSqF6iBladkqIUCmJCaUChDlq5xybxWDlx27IXrsbBMbY4/4ob
JQeSSesiycUZUFv2g+IO3pyPqX3BJMMz0XaBcvOycc3U7hB+0ABeUQPciYoU
ZoNUZaxrfU8b8Q6sZo6+B5dm5512BIgchD5paX1yhDkgCFcmOA1Dw0FJBLiF
Ti0/a383o2lM9Pkc52t6vH6za4hSKtqTcYcKlLXfM3eS6jsgvS93E3NbIV0E
GYTVmNP4aCPzP3mgtpet0VRTmiBpT5PLEeP4AAN6IBlC+v5X24qRDZC39kuQ
0WfNcEYqU37mio/m0ZvIUEBhoTwJm7JHDmzoA3sP99xpYll2yw1+bT4wuB1G
tdOYpYzaem60uEKL+G+0FeQ0AQMmwk/ZCU8o2e6/dZfa1yAwT/qXZ7r5b2Rd
iHRccw5gY3OrJLGCP65LnbDF7MyH6zatZBmZO5/EpQM0cnXhzCgXTs80z4uM
q7ZON2laYgNPKMDJzNPvFeP2jYd4db7xiQgwMhQ7h8he4me7LUz4DnkKvpHo
1YJ9g66ggIU7Dwx99KnkNhkKRrQiHHpWB84HqxhGSWpHsEG+VFCCJ/71lDoK
uuWYg0e0IWDyNPJ8j7aacEQRx2syuLA89CUQjkiw8dB2fAY8DeAc3o17sD4I
z6nvzwtEXMBwh43YmbTICimOKqxROw/KolkCTb7XoB0ESM9hm8QxlTEQTJLP
hW8udQQeI76TIHRlAx0Hz1aXzBQu8s3C6l16suXp2sYFpZSoxscJNuV/pfml
fiIjW4f4u9XkC+Z4l63dWP9+zAai5Q+uxnx1SNM/E08iuuVJ+nEt3FeDja50
LCUQi33utFOx/KMNoJL5cYDimm6UcG8/+YmxCF9CC+W+16pRn5rzCHKyzw1t
FV8QN0w8sBQA43A/8FaYmdoJmFPPBKAQA9T0mFT2Lg0vNYPV3zZ2nETYIwae
I2L4F/S4mt8PswCzYZzSqywbzIRMMg2WTGVdYKX5d62cxG8H++i//fE/654G
TKwUH1AY4puWdfjSQBWIY86v5cO6E9Aw+x+rqkugL7t9QEKuHa1N5yGsbemz
752oXYLCCSv6KHUPlkBO4s9TESkunlwgKYMyxSVGt+MBHF1l8PDMtndrI6iq
2KjDjw7tniksmsBirq6tMFTozKqKeYlg6NzpEWFLbL8Loj1y1thm0XQSDkpR
q5bLwMQPlX1ot9JQoUaFBgoi0rYs0StdvF0yQPtSHfJKKPD3UfSd0sh1oMpU
ylmcK5qvTZ7QG3SCePcqaKVqYVmTIWXWxweS0MeK2f2orHCjEUcqrXnqKeXV
CplZyDYFQu2crLuiU/MS1+Ax5oth96y0svwvzLwm55d4xUmCUur/XKqRdpwE
c8SFxvGLIOtx2kLrwwp4ZwDwUmJpfjX041MHvTmYdjXDTe+JHJsGNO0iBtrT
cG0FgVdgHmhby0hiQacCTD/odcfwVZaf/n76dxNstsIXzDmLM4gGUEwVxdbM
fREPj6RZ4APaIpF0DXQsenP3bh2kpzcZ3SoQT/VE3/KMr+Vvfp19WEac2lPB
IofHXCEgoUKjWjQvkvNiBBPRVP52/rfYVIMg46kwVNkUBU3FM2UDQjNiLZq6
kktlWEzwmg4es0Fgl8IbRMCPprmaxTOhEBpqQNr/WFsUomYS8Y9jvx2sVTKq
I4pWm9AVuMB0zKOUtTtWBVgkjS8OO2YWGC0R1u7fRwcxcZpp35oBLs5rm69M
CT2lwHs9b0kOd/W3TRhPz+IUZSy8+TI11ELr/0xiAEbrhuGPpC/wIffXsvns
Dzb/Z7xQo5smNr+mdIjxbQlcCs/C8i6X4ulXMtKcyl/XUnNYUpRtpvuQGI39
NgS3EwLJufGMaPc7Zo4X2bAGNm+83ZB3FVd00HIBcaZcIcxlUWa3Nu7mlv/R
wC40ph85NQmT7ELfb9sUEx5ohcdDfbLIrTCv/M1ZDKLsmxK+dHFApZHsVz06
Ug3F0s8Rld4QkCp5DsD9rGGZnWPtuKq79aZldbfBTfRvve+OUszrkxnh4Otp
JvHhG+LIrzk3CH53SpSnpZp75//xacu37oN8RL7K3IZtEOvbK8OXjvHJLsCl
8JBxAeI8/EZ9dp57nyFRbFMy2saa983YShZBp3/2ymWP0rI7YUVaH3iKWAQv
iMS1CkvYTekgfRaL3Jxn1/IHW/FVle4KJ+OulE6naFz2CRhlRKZBvY+T6HEF
aKw9V/VZ/9hV2rxsOziLHfAynGF5H/J6IECd3cQYGrRgO9rdKulQMIo3fATS
pxq6JG/isI5S3r3RBrnbfaJCNauTFncy1d3Bluj8/olKcxlLZwZmTJt3YT4D
10aByqai4CR7qnnl9fg2z7sw2sMj0j8HwnA38oDbIvhpJCI/yQBb4D1wVBla
mU+p2JdPG8nBW0rt7MwQ9zyiIwDagopwKQW/NTXr9EJjjRAshk7UaQaCyeTs
LfYluZJ7PcfyYs1izHZAcYgCgSvYu+TQe/khxK557rdIAlEel7qfrsmeMDSI
R5fQICKNKPEX/lnk8s1zS3mYaB06XtJun5o3PYVbt2QZiDbwGEc/LLbeZEN5
3d3x/jnLEpE76WHarUqbnPnASlEgfFdweSmrM5ot+gSJnM+shm4b5IqQJp+8
r2JQPdtchZ7MnPOm78/vTAJDKcS4f3ZbExLOVflq/gM28QYYRtZ3LbYUc1uP
FosmV0AUk/XFcchDujLj4ZP3ORaV1c6H5R4K4XsN9GSGc9R9oZzef1LCPvQG
n4RiVHT5WW8XCESKF6dDcAHS1XhuX55JCPUq8iTm2/phf5KnE7uOaW9C7GuI
BjRBCc/8qVSM8WQdDFod1GBlIrhClZbooBEwsIgDxUfS1/xBgHcsSio20SaF
HykRG1HWmYILVw+hnqIWBSuHQCxIxMTzSeRcPjgJfWcNF70a9m0ecYccQ7LG
/6Ge2Ug/UjWPFi4b7jUo7LVJkEObn80SsdSW7LnZ+fCToWhgu4CI4xyd09Mo
DAhi1GH/6qw45MKmdp8M4O2G2efHQW1EV6BWmlPGNAiWvCv3E07agXX5pW4s
CbaoQ9NmUObT4ETbaA8OLpxrI4146VcKl0WvmMem5PxfIRPwuxvkGst626Kx
m3Az9lgYwBXI8vNagv8XPvqZmNZXjKyh6FWxEAFjObzbN9iCvbAS0iNyyqAJ
n4TZ5aL5QNx1A2FV1FznIT0KFlHR82ePqZDGJAN+MV1AmA5VLgyyBh++VO+k
46Fw2TEGvHfNznOTv+7hZFS4BJpRLtujdfPOQ89ksUzpLrn17fsJP0eeyDEN
b24SM/1WgSYouHhkoGDWt93rh/QivLlbqYI0qITSnHE124jbasqCUBuwXpEb
Tbi8aEQiig0VA/xnAqXemNBvW3rou3n0mKt5CQgIccSPbxkmvF3D8taMMN/4
Pa51KRG9MYeZHWiVVB4CDr8l2+QyVftNy7LrMM1zk+DYmpmdeI+Jp8RIgPuj
VFAc6YfSQw+tP8j/MOtvVNVRs+mmM2OJsmaK6KSOBo9vaamhrEf8mvLlVTV1
2RKfoh4dGZF6BqhbJroTtqNdUKuCRQ/KRoP7yEosNZS2iJ+eluWAZixvBiJc
XNvjpHHNeHIlF0nEq5KKoeR9O2Aqgl4cllwZyVAiWyKTSutXxP+pulsLw4gr
+iePEL22ppOJCitrSyZ5Wj7OWzDDHAvyqU4zTElDWQnsY8JO7rFguFP03LhO
4tCYin6jWU9yo5swVUFH1WPm0qepDXFlukpKtXM7aZd4vDHK47BoB1P+x0bn
TXgXt08POGkZgnlFHPUCTwI/mwBZBazk7RHVEQ78AtWNEgmgsdYGfBZKPsH9
K4yTc8tyREJpIK0WYt8op89RxbHdi9xDytXfmRS8jwI6fyDhbb0t+cCCkMgh
/3KW+as6x0phCRtE9lMT2rT1ALJgwI6lbhd2R0KdALnwo5HBXiSJm9DcuoT4
Yw/hLIOSkOMC2gr+N8ydSrzSWaQy/Aa8EULmilbtGKRfDQeJyPlCwBElqqL8
4bVCAKN2v/I7agdX/c6c6oKJayOsyE+7PJTPEiPHiq7og+044d66SlppnUPS
nUJbzljx+/rx16IuinDEG7zC9IdZCm8Sh2S1/y+YKUPy2vnSG3+NOxjM7Vf5
GCFhkX5q0jfWBniem3VG/2GZrkSNvtdTchXfuOlUbAL2+aOwbLQBCmrZcrCQ
CqqsLM+F1rnzw8VfIKivLELGnUJXta/LEAFkPmYYSX/LAxIQgr05jZzSeckb
7J6I2jPODc8wnQstRLPsYJrQTTHJuy9l3P+gQlJ6xhQwjFeVahV9tJxMDn61
XDipJ76dQtm6rNS1dzswMHOJx6gtdSeCbQ8MZHp7y4oF7x8SBcbQfWldAlfS
9bhqDKncdvCfxoPl441fso6RZ8IuBa5MrtsXg8JS+WGm/KFtd1Rj/dA3cP/W
kwpID+HtFqwOTVNeCBlmvgpeWNT5l62TtYXXZ/HZUHsoOmmMUhxbB6NjTcWa
XCH6VI83L+I8t9m9GiBNSu7esHpcAiRgwbmyP7mmHj8tgOUvPljxa8Mmr7+4
SQ37lMDPLdJP4A8NhTWSR8BDfESLNhy4XF3hjB2xH0lK4TnXrCfWGoM+54Gv
2oY9ptYLWucH3INziuMNK8UyDfFWrVH96qA7ziLjGqXIPHbcOK1ManrbeAuv
M8DKeD45sLuHxQw8zFz2zIyE4M8TYqCTikiONLyMWzt3qb1hCjI9/3QosS2n
yOdfHDKgyvIlnuyp1B+Bn/wmy1ZH2BmHCFeOvRCrlkH70AxZu0g+yfxPV1ay
MSd0Rv/0L99kpEpUSCjPdpOp8E5oThoEs9vADgM2HJIfUwDdLXQ+DmfEW577
MK15C265tRFGDCUnRVBx44ih1BijaIF1hIL0aCNI/1PuDnXxVMs8U3uLD8Pk
GLySmniDaLCNyOZoEXAjGJnPHs8Gwh2BSBAMp8jGt+qfTKr+oYtJixxAQnHe
M/fIRlarKV0vW+osm+Pu+CoiOPToAzcVtS7gMIKpG+9w36v/JL1AZ6uTbbIp
rt/pSEq9wR5VkPTNctgO3sHy89BSv3Qy29kKf7qNsQNZ0jKm7nwP44cR9v4c
CSrwLlvZ7F57TrPGZN6Yv0GEbrg+0XKc0SJQynW8RSw2waxUyhJPUhYQ36nX
CTJ5SDH8/hqe+3O+Jf8ozDOJDebFgzpc2mFzHFwwBsQ/BvtP7Y65F/Fp8gsC
dA2+LYZ2X1h/AtKxLoo6vrdV4FfrnnqxNe3lZLqrlDPDbA7HTXrisdo5dZh9
nxFWizUV07/8WDoG/YQmcGytrzUXWMya6j3tcdkeoXUEsTYZjZbqKlzsdC1z
RmkgHP60hvCmxx52gqdouyThjQxWRhjpeN7/XwRMrSYb/CbIdBT+vzhhQJ3b
QuYb6NfmohfiQzVdt2HuQJ/BKrPyRpetJUbOkTd0cFFP/KnET+vmNOslToFl
3H3EKl8dQnFx51ILMYvSULnL/C6HxYvXbkSz/UETE6hnZLlk6mrRAyYlqRYU
3JOZKsVEjpkyUitwx+LloOa3HZsu4qbx1tX5L+V/E6bQU3mdWL+5uBGv0Cd2
mOlPOUtIt63MduSe4SNg4ZAXHysQjmD/iABRiqEpa8RqV+ETIBetSXiaf7A8
bL/RvmAJdkfSLioN3yu6mQC1MsQlydevDIFZZkm/EBPenabYti8VmlLPRdbU
xRfsh6SvYX7mls964diBcZNlSjNTZ+ZSRU1cgnqyl48ck+zhSfKv7RsFHwUM
ScNwlygfJSmpMbOxh8BzY1AJOqR3gnmQzgi/65AJe1i5+12m4gnyKZiB0hBA
33oX/7RHovd+7ZsVKt8xaS4Q+SHkfUcYh8XrWmF0HWsFdEnKc5TR+nVamaXD
XstnoAkcENj2+XDnYCoua++PQTWxDQ1HboCSurNMvedHnTlznzPfJOlWSfAq
IdS06sT/x3+7TEftho7HlBvajvlZbtSsMi7a28ojfn+QZhVFdER/GWIKqEx5
2wDj9VmHd7voFkUd4PCcU0tnN9Lfv9qUy0RIgr7puelRSQgg/DfEBcV5orP1
wN1Xqt++Fsl5BChupfol6vPArXuCTel6KiQudRZbH0W5WYAcQ8YlPvzuPeY1
DnpfWZN1OtxjL2kTtDAAjRUg+lSkUYiBmxFvuMeZcueLlzgaEU5azKrPC0Gz
1LO8JhADuRZnMBUQLUTQONM88D1wY/rOwemZgwCryrvIFRMeWHVt7udrKQmT
1j7ZcHGU8uy4em4qzJgoVOtXJQ1DzkiVbc/INSJmsehsBrmhscaOfIxF3bDq
4KrTffeoslavjXoqcM1PcQRNxPqAVkkkFTh36xrOD/SEkVjh1c15EkfCf2ih
D5X1175je1yy7OeqhFKbuOC4kACmnIzD4BN8Aqe0lTFZVvGvPQZ7K1cOs9Cs
+1TIXU9JM+px2v3qc+bUWAp5Oy6nczykzdpFhrlQ6UCUTX51mhXbwbWq/HXp
WreQDZqXg6yEs/Fen/RLy+vb01ndhT9K0Dv9aqQQZqeraDb+yA5flRz00z7j
SgctOSAFLnOJMiB1t8h36uIaWV8QuE6sqjRAdz7sbil9QHYkXQs4i/riVfA/
iK0ZnreEgamUTVxMiyQtyLwvzFdEU/A6cBmvGr6wOuJ+pcztjNHRq8pW1+nf
d/6t96IG7uE3xjpF6yE2a+kgdY0XhhljHZzNHgOpEdsq3b1CEl2IrNWZ0ZAR
x6hWwDKc5tTLAu8p8wMpDuaY22Unh3pEttMCdHbhuf72dX2b5kiQiKZuQHSK
BOjr7iUCwbwe5FaAAM7hjNgfKUEl4P1mrUxoV9Cg9PnBLXyrbhD5drhRzw4H
JdYtGu1JfvID2SuORjdoX+I6nT9Ti7GEv+rQdG9SnGIYl/GKCu0JdfuBoOvm
d2BWOR7yk0hqdsnzbGnS61+chzqdsVFaD0cNE2g0po4yfwOXVAvDoTq3ZKY2
DmYKyy68br342PV095MfNAADTT/MLHoXRi1FqxIYtohYXFYA5oGxpx15cthn
F0xgD2DTGrbcMxfdb93qrDMNHpFuB4K9RM6Y9MBTiF3wg/XSNhwPsqUI6zB0
eKajW5K/I6AQhp5h877OeijhM6cHWFVSDfLOdMdnturXp7dPj8omRhby7XQJ
WrGUih2ynz26Cy/9Z/fhSuDp1MDpkC7GtNGJZgY730D5sxluHOSyt+fOTBGq
HcpeX8Unbm/lGeraTLvRC6Y0aygehLf+8ZKLNJ32GFU7oaNP/iuT105+dCPt
ExGOy9aAC2V0DBWu5/R4+u4n0me9P3Hsqa6iu/XYKcGWLW4S/m+S+RZFA0RP
f2HrZ1dvV6AOJYItB+r9O7E5P0XX7kPYaGaLtUCU38lrgWvwjRvpFCFZPLKQ
W3gUByFCxWOsZgrQK3XHujGy8QfmiWRz7XjXX10bcEPhTyibRgi3O9nlraeR
lt9GDblisEZwh1Y9GQIDnM9ZwLi3//pKfqnbXC9TRc2muY3xszTrvV9jXLMB
sXqj2hxWK+jEYHu7pXBJ84AAaddf2BR3pFdisb3Bk9Vt2xQOGsw5wgXy3NIz
oj9dsTcv4Yd34rAM2/ibkSylHKS3YvSviobEg2mHxpYvXGRYUh5o2sUpXU/K
0AyH/T3Szk+L6EAtGcXol+12IdDidjK8GhuvjmHm84flmjvll7u99Rb/ekoD
2Uq3URj5FyYDGXQ8aEqqTzEL7a4BbwX0sq5CbjnhOiQXmYea0JWQeZOo301m
Qmhfmy+Cbpug/3aA/wsvcuMfydJgOpXbKRiMvlGBvMvHpSSgSGUf7ecGfrk+
2qo1oXa6QP7L9dVoHhTOHK5MNRwpM7/M/m9cye0VMq17AuHSsA55E2oesTg7
toj0wLsmHyshyb/f/7IUvxkeMQJ6le4focsN3ztrOGyqilc+QpBS/KPZyKv4
PbOwEp2OCn4Xa+opPEX6x91YJlxSQ5/NFX9fLO/SLOjpE+xGIfMMxXsh3Zjm
SIT/NCxk4wToH4vlsFGwwKFVJ+lnLAVbeVgOgL5JyDCG9Z9/yY/qS2F9qQMS
WvzPLXWq89Rcsnn+VYjzfw8bTt4ynObYs5NlerjTtF768EF1bfE/gDxmvA17
/Wwyou+3zUdgJEW7I+Jn5Rkp1JShWlBTG0vNhiRcmlYz5juPVPYr+6Ddb0mm
0pgAh1ljUvKByJSPHPefXrskjnj6X95tTTacwXUONUO68CDDZWJ1NTfFfs1v
7rPFA3A/J+imXGhaNpILIH8E1011bdu1N2MFeao6vt1Xz5hvKohALQhivT/o
ccPJ7BD2RtdPCh+z6E1dbzUoOCXGxy6CrumXDM1q4LtuPZ+rJfu8U/zNrGzg
m8gOPcK21YFUKBtJfouOHzTCycdSpvS1YJPN1S02cEbFw61w/Kbf48FSRDvx
9gulTcpENQsbLSCo5TK/Gie1KijPcT6yPn/6o6xfuDdGii1hqWxMxWChfkwv
ycffEy4Ym5y7E8eX/KfuGdGMsHZ2+nRa3RahQsS6Qhs/S0VsnHQA9KjiQWZH
me4q85nCaPNHY7qzkwVIN2pS9reC46iqP70bc/Sq30V5by/b1Va67nN2JFYt
6L00/O8nbWMef1Rvd/5FyhYbczBdIFy50u2HZiB4yYWHqtGWDtLBRI4kEzZ7
nHkkgx5q2nghfpriujb2ktPK7uscXOtyz2NF0jgFczJtNNTNGDjYPrTaza60
x410DWgBtmqj3CuxXwJ96ZHPRxXgdp3AcwAiF3dj7R4FCGyJr5hKiXMNAkoy
rxL7SinGFTeyeDllNZammOn8WaDu+RpemUY9fqOrsS6Fz1ItcG8OUVDKeVKv
KHZLGLOMmTwgfKda+w3oHYbGpNmjiJi52W9AJ7nIa7OxWovsa/jE8xLFIiq9
yUJgBmGRa+MjWs8h42gFvuZvQgMc288vqmG97H8oHC1/AAs2SoFqfxWdEfG7
S7Es/0Xifl/vQmhn/TC5BG6+dfPhUL+4htjvJ4IHLBp9scijOli4Wr+9XiCc
K/vrD89VWhu3SLus26gpa8+PUSrWLWtDHwKuNozBu83lUQpBV4dOuWJGmQ4i
j+YaFHDYIvLP76xJ67QTWakEXzj7C96dZYlB2c8rI2wLu+FizULwwLp6s0JB
CV8rY2Z+le0lDVdStIB/UThjtkG5b6wtmKn6VauxAgob/AF8wuv8fR0frXVC
yO4g9z1DvBdYBiE1wGo6/DUyC8M3kSWfjCsP2RAkJjFRmLtm9AOLbY+9t1J/
Ubvvv6Tss5dYvJcctmVPn7bi87GCyiZ7zYWC5DY22s2T8JeDz9+VHkS2x+if
xjA++7X7vsZ/Nc3SPWkfExwwogNfXR8hQEY/mYhjFgfkkOsYAKnO0SXkOL5a
rFgAERNtJxTysTqxm23opBtlQV33Z35UiCNJQQazQ4o1Od1vqqO3rbn/UZ5R
NWVZw/nrcDy/1pPlQJlbFWxgqRIuJO9xceNnsDR0y2xw9Lszx3VGIwJRjNWz
DpqSB6cQ4+u+0PCwUDGkU+WMsr/3MqvSPdqUGroiRE9A6AGB9myr74YY1G+8
ptRj3deWj6zxlCZmN5kLS1hD9qILE55KmW7foCJvkSiHeUpKgf0InjE/yxT6
OJOTd+2x3r+2aDak095PxwoSOEVlb2sEKBC7VnXiYpKAGM5BBoAh0RLooKT3
tcU/T6+vNtz31zsRql1mN2Q1Zp0ccSRX0o7v1JiHJGrXsW1bMo7f1s5ATyGr
kRo4ORnU7kSjKISk5doP6OX3kn6DCYSWcMG1a2zjV2YCpNS/Tdh7upTLi+he
yj640RKmib/zNUwJMg6IFFkOb0Z/PIJuaecSLxtwrTp5prOobFgPA3emp4j0
RxMZRFT3BeEDmenLMvXve3BT/IqfZ3aVQWncPbB2bjcJUimpZ2YDuEC9bc1I
Hy30IniFF92YvoV36EHn4ddkdWY8/VQ9ENauRBro/6pKxYlPEWeLICAW/O/u
T1aerSpgGmYtf8WVM+OQwxDYg+R2bAueDEQw5pHUrWjl3j/WC9kD3QlytkXy
foqInJPQvOXJUFzyI+ShIkPxvw44ETUPDJVeruQ1BeGUu+fnfHV1D2tKCtfg
80cHyYz+53rMKMzSVNd0FiM2GP/LiA12s99WAYhk7l7DP+8oOecCd9q3+vtN
eO18BtHHFEzIY92VbPFoaPUUXI/Ps4s8yaAl9sgsNsVyvEL7NvVeCmN8+MuU
lwW++ufWIrgXTDNNwxFoCK45wJ/OhqzCDif/cyfQrM7PLxPYjvoC6QIqCXau
qCQiUGCy/xr7v2x7HUSgEYCWlvlI5g5cZz1mOVmW4SFfProb+x+xAThxrOa9
7+JDV3qVntCDUPzrSeuN6AG1pC84t9QLfuspdmvOU20SsN2BbGoBtgFSqWcJ
PTgMQJRFqOwtvCWej5KhA3FrBJgS1yfhHUgGTuyckGNYmi0My9nR0k9XzYJR
qSe4Yye/EJHEoN+9FEWQxzapD8hY0/CtAHdDglsLpSUM+iXNe5FOqJN2c9AJ
A+y/RtmM3efTGura6cWjvCwyii4y9kJa2ny3AXtISkz0KvVSEHI3AxAQgOXW
zcsWKr5ZAYwiEGJUNmicRsoiJqMFQDIkqX9RMNPUQDIkYWACKvefTl1296r+
flMksfSMZ26GfJFEG4FVoz4ZCUwSDXClZCLyIZEcz5pr79XvGkaOvRsLVX2B
P1TrIBnLn5qs8aRtrJHu8yTO19yNxpJ37l+n0W6kMI8kUZ4Jf+Y+KC7R12Nd
7WsRUgXTj/HXWP7ltK8BAYOL/0M9l0c6nVyXyjbScDca5Q4T7O65F6P+M3yt
2GrUOhwbepWCMI5QF7wJT71mV8A6Y2td9N1zXnEOGoMfTN8IzLcWxhm0Zdtf
3gmTpjqXQpM2dRZ0VJ4XjOF/q7f1F4zpli8nWSjRPxpRfKqs8LTqMmqj0KEo
TSphXmlDVyhbaRCKn0SHcwhjPFRRXutI5gVrwy+fBB9sDdb4awmGQCSEtBNY
OpBYiQAU+Q1SciRlaFzh6mzJ470tOZY5WJZfR6nMvJp5M2rI1350MyOG4WBl
vot7AJ9+jzdaGysJcanv/2E43SOcPslus+9VfU/9IA7mETJcr2db0jyvBQSz
agNj5m5iWKfHaiFuvA4KR4Kr8fJBIfJfwZrOlHkkip3DpTEhyhFjf8u3Hmqz
CIGyFza1aNZl4jX2oA8tqBk15XDG+bfMDZAa5aM+l1tAJGI/X4xL0TM4y4RM
g0iC+3GKcJMACm87tZ1hFIZBAtLLxcXNlbERWpoKJCBrKKcGvXq9fWQkCXDn
y1QW9paGJP9u49mVTi5oHLoEgzDKZ6JSQh5+uw5czwXkaUo2Bv4wlipgdLyk
xip4+5fhFlyJvevT0/AxTv5mj0foIwPjU1oRnEfLOXaN+MfwuohRvhRBh/wJ
joZqzsc4KNny4M6SoLOvrJwH4gvbAo9q1xLzN8XJPXfI56eC9Nw3kP0Yl/b7
0ugc564JaAZ0gcuVNCOZDimE47jC9Rtg0AgDDmA+NsSvviCjfevsBQFRcLNU
gC2pufdSKWOkqZZK8afHdm/3Cg23zl9A4wnOgmQEad6HtN4LqSY1/ISTkIyg
6nzbnQ00fYtThYIKW/jaqAScMNxwGj7NSXMlqmSD0MHiigosZs8YgXLD6PkR
i7LT2DpGgDky705e1NlbAgjtdva7cXBXtir4AbOoha0hfoiD6QurgE+ptSnA
zigHYEAJw4RPtxyKAww/K/w87gpcoOGlHpzsu0BCE6qKwNBNDyjC++yjDX0N
Iz2oS37qi8J+0DREqN4aS5D5Ta+0qWiUZOBjfF5n9DmvgENlIQx7V/PshKSC
uKFIgeu+38potT1+qZ/DPZ26ZWDsLxilqN27b/TD15cbE5T3c8y9JYSrVbnE
KHd6vf1dTUvcmaAcfktAFdgtWQOxr144+IWSO2dxpZ4eDcNVZj1Ydl13DK+G
2lO+vDRplkSCBUVpPoRwTANOeL34kkCRV8TGCE+0hysNR3ZjyAXdcJM9tnhY
aI6sEcA3FRp+RvfgmXcffYKw9EPPF8vCiHT4CxSHbEqopKsdtuBRQFvmnwJA
QERPxDGRRbLOy/FqS7AWY9Zr6zK+oVg6bnuZ9dtb2mL28LWmO6bU1okOkqX2
FJgBubcXo6FkkoljMG3X0eKcpDtX7IbhdNa/jq/2QUyDoA9TP5e+anZj0tTz
ipGLOo1/Z60PnqScySkOfqvxbQhitM5DsxYwnXR5BKjpaOK4jVSOknFi0Qyt
awoWnp2lhSqshQnC6Cebsmx+ivCnouvD55rPQryVDuafxhoGNbWSdAuHYBFL
iy3iqgLT3MjZixp0toR+p2AnHeg6nAqFLaHSzY8l6c6X72hR9SDOmUQAcaZX
g4XqSZthdUrAoe0FGks5Ka0hTPq3tAEjTnC3SefwRpeY1fREvwGABqMzWXcK
3UNSRvrI4Qawb0eVBzhTfxnopOY3xKTemh7IYSmALouUkvdf3UPemZaeSoYW
CEQWo1kvpOfXuUfj9fA0x5QOYU9QEO4aOCicSPTJ4BEn/KZ+oMWI7l+GMIxI
AohDUN2/0B1uYid/tEiF2g4Ism1n/qymovNhbITvlncGCwFRaubZ0HSCX3n/
m254PTZIhxY2VHycMSSLe0FZBlw56cYZmTJNLIk3m++Bz/a8N8O5dsccWqAz
/J/zHbcJskt53rwrVe1GCqVMd8GH5s0/af0jyr4Fyyx/PXDogbamP4ZTPiHx
546Q8P4BxzR6Ao8m4Sg9aSFaZVcjr6ZU1wNtdEDPnVus71XG+n/qlEzvzPIl
w+RChJeOH9C1c13Z6w98l7N/gUCzBX+OuQW9C7AscXY62IZPdvI/kRnmF4MF
ydd3AVhXmJeF8N03qD2rGjR9ljqNA2eJPjLr2GSn3LibWvmnP//TXPXb5iL1
9o7VeFS8TSCdKc7KucPYfOygWGo5gnNK2lbtevHUVU5rcDi9UZMbp/57ODPW
vQ1i8gRMhiZWG2DzV89fvETq4mgyAhYt5lHcIaFNVT2eCx1VeHwAPuu25AaL
CISpNPg0uMMeRDUxVw5srY1B6f8KpEo4y39MrbGPd+o2pxXXUsm9ySkzCw+5
JkRJrOd3Z77qXWSNdwtUCQ4WfAKFLKF9p+nUjLnzHXmgDhIxeBsjqyNh2SMt
j2lFFf2QRLJZupjh7qg+F7HbsPB9EnFJofVCBs7NEsMZPQJNY82EKSBWSf8z
AmJCSALNhoH2P0DKLkXEuCqwCVDlbtJlnEoMejwogtU156h8tLnSI2sKLBcL
9JDiRSwPhg5gv48XIYuUd0kr57unWQkURCoMSPHKG/+cNnzw5HMsZSgiYG7C
x7KElSWyo78dONYAr3feAVusP5kioPGdE+f2WVKB6vjg0MXIpSviS3Qlh8Uh
xuiIwqBjd+K6zyZjnyaqgAgK32jS8Zm7/AmipeGvQqxjSe/gGTfCQ7BrDts6
0ViZN5y7JJALqud6qpO3hNtZaIHsSn2wscnV8LYFYMce+sE1hUUCKuSvgERU
bmWaoYChVaXSihIahBB3nInKdOlmquufmPxmUBlPD1gXDxpXPDcvz9RdMc4q
bc0Owgoknaks3ykOj0gzvE+hCGi1RBw0ImPcxPBWtnyQIuHa+HE9MFeOHSIx
7A/SeOlIxEGNNzUy6s4X2PcsEXKm/G6OZ/MObSK0QdFV8qQIViJrUgdZVCtw
8Y1h23+k1V0MBPN7iH/wWaRAEA6dULVrFsEWx2s+IYWHvD2JuQlv4PH1u9RP
SOEDWoCYaEAoTidboa2Cyd2gmrzdKVsT83LI+MHUg+zFiqOMTA/PWH+6E2vy
OOF5aVosKd5aUmYDnu46mWXuRaNvFbJu1x5iK8qvBZsVeSseMpp1ixqgYQSH
pI1PWLa5l4Sk86mvKSe+lNOYjHlR8XxOIRokGIQKMZAQQpF2/FTWJ7jo7GT9
GzSvyUe7SpgrTYj+m7Kr+ufTF8MfogfrdwOQNf19Vb4CsOpULOF5XTvBQ7ey
X+ErQU/86aU2EswYdgLgcyjPWWd/C8K29F+w37HsXUOQJJ5dqvRSk0Lnpu2Q
O/ecnaR6IzfvIEKVYmwmHWY64YBqzSvy0KGFqumw6tTiydLmZQLGqE3iwuiW
JY0qVa+ZRgHP4Hbchf5NVlDgkyEdJ70bV7x+naBZwzhi7wqD6n/FpXAOCgBz
ORFedauGTUIiXNJzjgcka3994hISxy1LnrPMhHIFVkStA3Cb+PlCG4r6Mhi9
hXJ43x4zmgQ/Jg1RYm5l44dUtyRRvWNmkCmXCzZpSp/1rVB0K+a8sYbwNS/v
JrFT8EAyCjmyaIQPOOXGTSTpeyBLRkMI02ge0SIQ26qdjnkdQS9OG/PbwHDL
XZCx+FZNZeiQZrRw4PzPOL2uJW1ghFemQ04HbwdeW7ymiSXDx482KWatT2P1
0mIH1tZF+A43vHrM8JVsZ7/U0mmT6ligmCPYRhFMX5p6bVUk9OwT7i88h7QA
HvpoVMYM6nENlYiDLfJnsHs7B3nFSg0WBY1RwBzZEYx9IRVxScaAVye6fKK3
mczFY/aBtXLMjP5aDwRfoZG8kvxTj5FB4w0LwuLGP5EnUZWZjS7c/bExQBji
tMRYPjvkqoyYXv03FHmY4K+z2WcK1nNcAvrBwLqidxS7rtx1xOnKYs6xVGd/
gpm/36oRU9GMsoAmFTHvcZPuS/TD0SuFs3XTM/b4wmu2irrt/FP0rPjmeX6G
1LzrJbzVvqwQCwr6YtHwTOKFFiidRmZg/kAPj8Kn0b6TIjSCHpvp5r04Emoi
Ky494MnMKSXS010CE1ns5ViLMUpWN9u28DivRtDJxAAWESptT+XEvivvALP3
2rjRDdS84BNY42ST18Xj7RhcilaBkEtTDkmqZjn3ygShrRCSAkRohDeqBOn6
o5IET3p+NmnxiewvEck8T5GDfgZJoqaBoRa+nNMWjdcPQwDJ++2uOISYWQ23
+m7ppiXn+yuSO4cHLBEKk2nVNrtU97q+S2QVx2ypx606kgKEBmoOaFCwDUFC
Au1pNnKJ4l7cToJQTahhXGYfISpv6P1TmQevLGyyHt7bFD7r83W6t6LZFQmg
Ur0M7sRq2yGlZyDNMYOSvj7ElnnkMN5iPZLSrI/8O3WSiBULCFhzUOp66ADJ
dX/AdgbyOtC2Iu1oEeSExvT7pPfV+Q+0guGAfN4hiYR82xMcUi4u7Hm4ZDiI
gLIvfFtzvVFyrYE+badG830BAiJCU/IHeCHAzLLbsnX9jiB4iIuCjlDf41l7
a2IpQfXf5/DItAIzri1JLsH/mjJZGNCstAJxiMHVu2eeM72GBF41ZuuxviOF
mlDC0bkASH4jZNCXse6hvj2cp47neMvu7fp4IYdAZooZoApVzAfjkYEFPuUf
VK+D/RATpDSRdJCEaUdhQSIMZdJNmQBCOzW9hJAfCdgeZdjgBvNpp/T60mBf
mxKrIeNbAceB714ZyqerbhaOvr1bMWBI1oPUwzIllXDUkOPe1Ebi9AgzLgb5
jpsMzXojqy7sMD8g2/LYjQIBXu708jsMc2z1AInrU/unjEbhnQIOx3MMfaxQ
xBCZLb1myS6iXpH6+3CsHwFPzpuc6fJy3+lJoZeItf33i5fBV+753nSnRazV
8AHuNSQqXD81TQUEzhUXR/egjdM1pGB7GPTFY0xOBz8aF8l3TH4mj6Lmsku9
45kZHaUKaKaof1XbUHGE0qCMcdK93YFoWRFGOouzSNnsPA4fDt5f47oCWNUR
haHPLtsdcFDXGHObmpk8xe1tIZTQ4brRpk8PIOHiH3DT0BIdfTpgjVPGEueu
qHqTtCLabHz6WsJdK+919tb+isJ83uvHzt5jbDO/NmDryS0pW8hBxKUp71cj
Q9W9wbXLfqP7O6W5WqoF+AOC3yW44k3AVtwMvCelbwruB63VlkRfm5UKsWY1
i7JMkKmgtDpJk90UTI9qOvein8P7b5SbE6o9qvlaksm79LvM1g99b5d0mwcj
dvU8TPWdNdp290i94i7FwacThnzX/B8pMKISb3fSH0tM3vkaO+BAW6wsDcXq
89zO6xk7GpU9a/BY7vujj8tvRl3/Jrj9+G/HFnwh4YK/XOjCpqkfgtFejP+U
K1+NtUDE3qmU228ClaEwyFWgV0CiE3S9d59hAY0ZhnJWr+H5JRiOar4Exdw3
WG72/MZ5IA7WfzVGgWQ5vB+8gaAZSw/YVi/e9MIUizZWFkp+RykBbVmPneib
9EMaNiHzzd78+7MCrz0PJJhrynXyPYNv00vZxWxVQz+J6I/DSANDyTJ0XHqx
/LBGxL6vPyIgmFT7joLkemZJORK8zKCmeMO/vWxRvr7+gP1SEFF+G5MznHgL
q/JWxpUm8yoviVy2DW5CdbSzt69olwo7rxyaxrP/dfu1HcBzarfLMwAwL2cM
6ehMdomJl84M7OrRtA2b8TNZLxcJOrde8X7cncMwnn5jFKeVpb62ekx3ZX/j
A6z0MHxgDkDiExiKE+yHzWprW0kudwl8RzxFAYHhzgcsrdaqvt0VbeXlE3pg
pudAhXmooZKUwTqnhqKKU137iRyaGyvTfD4KJDCizgWK33oxLCVSZbzzIHfR
5+nx9vVnpGrX3RS2Iy57CBrE1Ce3BDcIcplItU+AsuvevsAbJt+/ZktAt0la
gTpZB0psILDAPbtahHb+Ym/twx8myiE00F5/zQmYidzvTxs5zZw1Da9pQfLD
M7f/7QQKc2ycYa99qG938XETS/MwyuZKQTEuatAbmMH8tPZtEPvI0dbk1pQR
r6koLF16M4uNaZjYkadl8tNHFkoO7c+IjrOoxiSbPAdk+wW9uLFTV4c2gte4
TFDQCy7J6D2Yb+B/MBWjXMU8qMgVuswS2ilWS9LIRQJlYzK38tfybhnFLFMb
GvBimPHH1UWkFM0hzCWi4xJgqshgmbK7Xnh7b2bJgEXfaapuXrxzwsY7jOJy
msIYydLhzqDy6XstozPqb5/+9J+sokv2f4f0uGL+TTHFZC6yVoPcreSqkGa9
+JwtrpJiObQ8oTWjHokOAhA81gsiemW+ekbrgYskk4iunjyfh/gFK6yHSspH
7eWHkC5VtVTITqKWsDRrr4QYIqUFEtjq7KZaq5C5aCEfJA9hpfDypnM7+8r3
/rpRDjWUaBmPPrb4uafj7AvCJqQ6jKBsF2v18yd4XhW9d26N4E57oTrsaK7S
k1WwkOQCsK2XuwaZ6IbV0w/1sN6CbenUNHkFDO9vNFPdXlX+pnE/p8gu2MG5
HQr6X8TvmUcvxSsY/6tM3HPPVVzJqlZHeHjR001H3qu2GCA9h+48gnRNFIsz
A4ZWDXMk9WxZiuoHndZZctlv+HA9lVM625UI08e7ZdHg29ZFz5FLR+UuXvJR
pRO8yiEZDsKeG6/7JT0kObnfQpClaP6946rAO+mh2jUIM1dFPnX1kjpY7PT3
yMiFFuAkdESThLwoHisJ7+li98xDkrj5aEEY7jC0axU1eskanUkDHThcM1bq
mOl0iu4WDUgBR+pwt3OueCuNODR33OBSQsYopxGVTV5gZAT8vFHR8J7UEVSs
mGtZ0t7H8Qt1CwZbzHbYTxs8CwfSiQqa9+/PEC8ytxNrte8aq+MxtnWHB9oG
ES9bwrjf8JOIT7HxQhRfV4p1R/s7KZBD/NY6CpRtfEwu2bjqqwDBoaKS4lVK
ST7K0tQvUY9sTnToRKOT7ikRBaMQuqrqRKh0sZI1hx46wgl7IP5zTjLp9TjC
NzPVBXRKXgjn1L8TZVPCaEcyiLgWfMh8UAG9RDNFOrmdppGCTw9lbV39xVKO
YbP6pXxiQ96ylHrav+w9C4vsLMmLFUXwpNDO3V0sROthjPQRska+UX182lu9
bi2WUEWPqSCl22QP7/FcnoClIWyetBTqqeiJde8YETdGduUugJatf6r5nEgt
FCeeq2DzG972FQEbZojOV5ZAYS6eHbMh/m7+kSZxOaTnAfgq2JvZPCIq3u/5
wxfZNAJdBnZN23H9N3wqAMDhImwdCwGn0g6q0ALOU8po3az09oa2gd8OiuWA
J8LQOtdT4/F8mbgBBN37O7Cy+GmgSmuT7MxY5vzS+YiwcidGgk0jp7tn2xLu
rBFnQr9tC+3cS7z/fvOZqZyXvjoeUyS2Sby6go6kw0JDa0Rhdgev2BFvJAId
NcCDRyXC/frXHxOw+eRlOKlSvXfwLzqtY1dHpqoXpCNIQ+EP5IRyRTakiHss
X5Uic7xrwsREEOtwgSB7BIAzA2xNMz9rn6hRxea7bQYC2TlZoHmVFqlm2Phe
Luk1UkBhh4ZV6/rQ1UVBPX46HejE1n/bVj0n2ZjFwBNd3pF5m1LPfG7WCnBv
f8dOy0sToOQ9Rk3gwgfAQdiX3Nm2a/nJAbOK6SzOOy9yFL18ID6jeKM28f1F
Y7y8MT3UEVZwS6KurK3t54iWp4UHRhZkgIxj6F7PraSk0WCjNhaIJ7+tL6sW
by3QkrS6fJsYEFJo23kztNlWucmNbCQ80RqJBbBCBEKkvnobmjYtGcDJzPte
ZkNXu3MXTz9mc8/OeiHKFiQKIWu3HReJ5Hx1Pjer0udkFSlsr4CD4MQnB85R
yOXp9eNhNeNM2WIoib/IEgZlSAbzqmxlCY45qK3YiAsR8lhSahRTsz+raVLi
Jkg1/suyxsZN9iHnGFZwT1FV+X081zSIfwxDdrkj6qkkKIJLWlZZn6x+lx0F
NPaDpDg8Hs/d8ABHjYrFkYcn1hlLM+QXVP5dM9kSwbMLSVHJ19PxCOOGICuv
a0f7VZxfixc3nvxGDRk1CCa5HBnqeXG4Vg96S1spVdq1V3SuPgF6nFjyw0xx
Qb6wqhHrw6pv9QSf7XSYHtskLhyrzZkVVakP2upzBc2QJj4MUGXNDSaFg7fm
RqVzWn+GKcR23GzvwmUZelowOgMu3tagPLRPxaykmwQWMbF4ThihZmlU9wk0
C5WqVkSOTMob0GA/RS71DxiuQ3zc0iHsi8TKRaeo/DiV5jbUP8Lxgomr5hc+
qISsUq/5HCEW3NXU5N6fZAUrUASF29QYQcxYbT1rurDE3cFz0w3BljIbqV3j
q8k5ucxAcIT6bjnwj1KfWyMTY8lxmmlACgIaKzGk9wUhjDz/N5XMBt/T4mMr
KodT6UUxWUVkXWboW6MBPfH6xve/9kR5dEp77uIrDkHld5zcHvn6Q6OLW3Qo
nitSYddrYdfCJMcK3vljh80Q3qdRHMoIl3yEFvf4x075TsjGSugHhYyerdWS
ybkhgNJ/eyX6db/VuDW3w5oLM1X4pg83P55tNoY2QPl9OTW4OhDCvk0z7SpB
3Wwe7wmtq2YYvr8hl4RKlJJsPBqoZGP7inBQYGRizx7+k3u3AJY8vc6TLFvq
fe/bCYR0HGUYIMeQdm5D6O/q4RAZRueJQBVl/scfEqj3XwKKEH0N0m8bBBGP
s5qSVTa5fVTKcFbtPAdxZTAw4wMA3sqm4uw1MmltHfSMGH9aMqk60dPGA6dy
UtC+aAzGHpf+lOQkq6kXo8iw9ydgTjUYsLX+BVGM4LDFHqFdqCVe/huCslZE
A7kyEXXpxVArK3mvKAmybAwpyknQoJcIcX3TvGdphty34PajwIwwsvHEHkwe
/txM8A1lp7eUw7rh5wVfiZT5VV/CpZGWvA7V8gYc3Z2BKtWPZ2wcavnrlVDG
gesXgbRUB1IGL/Yh+Z1fezgiSjIbHa9yoLenoi8pUyNgHOb7CCMa7As7MQat
obst0zA7Z9i0yIwBiBxQ7r5kmiPYZrb0dkEYjLdFjC0JrCmFqwbF1n61Y67q
hiNvKxY1gAVhOCxwfvLeQ/NZzS37YRjTeYqWCc/JQ/tAeJP/FloN6hhzqmsq
CCWLfarq0VxGKL7U+BB0yCIHCzjfsWPm/cfKkKjhljyKf6UrgPe+EqscLcyP
+xKGKmhhMq+tdmjf3POP104kazwMjhv+2ovpRo6vI+Pz5Y2nW3AsUu7z8B5+
8GvssBPse3a/yj0hyxnxiYOpOc20I+6Jmo36O58MM7AreZqmca9lZqUVFhXo
2q7caUXjRm6spAMTs0E9M8qZIvWHETVP8f9Ep6KdknffQvwuM/IaHX2JQogu
lt22b0/ZNa6Mt5TlRMH3d5eCwZt3/jSFDhevxxjO38Be0zRu/lGBfNWK3ttY
fxmIqF5RUQKdrsxQyCfZRgmr2Gop730iBPDinejXsdiytxsx6azEXFUdFDpE
IaZjpoHi8LUpGxpDGDfqz58AVV5QHLwejMCvJ8ed3ovTx8Pt0O/fFKgnn2/O
0e5XrbKx7uXQn86WZ+HXktfZbF/sPRHkoK2fBJ1FU/UXqAR49LQA99XKYgXF
vr1CESfQkt299KB/wqFDaN9Rdc/7qpChNJuZUyq3cQ72UGGy562cNnCpC5eP
QpUgV0SsGadAjp8Oenwxb8Z3X9s99QkCcgTy40ZjKxCtcl+f7n8IM6/e+zqg
rtPZDKTbqV3VtfCUF8hdY+5TlG8AFCqKkOkc+OnuTTyVGYvvnWU7BXwCGdzA
QGPdGUM05pmnJmDwg2bMiTCEPquVjDxWhGZfheuq+mlMubhtCspRY8yT7BvZ
ihrNf3rLzszeBlWRgMtTTMtlYJj3S/JQ7gSeUn0Ph3B6wiDbvYc2onUnf6dB
UvxC/Dd/0pxqkwT/KFVSNN9rRZaDC1X7Dyt0mu1XWvx8I5bdaIIuzVSPKUrq
5B4uYK7X0DFV+YqHGaCsgwSm4MVz0xoV1shXUnvZmv3EZF3ziyjVK+EMGVH+
+/wMYUl0103JjjCdpLaRIHEQp3QsXN9owUAehIe6N2JaxySPcVsCPXtpS15O
RUfGtzTu9Y9xjX+vGbRmGedggFmzZeuvyZWfFx1A5aTr7plotpiwhcgmNQYB
5J0ddjcH8P08px/+1pNc/Ds+3BA+JkTzril1b1RB9SefUsKLQ+E0W7OM6quo
J6BLjU3Mdo3kdHWMEIGxoltOcsADrB1a6mVnoIPXG3lsCX3N7fBZ3Xdb2Zr1
Z4Z30DSwbY4SElrtk2HF7Uv6XhUcpQiVPWiaF4edKAeVDo9o8pHRgTZl2Tmo
xvrc6uNIV/PJmDjvqnWnLdmB4BR1/+LBHie7cwl1Ej/213LpAty85hHk9JLN
s2DlKbA3Lna7fmOwW5/4JnKQWZrW+qFvvUXt54lGqFaXKvs1K3ourOOVUeEa
3ohPxf2dqIkWxg7yqxtxagX1jEqI3tRP7OG5VssBCcMAIfSRvP1MPaDLVa89
U64SVp2lDcB2OqrUTLUJhDe4hmcph6tjTdy+YuZimdzWYUL/FdMY9M+IdJX2
CgJvSZzpLeRas56I6wa74ucIi9peW5JDPF0XrWv92CHLo+5Y8GIKuM/I4B5g
sYo7Ej8iVoOeNfR4xpKUcJ5gB09HW5lr4BOgD1Gv0jb6aUjLjSU4f2PlmH3y
GFdU3l43boYNAahZe5WM17ADTXOjSEzcNWGQbKJugjGDt1Wzksiyuj8dafmA
g5150VucUaaBbK/GVXtzs9xCWoSMkvhhNMVIm4gwn/mpy0SYq/GcaM4f+FsO
MAQbX6SC0cka/7BIdGY3qSBNFm4Wc16f/Yo21m4kVdTKXLIqIshAKrtDAjsK
IMz0enS3LZczofZRBYoE0F3cB9r0hpof5P5vN53gefJhouftHtZ6TfdA2LWW
WhoDOd2laE2WWpBTxn0kRhP4CR/FS4rw/qcSftP9dfKw31aqOWXC7/58e21m
C5Vqy84HV3iu5wFmRqzzwA9oOMXIEyJfBWTbAXzOlLkTxQlDJCYTO2caUFnC
U7FjGJV2FNu9uafRg9fonxUkkvH56GT5NGVxnYIlEHo=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "B40jvh7ud/ahkCWXo8CJP0S9JYnc5+J2pwOdONjrEnmjRzb1YpxBEP/gM90XdEQFf8e+9j+GJABVN1VA/EUgHmy986oXHU6n9uJJjaeBsR8h22iSaiy//95eH4kKFakRZgkZDqWp0dX7AUTwRg4vZKk0rom9cx0xsiuc1Ki6fTzxDmmuuNW+yyxk/luKJogixDl7f05H1PhFx3JTfD9y6cRFGovJ+RtyYHOBbLpk0wgQfkH0OzPj+/xnj0AVtKROMEir0zNAKk3a9yBDUSAxL6mI4Lxdz5oN1T+WL8Dy7VHsU5H/eNMrckvLCUoXHakMik+wasTKl/6CijM3xnBTnoj5fHOXKvu3P33I8JTD2SHBbV6o0aM7v9YezrOM2tAFiD/30BTPtuwzjVWMLw9G5M64+eo2cOlwwhpuj3XDSGsF9b5vmOwCchrgUvOf+w1L8qpf43gIJwkLG7xXIUpq3mI735dgPrpWHKU1eiqTE4vcQqDD03CmQ534IuHSA3fw1kBb1T9oVQzj+pZjVpo4f3llwFXViGYbbAy7SuE8bJtlBwiYsq6uslQS259GMV5RH51qrmqhsy8zu0sOp2/s0ecf58R9xUvs7p8ID4GvpUIhBQLtb5xwbONYiDwzYgfitny6iRTn+R1AdEWvESP6HB38UOnJsNG7pIm3lEIH31j1mm58dp7V2t1OEJ+HffUbOUGxji4rJewlJ/8yaRlAdEPAvzV7qgAgJTSBjFZKoAQH4041+S0e9mVer0IZftdH7MILPkWDql0o6kcdNtfJE5nXZhzZFWsRBYM6neUv9uvA2HMvqyLiSHlEzgnyScwk65R8ZLqGomUqjm+D07xH2LfMdDY9qYOZhAbyEDJD7/T/Xdj+l5DGON9ROstEQGE/7fVuZgEQaRxoV4Q9GgBpazYSuhnw0brBzrbFJRktWKyIaToLs29cRnFiAMiKuZhUSGKfw/7ivcim1VCy1b+l6y5nnmj1nBhUfhYHHYIJZhHvLh0Kw21R9WbAqUDwCxlt"
`endif