// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jmJnYvMKSr5B4UNaU5bWQch0e5KPPavFv0XHd7zO+Z04Hhdj3vch0I+E8ly/
wROSav9yg8YBl+OKUvbmZ9aO2PGMhhzFYpJ7tauwI9sUBTpbNXRu7FK0RDqA
/eCzbomdgEQxFoAXm3f1SNuQbXIHnTkyTeLpa9+IX1NXFZFa3J7KqBvRoExr
bOMJ+egfcHlIB8xOGWNi2a9f+BRadtjtr6jD0NWOvhGDOFno9lIkUbkPiSZW
K2UMb6+dF5Yyf7tNG1g00hnOAL+PS1xoMQ55DKV4y/fb8yu+l9m9a/s/w9dC
nymivPXsnHjacnh6M1UQlMxvLj8bHtTA+kGq82vvUg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CXmOn+HD1s8be5yJjQRDtdV0Ec1PaIP1JIXrOG5sm3VYcoKn06QplGqpyoac
2U1IksPDHBqdp0y0eUT52IDlllitTazCDkmbiWR+jieLo099/YsFpOUKrS1f
wxjOo4ddy4pv1NU0Oy+v4CaIlkrfWZlGFofMTYn9wssVSSTQR34TS+8IZUup
Kuw6fHKNFyFQf+UD9+Ij57nQ8ZA+7uJULTt1S/6UkA9usGh/sHKI01gVIOsA
dpEM2Q6RLzQNreVXbrE4Nru2OvqtCSI+MmoDLyU8oznv8R9trfEa4ahgN2Gl
DyvIuFuAuKpjUBHfOu5mtZZ5wdI4gSGpRvv1jxqnSg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cXaoRQeCYGofHtMd0H44Fz1n/V8wAnMmu/zElH4CLm2f8kA3T9pn4rhFZk4Z
DOoKllqdBXMxETfhSHVXrWnWKpdsxYacovJfqf5CSCLJy+Ktfg3m48puz9CV
Zy0qFNUykpXHbAVVrgSCIfER7ysXFXJ4fM1BRl/XmvrlVWYFB06ExpQuqzAr
7UUmjdOXg67MliHxy73aVOEU/woncVBXSZmwqAss9aA0kNz5m/lwMAGSDBRU
6jQGZoGrxofKBPYQ2O1i0i2qisbfWrO7SPV2NLBHWvTVCpUwz3BxGVM5JFeg
z4MxjILDXLYus/iNMEtt+aJtc26Bx/cfOHEXaczjOA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
U49MBtZSi9sdg+M5g+EHccVPap74KEwR26TB8HJnzdhKvUbCDNfAVKEEoYki
JcfC/ZCw/306Aao5tVNmZPRlnaceXO71d5jVnk65SF4rq1ARo/J6LA124iSO
QstSx2doRC+jBIaEDqEGHSYLYS0oML5bvWNDO3ixqkVIly+3rqjsEPvJISBd
xgfK85sPjS2kyvkfaBEkGLzNjeUXa0HYcCX7pcNh5j2EqBYOoaVyzcWcNlrb
VlYMC/Qhc9Xxvn2K2HQYh0YTvaKb41lTAUQiTXk/KuIKzBZ9yHoo8APigxbz
HH/irBTDfdyPvygDssHHukCiUKjyppwdFCfROy1Gcw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hzyWa994XyjtxF1Rf2/w5XFilyZ6l25v2VvbRGb1XaMiaIYX69uwB17fzT41
PmIrxpl0W4VB+/BZzfPStJYymJeJ0/t757tWNTQAf4ox4rLBZSy+VZqoHyLO
ltcpUJyEYr8H69PtxCn/tg0J7KHAFffP1z0vi/4LSawPBdMarOQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
B/vOaAu7cD26ABl2OsIP/3NJSzmRi3Pe28iyKSRjEHnop0PplX3VGFmMJgIb
iO2M3ewqxvl4Nrux/cIJXOKudTFCYuYKZY+DYjugVcpmQdkFa/3woRNLHRiZ
HI0IvpwgBRtB6yGIas5hNtHmzl2vcgeSfdH3hES2upkx8xJJ+DZ2CVwzxdJ7
8AqYdUwxQSP+Nzqzncq94BnfPXRu+WyvQJmZzjV4zexRAhNqJpuflKid2Y4t
ku/C0+2HXkD+AWWLbkAarE7cUbMHNMEp6gJyFI6Jb3v20+3V3OkV6KaRhQoQ
Nqtxm7DQ49gkZOqJvrsVi9k3NApD6wv5vLSf5ByDyi3HTnuM1ZeX04EnsDBy
WTz+ziaz/wRSpOKuwexU1Q1i/TQXxeyZ8elvv8jvMqL/X3vOrDXrbWDfh5bL
5rNcUjS6M2XZE2yd4kl5+NWGZp3dnqvPBlvBY1RYOdxTZZA5MprZItR2u2Mc
iLVPNAOWWXpEZvivFx+9X6JVE5/PIyct


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ls5ZUJO48fr22a2lRco+omH5DQ8v1cXg0i3uLnuH/ml14wz7mUSAMCgZwku8
nGW05BZHbaIlEOLRn4rUArchLO6yXuPkWVGqqJgsHmdRD/MylTrPij+Ee7uh
BorhdJYekeExuU2lpEWhFCZN8AErd7m+VwpGA9o5tP01ILDrVSA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
q6AgGuSAicBAbIotEclancvdHFK7uW/lVCzSD3nazC+3ufEnB84wOPfE+ta0
fwEraRm5/ymmQm/frIfqoj+2pTG6lKHejob1M034Dy1k2vNljMQDi8fkY2Ib
BVgBGMRm0tYGk6LBgwUBGvplG8VnRSYvxvh7/HhJ3IT1x20/z+Q=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9472)
`pragma protect data_block
mUXUNbWSOzbXTwKl4FnZ3gX8h3Dvse+nuiFz4Rgr/p2KXVCVgu05B2V4SFlO
dbJMLsHd7+ezlIzRVK3daKn9oDGBwANKy/idKpzSahocHe+SjaxXNf1v3FP0
DlwTJlho1qHVL4mJA/Gg2KBdt9CgskbxnoNPE4y26d7hona3rx7oOKfPyq21
Q1+EHV8ZWjszisR5JN8Kz+NNeNdmTmMnFjjndXrmARLKhZ3Nb4buNrjYrXEU
lmqLwjH/BntWlzqW9GGxQ9pMjG3xeN+ZFOnHsp6+iLaxdXsZ0Y29V5oAQkDm
fmkreHa0VbjG8tLLo2b+7B+A3wlY+QBOg8UlKoZkSIX/q0UZLNDTcgFff/S1
XR5U0X3oRXaHaCnYKLVowuOnFuRPc3+ba/rcXTPElG4CCeOi7KpLswpQO8KN
lsq3PmuJ34R3frX12d3xd1XjiC2nwuDawek4H7g8/Q5ChhkPDeLTlms1nOCW
unYWyf9hFOmWjT2RNyC4Qx17MUQFa03bjYdsSyfBZIPj9M3vSybK+Yvys2I/
Yvs9YJSlpFrz79pPoBsD6l9cHAeqrkXM4mqHbU3LNWDbLa3QOe9pZXNkCwVi
2j/9ivFgs7SjkO4J0cvDQYEQ6ssUEeOLkeId/1NttUosxI1m5/9UYpdgtGqS
NbkI8XrkjoEZ2ngKzKOt9qBTjSfpZDHe1oXA+PrdmeOKNnlBuLOmNX2xkIHL
9im2MFpJmj/Af1xooOMv/BIcrHkwB0qfWtZaRJy9Ulo9xGiRoT2BzS60Xs6Q
lv8uSPU1Xl3kWyMTvKbtEeeLDOJ8lSHcqCRbL+tI5kc0h3+0vVb4l3WjiViY
N5MbUgjDsjh/j0uqKvsopFBQtufcUXSRHAQgRg6P4wMdjfhkpNRcl2M6IzHG
UO2oujnpCZRcCnMAYZlZ/MyBgo5RqnWc7ZjJcrj29rxFTUq+J1NePahE/RrJ
VBe08RJDqiUNcrz1LgGm9UNgKUkT2Skl4xANivaLynqSzYxgXPTZAiiNAy/8
iy612+hOjsP6PCix7xoNg5WDpZsWgjJrULsv5RD8j9HgMUQUbuuRWvURaZnw
l0ab9uyP1mfUB6GGCuTItjftr7pyaqs7V7icYM3hrK3NuqhHcF7D7QIkHvH3
1oKUPsGI+BzcTzQxOlFL2Jf5ic1cDzpOU5khsvi4rNmrwyN5ifzrFzfyjX8r
cRvdN4oW2DhZF9VtPvB53dk9m0KBZ1Q97/EtAuV5iBS60Glk7J3cPwbXlNWp
BY1z8jKqxTl/x+V4CuD97/xbsBTIOIeMZz4VivhH0/H2UdaUbQRuUoMgS7wA
PHXGaQyFudotmWb9iX/swVuAoxd4Ll0J/PAJFuPvlsI82D6FTYV3bOFWqzHK
kW+gQej2zooNa5eR4qEHOfC2XAHPUTpb7af6Eb1GXPYQ2/hHsgUOHihwqFDM
sp+s3HfOUeWCBOoEf0giJboaiwe2XkhGeCcvTupfjc8iS6H8bXQ7EzRF94GS
IvzUeESAiPDwM0JiX9YmNvwgNs07NOd9a3/kanmF83imVyIP68afyszk41rZ
q37rPocoN34rLDOjJkv+4uJLf0FvInVlaH8k73khu9Xahk7etJLwA0Ig8S2r
y0QzjB98YUz1qorT5b4FQ6AH9ihTcc5Nm+BaWu0BxaHh6bID+GVrTQ5b8XIO
MGriagDn9a8kbQnxdGJ8/F42S1JQ6pNUYM1D1t5z61NX24gog47GMRk7iWMU
fewtuB/92NVvEYSqTBbyWXQJZCydgBuOxlg9ImZ+A5HPymQM2vnAC4L48Yn8
Tnu8DLk/7QDkShE6mN6Wj4+tXfxIVcBMNHmVs5SiFybC2V4MP9vTU1jZiBHA
hD1uv3Qw8FRRXTRhIwyAWy2GG/OL20NJn29b6zOngidG5B0DewPJjt7Qmmnm
cxBm3zEuBU4ZMZVTtHf9EzmnPD36Od80I5KDNn2BWDAEu5NODIiQSvtamBOr
cWgKLLsPFQQeYg4DBAKVQ4CVRpi8+8e5LKovFCyvF/CJvhN6GVcTB54E0UQz
mxl6L7NjH0GyTEefxowRu7kMi9cFKRBkG6GI7fwZxkE4u3Uwfm/qjHH0w+CQ
vJ/BSa++1/hLEcD50+bL4NkuOF2erZ3bSW95jRq7TYYc328T/KvXY3qCKCPq
MDPRi0RVrgBXG+8+PQtk2kjQeu73TZg5SWkd1m9nlz0OYAftYnjhl4kDYrZ+
aMgnoMzuxXNJuqJ+05x3Y+mjrgW6wXLzbB6SQ31unA/9aAzpHYy8mnTwoq+O
a0+kziRuR8ryJHT0cpF+ZuRPAZYJwfZ6dCvc+8EYT+lKM9vW5AgfXwr4w2Xz
gFwLFXSkwIO2onGCT2PsRWsAyqNRUwIqcmkf/6Od1MwybApjSJcPkovvSD4m
pBW+hqGl7myyI3s0lvPw+Hri3xKl75Jch5t+3NuMfnHai2bvfmnt5X6a3KQo
6wk+W4jHSk7MpWkir/pOU5DVA31rgmd7cYDtRAwsMnxNY2A4Bff9ApFCnhJS
I0X943rFSQhmnUBqT/2N2A9bBawljd9wdZp63DHvp7NEl180Dr9nJimKXUaC
+QzFX3c2d9RU0Lzai8Pfr0mMUvD7zdzCzYwXSXYgM9l7Aw+p22PqMTZrFKkr
fuwDtdS0x5B5qEFPs9/xnTfXcyvAg8eKY0OC2jGIMsF9uXwcyWgpIWPDtB0x
Lc9MNVRsNlRIWlxqbGXb8EH4ZEowUmaWIMnhCJ8OE4UZctRGC+kIR907c6wR
HuX26MzZcaXkPqPUSJk63JviQNVr4mQ22fsrqx5ydrddT3BZ1+dQcqe+c7p5
wu7LeVvWomT+APT6zXlffGvCA/X/g5xwUBpIlqf7dNDuvl+m6IsJkN0tq24q
8JezOD1Z8UXuBMZelnO90QBWKtemzDUqPVpD4v7BeNOOK74Bpav6oqa1z1+6
2n5cODMCfLUdWlG4dflFlmPE/5aB8XqFXkfDqPQqeUGi35A5Nax8yCX6ZoG3
6cDTktsk+PlL4+73FZocI6z1dGHkSEPZG26Edk6UJZ5vxO6nGAwUO48UTYAX
Q3FgEpuNyflbFoepml6Ku9nSbOee9UFklT81X3zZiSkOiZLFEdLdFv1dKQ04
AzkqVZfdXoLSYS1hbtRe+DEuf/ZJyIhj6oyyrXLseeW97yakO+fEzMb5W1bD
oMZ7HA+p6A3OFq0zpsR7lAD3oKpDiUi+x/z3E3YtDIXHn1/rBvxdhI8oBFbl
clBagcYF2TKrRc47E+dUcpAVuImrkJxwu7mNxNv9njXKDwIjuHrn9W8cOnUS
yGYG4bdysEX7VNgPhFF7cHMGR1n8MpcmU85yty/KfJxp/naWRSeES/H9Ndul
WtZsykpl6neCrPaYn3KogbRqpWa7ZxD5MklWJ3oMtbYX49ho/o28ryUYcvHg
5g5DUu5cQN4ni+09RXN+Zrua7iPbEl5YY3RFxu8ule6h2nim/VyLwJGwCh3o
4rfm3/B7T1KU/wIeYVppYaWnZlzuPM/3uibzrWkfsp3InEY4x22RZimJjkO6
LWr+VF7W4CK8Jf59eNpqQQ6eTe2H8FxdHXV6UFhlK7n5M+a5ZrIEINABNg6N
oVYkocJIc92u4lrdrEef4v0wMmd++gDd+RllUVR65xMFRMzxCu+Xr73hO57N
TjMg+oyRIheCUvdUSXAGYHN/aZamhgCMT7zdEnZpYIfXTkt1wq7CtHIxPpU3
0lWwXlIb8CICHN/5C8sytWjBHkNOaRQHuYCV0njd6r5KUFUaFQFQjdfyNLP4
b8zZ0wLvlZw/n4/ljqZpBKyDS5XxqwKZIFUnopZs5BRAl7SC5UiuhVmZsO+N
hkk1NfAalmORFCaClAawqW09T0E3qWIpBUmZtU3KaPpK36h8JhMvXM5ijq0j
I0pziNxYCspB4qPQxC0EHrL3iFYlTdMz7P+F7zu3fJdiM3XsxVWZ9hZXDKiO
iZAh9BlwuqVdsVRLq0xnzhIZgbSz/n/2YUawWk6SoIchvXNjkcbxgKRMvxC2
2CCAdbksQZa6TcI4U6JhhR8jN1YW8hDfvEJ3e8fbAUtQvVK3ODWvaAJSitiD
XqJ2GlM0zYj5sPLQggm9WnXU/ROFC5Vixw5aw4YzfRynA0h1gSEvzqQzA8n3
uc+l4fwEJ5XteW6BfsgoykftOAXizxisR+YkJ6QM/fI4ix+9ZxsiBQONpG72
wW0bNVYZSWBhNaFON69mOJwgeFZWNt7nA9kRGFu9u23zPyxgdskJCm8cZtZv
vCCxuXLZa3AIuIHtKbbr3XhVSP4TI0Qx0238Zcd+OtLIfx1U5vqCzSsdVQF3
FpDMZpY7nIpB/4sfEHsymVFS8YNm4EYghVB80ELxWpSSqlA1TrjoQYKB5BED
DhMeb7VpNl6PQwwrRkaw5WPE+PAveIzZBUSlCWG5zcJXtH12ev3Csmm9Hnyp
Hfs9xkdc0B6T6W4yfB1GOItmbCTZ/OaZohV3QI5cHCiw9QMqh8o04C2gX3xr
tGwUJ6p4th3VBQaffCSW66VOWNsZjVZHMCbBMgvH86wu19II8JLcJCtzxU98
tmXNz/b9BjHtgb94+8O6Fa5FpA/n1Aos37iMOhndXE7UzTqZLDFSpCeXBuh6
+C6EB/tSISKHuFfla1SwqfsJsom3k7IftWZHt64wWTVssOvKxYixx/tp/MTd
h+oZepCCflQHvnowYl8ipVmZ9P9rU21fu5kQWQ6JM2Ie8i7rS7T4RlyMGhEN
Of+EGyIbrcvBEInHSci6ntBf2WAadlFPvefzbx7pq4hORUqCpgR+9xl4J3yZ
rs4yFFyILwyJYtiCUHTf3XSxfsSIS9iEdrsu3tJWOmCmkSR3Z6ny3UuI/i2D
I+XaVX9AxKLW9uIP7PbA/HRo2roVPW177XnDkEiBIfeUF1rVoEpruJiLR8ej
04AcbslgNF/VjLma2vgxXPXFMEVmmClpk/GheWo/WJYzTnaGscZl44w/4sE2
EzRtgV8Z+YT5Tu76vtQT3McsvOgmptOl8Pi4XjUawNaq6cMxLaEZsCvXI/bY
3wZ2uJi2ToAUxRb3XIJihCSonZaVFEawO9hrlB4/HNPwsqWhFzWxcU9SC6wE
+3qKSlFCHEwdlhOmmBkqcY6oG79zWQFuEg9SG1ZIDu/FQz36RJjeEOwpEdbi
nE7PapGk9yx+tUMNcvGArw01pK9d0cN0jJdCNaafn6cbMdRBrIqF9oWEO13F
U54BsYxFaz2hPzqNK1h7yaSlGvwJ0e2Vkx97cCIdjgkdw0YTbiYN9yEXt3/M
VyO/iZ6/iqZghowaflGZwhmA2YeGv4m/qNDIVWkydRxYdp7GAG+bxnnZm3X4
ht4D3eAbIqxuQOVQgrdLwOGaCBg34pAqUt4v47mgqFF08h0QO/gIRncEqJHj
EdPw19xvAyhVeH5RoN0IrYBmn30g6mrmVJDFYT2BIVjY8ojiQ2iXcyj//BuJ
s5DPXewwxZ6AM1Vt5CmH7vRWoSJ/Q0VsTOa7kEFk9cZ+U6QioRjVIUX8SkKJ
mUtUo1z8aFzww1ciQ7/InT6HXgRY81qXe/lrUxzUMqAKtDm0szNyDLfXG6wv
uRZGSTQYOrCl/qzJerf8PtcUPuxStgHlXAuovZQwT+EMAeGpv8VGUK6WUd2J
PCWqumuI3eXNEhXjqu10Xe7RI6z8qT/R3Kc4O4+zZM3BwI2XdFjrqeNyv0P6
tjeTRuYY57ioDsjMSsPeJp+gHRVz/CYq4JHlI11Ujulh1kM5q9ixf4h5V/vM
EMBxHTC9KJ1j112Mi/F1eEBgrChvRaky167rbsyzkNdB8BBJ/vP7mxoo6ARc
bUnbr0UGeGIVedTerCXkl71CA5Vam51VVrg8tWC5aZHxMwWeb7p8JP9DoFQi
YL7GuU2btUD8q1XgMzIJhdcT4ZLP+qlbgcUOEuPuP1gqe53ml6uypGKWZL/b
XNBy21tThGzCxj8J6+pMbJAcM8pP6qqhnnbQnsQhqsMy/7csNVioVO2M0fE4
8Gk7Z+hAl3EtBAaVMkWPCJtfKKCApY4fzCq8n2EqrOALVENim1H6p/FYUSz3
qNsPPwUQAQXvc1U01lNOM8m9JnHhxONzs5JqDcZvOLLS5o0G/exnWrA9KEGI
NJ+r9Jmb8uo8ZDaeCN3+v0mLGp7fYRIOQOpIrxiYQxl30xS8Igiqz6EOssju
Eb2xwJLYQzni7CJxDvPRWIMB+g8n6EZu1JYzQ2Eipctvo8Tit0QYgc9WbOqJ
gjkpavG90AzeUxxHO99ii1IbQIdpgrKV2oTD38wJLYKl0cEv9qnbnzWD+8Fa
qIJGi0mzVTZZp05UOVQT3rtoRndJmJ037O+SpLGJ9V4Tcg13HsiOE/zZfY/Z
K96kXTLWb/m/HD2A+/y3JtjGWC5b6rgfrtlj0PkdKGNrKRiyS5q4kAOgKHh0
5Qx2EpofxajHtaks8dCoYGo2MbPmrpT1vT8o4GRC3+oLIdUhhkRlk2GRjzo7
0ebmiGWIMWZkMtbM7f+yUyFf6L64tTvayRZb5wZkENVj8Hjr4CI6ZrtCWrzm
CGD3ko8Lrx1iP2KjnitMVhBuLR7qqr7JK+y9uPj6eLpyvHThVY3ulN4rzv/Y
OLKs9USgVwXHCG4VqlGDKCCaUeIyxcdwlz2YwybenVc1VvaLcvWeTIL+EFX6
eue+jPVKmHat6XRgt7+vL4vK7+uVBO/snXJ4Bj06l9QiJyj70Q1cQ8M5gW/U
Q0van2rZY38YFPrVwaN1reMbJxDzaEQnDAf69k1vigTBjql2PLdk76pCImuI
PjREfFX1hY4J84t3Rrs2ZdAy5r8vCcqC1j71+USV0klCAsMHNBdi0K1Ubjlq
3VfGb6botp7Uxr54KZtRp6YK1USEirYtInCf2YMoTxO8uqEr+W9emfQROtN0
QuhfzTpPF1JtS3+7mIOzjzOtQKU3OaQ8RIHJlBROlUGhVjWWjzPnjeUl9TDT
8o4HXKKNBD8TBD1rkntlYUYoCtwzGvyStv5lsY3X3ejKMW9GTKg711EwPkbi
G6VMNWKusVVrpmEvHRL7k7NJU1M102FXlFOvQsFCLbEFzaq4Z2x78OI9X4wi
EHdE4ToY/i0yZNhVOXasrlO6evhZOznBMzU6MgqgmJaQdpPdsbEUTuaqf77T
LdqFUeLIlpRkmt9ZWdTZRGgDt+Kv0iTuhVzFseV9GmWVYUTn5GU43mw7pMXJ
RCTz+acvW7QtB4Boj2cmCKvhrwCYVSnxWVNUxpGfLewBlmdAPeV3ieoSwyR8
L9JVGzVzPPhD1SM6ovfCirxymxtd8dLl3BrKF0Cw01Q5g1jzxrDsWRZaTKQ7
4XU580R0w808rzb+Xy4+UWF70OCzwd5265qdbNyqtHzotE/7popzdC1XiPvt
mG5yeU350DXUPvywD5Ts9Gts2B/pIwjOkIrasqnD+aos/LXY182AYXQE9zwv
0JTk3k1JZvFOxG1LLwLSaY2Clxn1ZIjqeWv4TxouPTx5xGgkGRUj513pYOry
H2xi7055GfopFafqjib01XBoTsYBTTvKMRDIN0TSsXo+LkPk+D5cQizEbSse
qbxRUV06k68YRpHS6x14iDF2MhWYR3L20DQy59ZUaRnSkqrOWjOQDMKUHePu
5erPeoDZazwX/fO6zhx9ngrpo4PSI7i8q7FbmQ5BZhQRMw/daWYtQwr04VHD
grL7GpF68mTwaJrkvwJUUVJ/91lerzUgk+u2HR2Po9GqBuvuqLpyyZCVcgtM
FswEfbFXHoDxmj/YoxSbY9uk0q9JHn14YLyuX5Y5BhZpj2uOqCKl8ol4cKfg
xqyF6qcdsHTZ0Z5PwtYZ/Uc7d7PqfobR3V5XAsIL6AiBNNNjP7NOLhDqPjUz
CVFL5r6dGzI00Kk6uGo6XMqJliJViudW7KmyTLP+OhPJqsCpsjOeu7YOlde9
GAjY9kyVWWQV8lB75v5BoDG2GSJknZhpD3fJZmpYkygx/bWQ52RVJda5hBeJ
PsOIQejjbG69oHWpeaU62rdlvetBhP3I5P2wdEiTrd4AVlHSg/jPSSq8UG4J
xCYCGzxIqCuW/XOgy41aVB9aYPTzJFh8cg08z8rTWElxOQSMgvdGlSoqT8iW
bxhW+SkqIB0KASYfgbin9ie8CBWMwg/7e7MO0cg7yqH2JVmzQ4w29hRtu5Kr
ConOuWvoMrbAgigRodhQkNkpxVAvZibd+JTUQ3IadoiVUMK60qVEIzS2bJt9
MdiIabep+2LUlGpIeUFcORkicSr0yfyDHVR9KPPYJM0YlsGe6V11jXpEP8hg
vZyh2hdKiKu9JKfK2aA0TI8+2d9BVvhhb8G6CvtN5BKG7Ss0GzinuJPYBsbg
QvF1YGcE8fPt02ftTOL/qCTKwful7O5KFhj4Kn6c9GJvgTe3Sg/IkD5UMo8w
GZVW+zNOFt+BIiD/tbP/uxayBlyg17uBfr86HH4UTbMfw9/VRfH++jBf/d23
aC/R3SI3js3L4TE9oK0XUsnMs9oAk4yHAk/z/OdjUMatMaEtwljy9BwLim2e
rbPi2dNKYJccOAK8dWOKsBNLmeajKOB9xaLS5wcTujOfyPdtr6u7vJlKJp4e
NP8RSKxdbstUUUbYhbwtq14RcodxRc+eeifo1NJ0vpCBZS7LZMsLGdl1toae
gdYkkNgf9z7vofv+c43EYDIwGhDufxq76t9iFmDccKVIwsJ+URLxcG06Eyns
H9inNu2o1gVuU1PPwo3eDnuYYJajZt03NyY+UBoTw48KWEAcJE3ZRDp24qow
gUPlZWHOHx0fAWfW9hoZK6QLTLI2u868/FYkskHEkACoF0yyl0xJj42v5C/K
Th5K/DL6bHdUAvhgZzY0JH8WNhQ1fC9TXI/n1cq7WqaSoIVWgb6h01tEe6DR
P6Hc3MQCIqknONK1kcw+Tc9c1cN/K/GWGSL9Lxlo9a2q71M/LO9STFKN/r1Z
2oNpmZpT36H0l9byGDYong54cToKtGfJ4I7Vk8REb/DcxwSgipAzAbxXgI6y
UcSgktQemBgFYaUS51Hd+pmgnimZ923xTU1WNrhfs7xEm0AAtam4ciD/EgT6
ITUP5JJKxV8TDDzV2F/NuP13OFsBAaTvhUZyzf5RveqPG7kTCxNU/IjkoLJx
8R368pvEvQht/0XyoLYAGRx224fkkqDSeUAZ7pKOZ83+5Jc6M6Eo/ivmKDds
29x7MAfFQdJD2CBk9YxoUafICM5/ECYD4R60TtEe5iAHekyXDL9/SkKz5KBB
VFHAu353CcQW/L2PXRiNioQGPfagv/SDWurlgjWJSvz6rHqhs0gkhAZI+kA5
SDBeW7iDt5XsP5Oa0R0UZwEzsS2WGkXBOQjpb2oCqhPqxbDNgc7Hrnk95kLT
Lj5nauxVf0/RfZYimS9WFTezFhAfth4/x4e3nsMrodZagFDR/v3CeZWP9hxe
rSKD6Q4dDuomA+GTCHCbhoSME+Xc+QAiZJFuc8pcIA8uKgFVImOffZudfafj
N7yZ3PT9SjNihyFUB+vG5t2zhxlV1u3GQ/NOZxDKttQxX97NWybXKgZ3jtvT
28BCqkkcaJep+RDi5Mpdu2/sexbJcF4g/b8fccmNWW9Ul+lW/Jc89Gm1b4Af
bqNR0oQPpaYWcnu2abwTkUCSK9U5xi/Ftq7/ztOJHjP500mg+9cq8u9fz06G
jgN2L+xiRd6Bt2QWpQSRAeK72v04nl02Z0i06yPZVsb/mAgulO8ZYdLeuOdd
QmnIG4MnvnmFNfp3JWxyoUpVcAqCdKBs6b/4XeykIH6KeSlkLiZztsbI4HZU
Km+txh6VcDsBSjLIWQ/nGtG+rjDSu5yXFp6ipNwY5QZpvh/2eExexaVeDDed
7++Wnixv928RYueY5btu9mBBvLdC0VIKAm3W1cXksB9f8gsfHUwGBbBMBB7x
TbgByusVASchqD6uNiwgjAM92zf7oQhG6pf5ksVi+1V3NUH1WlW68moSGwId
8OuIQPzjhBk/DN6l6nOZN8GPv5IaYUDZsWi5aIDwe+nnkyK00gDpSxdCXfVk
AOo/z7SXYRkJ0Igr4Ok8zjHQsAkOqS3rbyLmlJf6culX8U2vMQaByIiwH6JY
JGzxUk5swPfbRiD+YB/GLagx9mt+ewQh1RAhy0Kwu16hsIFhcKAYOzGa/ViU
Pp5C5L2lKA9Lk7cSy3WFSZxpZRMCurWVQlnajVTqHn9bJQTyVl/hF1ZENfBS
a9KkLtuqWlUmXZhb1SL6j22EG+ZzLctKAIJTwsSIXRMbTIxGluKVP5nCUTvx
qGZiH/xKbGY03LJ8roN7NmDaQ9nm4lg8HF3PL80cqamoTyKBdDrRV15Has0c
q76QaCs/oRncHM9al/74CnyXdxVc9b2/7/H/6hJdR4fEi1bCPITx2ovZhAr5
ssLxj+BlH4F9pu2LY4I8fOU7nDWqEr/hxnhH7f7X4j90ZTOYCAoGW1cmmsqt
kD49dlRMk0L/U4j55ybtr29k9EQG6RJbQCTWxU48ETZNzPjw+lI44Hg6FUmW
BgxP28VJruyHJfAJmC62BpUIlQJ0RL7mxEHFb8KXb8DL3YcZcD9UIDKM9xZq
NR5V+KYIToHilvvN9oiXNbdmBY7BXskeNjAdn6Om19ZCNGUwMjQxar8ndH1+
Qzndx1eQ1FPgXcKTnEkihYVfY+mcKshVQynHB0IILitjA6ktetxrULSzLtwS
MY6VztInPHQZzP5GxQw4rkuibduCCWvsLhaIjbQKucDOY1SQxufwu7v+XEXs
oM2JQDyngdDJ43SIVZKesIpZZtu5Dzx3JyZadQfs52Dwh9OmgI7/UGYqGuff
vB0yEaZ9Xo9ZAIsdVJ7Ur4vmcgYq+AcjCU2ZmeEYSAEXtzObj0c9lzA+a1MM
UZa3nFjelloSW12LT2CytgHBAxEL6nZuDypNPi/S+1tH3uNZgkJblQ+FWef2
cMU8WRKcm01qaY9NFiEeaKO0q2nTk/0gBrA1vMEF1ZENjKqnpbbzsi7RCVtZ
bEzgLMrPKuJ3Scr5ESbS1AiLUbpqQpC1FykUuNQFHOhfORda+VAOHAFJjgfN
jbzeIXJdOFHGykfW7xacie11z4lV4hV+OeeXWHyKKBvlyMS0QG2IKuLDccga
4XoMzMJbwzDlCpFNlUo0hYqDnwqDSHiNfyCSJ804aawSA59B3kb0fNfwt8Cq
nINnqFbyxs/ZY9ESNsGu3qxSrXsnPNwoasVMvYvQuTXrhMALcI+7SkwuotiZ
jfNnrNL3lCP4AEQMA72ANQ/Nd/5TL/X2+bkBzFfGHgHJiVGyt8cOe3w+xn/r
r6ek54+QsbbN5QuufBH/60c53Dobzgvvo6DGb2Er6/icprDcMAiUHkYB0Dwe
M7ASs2N+6ZoNWYkngUbRatpQYGYLLkbqSeSATkzZi8e9ZSVQWVlFiaOppX4t
hD+Cs1LE7Ms9WtiiXGVZfTiYxS3Tm6oOI4cjouYRvBwqvwpZ/hTQYaqCPS1W
8dvgCqBZCamYjgvBxTn4YooFeUiMRrQTZSuwwS7C+84uQlGO8qECxs/YaIU5
uzUDqSdUWJWbD0wcPBP3kMbvE/J01bN4dvKVLol8jAOJjt5FskfdTlmWBTUB
TWRWZ3MBXGzssopNOWgot08+Y6sJf4htOwCT5i9Glgy3oD1nyl5PuZwxrWpj
7CiWTB8yiF3qNPyLkM6G8UrdIELP3X2pB3HNczvV0/037L6OMe/1ssb3gB02
O90aeQlfbmSPMWmPdDMsqlbgpZelNwfbWTiXyVJdjOEbCCkDIcA7laUJKTda
62/z3Z5WvwWGcE6rRiXj/7yZjqJZpGzCvEAG+Eey2DKxiTnYpZGN1j99Z0jX
gNdl3bAdyhCxk72thfjcZXbWeKkGt0lSo6hcXzdo0LoK2RF+o2u7/7bGQKL6
4zB74436dHWRzmfgW6zIoAGxbXTTEJx+l37DE0p0Mdz5Q9pr3Z1Z+723Xf98
K5qT3ch7Y72wILvQt48iy2u8h7iCtpSaCvu9KzyceJ15mNyYzg9TDVj3KLP4
A3o6VpmSJf8utaSCSREa/nmLDiqF8DpdlenPv342fh27zfpkAdnR+oQ31t22
cWK1igfscLfNEh8xhQfxhzlnpSshK46+f5OAZ5O3AZc35V251TXkZFsup+rl
pARTh4aNFpK1UGx2aeh004P4AnpPj+0nwy2E5vFHF1zDUhXZgD6Pp4O422T8
LluqDwa8QY1F+LFdAqYLRA0DKkH8DCHhrURcijOV3TE0KC66UeTmrhjtNN7N
98Ubt/j9sMjjVH+EnFhBGmPG3ZaWn0NXKyuJrCP4MwsNwSx0y929x6mjLVEA
tq9ogMKscwxxF8inx2NMhGCYH6Wn3r6EIaN35LZg9eTm7bvmAbAoC+xeapZf
nQLKNKJ+E0E0AgO1vHWt2NQf2HnPObzy4W5F1DgpCgTlF4L3I+0Opaz9D928
M//GRCKbsGS2QJ8Ja0P5dKnpsyNK9YXUkVju3FsB4B5f1gk7kofNCMrB7dSZ
nDO5aIaFnFxQFkx4A8SAc6Ye/M2dfU7OBhytRaRVzh6CV0KJiFv0Oicm6Y0g
MVkBYJdc+PBydcKh87JH9K0m3PRw8kJBSZCvYq7N/2gHYoZdc8nskRvrKxZF
i5ckSVKk4PhxZ32QWFGGYggeUMzGVQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQozonIdtulbSjKTkzRhQnu198D6t9bzEM+6lgdYmJYhG27PZS/y+HSM5TaQS9UIQ4O6K/vDhayrCGxegiB+2yqKNx5EciYBPzxmlwLZwmOFhSYYzLi2JLIHoLnC2LYGXsVprViD93RBY1juIVXfOsKDEAGIcyP1ySRFrVpvMBagP+ZSHbnoWOn1n5ywxhVoFrvkop8Xnchm46EYs+oiAmKj9PwpxaZrYsPoPbUhUAHGx4j2nflAu/99KaP3AMnzD72EiCwKLCu3BgveWby3Yt+W06z7ORq518CNjdosyFc20fGH70Z/B0WRoxVflB9QXzQVxs6cX8Giog24ljPW92p+KfcM/5qpYQJlCguUjiFmZLv6Znh3sJnCJmlM6SXdl7BaZ/GEQyg5Ywlxvp9fYstBwsIwvJW9LCYlTR/00MV6Y3lT25NpK6jPN5QkLBv+pDaM+xJbIs3JBVOZxTZh04liZaOAOzpW8433mDMMwlM5+l5DcrHFzCc9q3QBlM5v1bHKSA9CRl5JusSb9gVashgHCWL9v/mvGoD3x3f/syZ2Bl9OjJNtMUt+7mM4ybPC4Bx8gCx8Dk1zR0pmnw1xDxs1YWklDt4go9JUeUIykzTiWjuGLgJyNIbyS3m5MjaC7/5YwFPnuR4cH4SSPEoLi1al2E0Zxl3auluP3QhGRcU0tJEoDBxA15zkpP/a8w/ysLYObDurEQCRp8huMYn1tr3MBWvLFQ85b6s7XNmLcMcGpEsWu38CQMMtrpWLYy8Wr9XUkbud7mb2ohDeu/vTTCLg1"
`endif