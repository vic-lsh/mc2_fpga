// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gixnoT0P6k5ZM6OU3YknHS6Gk4+p5W7wlq89oIfqZysccQtn5atSUTXpak9h
XcYAxMEJtOFn3/6SO6Lbuxq9ihCzAH0oynQnHDFfZN1sjI+cugGFeM5GZNXe
++Pi0M16HPOXQiAKGTZBHB+ubejwi46IttuJzulzGgjcC4Xf3cJHzVYA5qzI
GqAIq0B4nTmTNvt/QvUTeHijQ2YXntR0JFFeIoxW478ugJtBSG8xmTJK2osz
aVkdMhOAxKNS9THlQVUbl/+FQjbfMYm2lPzbhkfhTxzepjI8TqDhj7nM6+li
8fK9CDOrK8+YlxwEEGCQ4WFUiHt2VOpeW1c77vSGhA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pIQSnzXhMVc8rxKwh0ACUsaDgr+bx2aKtOTCin2rEkQs1dHFQvhqXSDyWAld
Rh4wCYGLhAQ0J/CHDnggPSwnYMsJB5whwnMpScPBWMe648uZMuCODaZhRHz5
iVTHrVxheJVt7GyFb8nAaNZDIJSf4PfN2iNSH/RXcjXiPgadYYreVpaLwOPi
plmgeSflgMZan5REMTElKMqousDPSM3moin+9q8tSTLl8ac00z1LAOlNSb0k
IYWaXbpM0NMVPNpRuWQVPat6f/F/cg3yJophadD0trGsFfWkFypgk6/UC5PT
LObcxTlt/w64YvAYXZCOM4k1L1O/QRFDCZPJdnmqvg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
j/SHYLOW4Wb/Ru3LQOk080+hMeQDSXaTTW8pC30u/CAHMbjweYRxcLiRh824
DnerHccdERrVWg2bUGj1DKntLjYCRMOpXXLBLA9O9SCbaECT+g6/HRVkkGtr
ezHKXMfyQ/nvo/w4dXzop5ptYKpfpfsOpYnzrddaJBFrG0o7mqzBMYkW1t59
JyVq+N83bIisqztHp98g8xoLEZD1OaImTPJB8CXwLTNB83ofMKzrXtmDjVN/
deIKDRekB/RIwoI7DUMLH7Gt+0KVXgBXo8JhMSHvh4fpF7Zu9yU9z2sBqIjI
NN+gGjIzGn0+oCSDDzMfBKuZZLnR40LXawpT3XxNaA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
X7yBE064dwn0lKYiSeW8dItCHlI1GyObuc5iTlBe2CnyoGD/EZfNelIfbxkG
uHbm5dd1I6TBhrTiEj2I5UvDptNePMf8QPZjAPcivWaQ0IKrnh1qgCWaCIsf
ioGkq8Oxpx8V57JgxMv4Pm+MMVeGHhjUw7+dIOScQfy852eTYeZJZQmaeNJ3
2A7eNWSCY10UFEoWozFQCb81QToK0aYXTfH+ihzcWDG4MWuyNR+Lz6ErVh/P
5tF2hXqe8F0o97BJ/cnSRRUUX9Bv2RJ6NvTY+v+Rw/+4HmNjMTlOY0esMm0n
CRuSR6nz5tMMdaSdOYttoXu1fj87LlzsOxr1IkU7DA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Fg3v8S2TyJbp8UfwDg8O69PknIBHldKXkkJCFC9pONNWsmjbCn6z7xS6NPBT
y4fEaVCXuZe8p4VpCDIRQIMgB+577j80xIRg8d+4hMtNIdDyi3wLVWy12/2e
ZnHmCta0jktkkhypFtFMWRGnTF3wY9hiW8NSM8ZVHD/Y2RQr7og=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
svvi0MeJV5TOhxTcw/j6V63qP7cjAqlSe2XUjIh7INuuyB3fMMivzzqeurcJ
kPsSMCd6IajWJ/Pr+7NtopoPUMHcSqUh0ej1Sqb5vn2q5XaOgtJX4+MLKob8
tWhjStH3MmhsfXE+8J00RKAXcBNIX7C8GBCMvjh6zqH9h5WfEKf/UV++Fof0
PKIqDrVRS6pCw269NKpkMuzXLYknVe52/aIkv23V7nkFACosJmgFwr8pTgPt
KmuMDNH5tC9WZb6YvDzySfPCFOrYBbtSIwxBGoIF3hUD/SlZLjPsfHVPHpNX
R1Eid95ac8mZmnRPEDv7PclhxdbpE4eZz/eMMVUTgyWjNg3xWqDZXi3LVwHM
YGlCicrxNQQcyQU1Tu8ulbqUbq3FJ3VqxQsNx0iOL8fgitYz3kZfA16oRnfx
UTjkuN9oKjd3nRzTxEk7PdIq29sE0PApQSU2NVLoukzB9pK9W0oTsVJr+/yZ
cBZPq4z3JScS4A70dH+yATgDJQYgKFPg


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lWy8e6niGsieVPVHTEzplSy+Q1ltFjkou1TCWi/+cZ0dKEtH3F1s1ZXcrTk6
FH9hjDWr/5JFuvTqybcH57W+ZASi8G5vBcLIL2rCsybhZUlbwSilvPRm8V5Q
k+yEPkB/WEY6xEBCpVkVLQwb6D206I+vRE6Py5gnapowM6fpp/4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gBFba2pTQgutEXLaN6erAosCPR3WMEp6myybcId9UFGPVhLlj2Fb31fVLg+O
yihHaTReomS5OC24WEywvMOIeqGeSZVWb+achoeWnh+agnHmFyqMu/0XbbBw
iGZKCztIl19CqeEXNi5OUedftru+0NSwhYVQ4xFMeIKPbIVhF0o=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1456)
`pragma protect data_block
0UivgcW7+WdfMtK0kMUxcBQ7lRRnBVPovRntSUA9g0azWOl/tv+3w1jtRIXl
N/zdWxKKkx8t3JO5G0cbNanZ3doxbUcx9+RKO80/U2iplepdCEi36oBH6pFN
+H1bzS6PIh3fRFFYvNJXk2v3cQoAJ2BixuoiOL7wQO3jmke0fHnlJxgc5SeB
nJLcx5jOBGF7nM8dj2W9Y/WpLWtiqZNtSqwm0I1KXUciWswWXLw9Md1C/G1Q
kx9LWRBf3rUkhFTGCQmuN6W891EPpZlzYBK/x3+DW7RMkyXLJq39xMGaZaic
TUY4qlbeAhyw4wHNtg2B8jZSlQdjYYPBnXPeUaLiO/o5F3yIwAXPKDSx7IOG
kghA4pppu3ygn3JzOFlFtq1IxaoVlNZzE2brvQq8TkpQGxokuObFaSjUB2Zy
0vXwff3i2D+qdvBHFz+Byzb/xY60QkH7e5k8DV8bD0nfICfR42cps5Fp5iRo
M5WOA1NnJth+yl+7Di3j9ROWJd7rkN4Gsh2LTxXuLvDpFumCM1WnAIeC6zFW
+NI+ScNr9WeckE468saD+cxGik6d277btQrCFcKb/bNgrQTasUcmhAJp62Fl
AbSYCLWHxwqDAmiR3pllAz2Rze6bb6DdnOEyPsQ+cZiuRAXSglZZiCTczguZ
gRY+hPWpwkO6wJHqGrLY3NWUkSIccQcmT2YnU/en0DdhIO2LjmnzUARV5sMZ
esBW78CAh1XfzCtavLu+kpUrh9bfqGGoDclzXaDarPBXwu/jeqD/Lv9lRA87
toK6YkIsrOFxQGUQXGRervxD6gYn44DJhjQW4VVaNQToYdoDYIgqOBbguBJs
W4oPNS1A1ExPHbrPrS0NTZMAo2U4xauPWT5g13K5m0kXpOj+1BSrg1Czi1si
7ujvPnx9sB4aR7PFGhjO7DsA/IQ/TjfCrAGB1YwPi/z4+IHNtoQqyrRnNl6R
xjf5WLugrLd5YRUpzIAJDvNScF+n2r/K/HnBzHFDaHmHpmigR7edX+iyGuGW
GfdUidJ6fUQc0ZyDS3RHL2NMbIvLBavUS81zkqkGe627kVZHLrLlyeKiUy7h
JeNi/2urGEhocFmyG4bQJBdEBiyiQDyRmbzzSkZTbooX4DEvHyYTphNw7Nfv
y6sNOsYT0J5qb+IPPGEWS+dZCKoj0lLm6/DxfpR9GwxeEKL5DrwXrlT+9DNN
P7/Mz+HY3M/iDeYGOMktxfi0HCjh4YGAPiGrAoNhAlZ6Aelb2yMs8q7jssLu
2POHJhZO2VfUTXFPUtcnWu2QSlDExPC6wSYMGdQJCRh1aFmwozJY2G43TbzU
NoOSrY0uL5NcDuobjN9Ow2iVVNVwOvcyBS/H4VnbN14OFhCu2Sp0Q5foI23W
YjG1Azx4GKF9kZLf5OWr6k+3Wa5M2kuLt0qky04gHO3q5SBrbow84sA4WMNu
ouQdXsLq+8rNmTbt1qCxgiDpqYBUBfnhIAb1cN5yQWab24qscXhjKt2m/eNi
zEiHeUDqhxeU/si18IlLYd4HZ4428VX1VRHzaWpulb47yKjLpmeMY46Fa/72
ETSO7jMM4bSdgbJRVM6lRHhmrTycnUwnfpP9iGEbIZsbYvhCUGJV1FTRQuD6
R0d62u8oXWijYuuZpqhZwl91VDbb1HF5mkll9a7FjLQT3Mr9Cg4GAZU6mH6c
c6FzGP1cICbdcykHKRnfm9yPjlVT6pfKa5uD2QKkD+cvr+cLIQ4x9XcSrqcP
VmNFIQDG8QBCzWd8fcpKDLPF7WLJk0SvaVGkEn7DR4ZqGJ6gl3fqMqo84NiX
/+R8x9dtmc8ggkSEPHpovdkuiGubTIXkaG+416jgDCiOyWa4uAZadVeQoXRn
to4DlM1AL6dESvHXJeZu3NoGjueyg/VxgCIWnEwPAMftbLHpmyOrLWYMBm2w
plgv07o+TB5+mw7VWE/dMA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqc188zF0mhEAwzxJcJ7cDo59ENUMtTPfkiMKPCJDiQPPzT3MAA3vEkHDXbGiCWtuzlNVwrtJOatRA/CInXFr1EEckWfLnjOW9voxjRj+fFPXnZp3QfQNWoYADlf9F7X+mC6LstkoGpOb+hqka2t8YOoxggOI8kU8s3rBE6HmrSBAl6brAve+6e+DWYSZttdkQaJUYTQfvk3eeyH2OSdSUOUBeg+gG5GhWwPI6qdSzc+GBplEXttZe7GOsi7AlL4jK1Gx/zTJw8+UDzowyRRWhp64ex8mPIu+YuTipF+ACrjTwka/DEW6l+JuyEg6qnw0dTuBBYfNuHb2kv6jwQRsfGfln/Ss59VnD5QCngXHZFkUw2e1BORLuL6/Qz13APBXMDbUXLG0Jy140FXsBeI6W6otJW7uXLLVvtbkLc7WTG5Lv8LGT/HNHwSO0S9+G7V0AYIHNgiDY44UEikqgJrWdxcfBq3OKG/JTqONgRosTwwHWCs3nbF2ComzcAR83oby/XZ31PxI+Zz42JXNNJa9zyffnNXYHmQkJU7h9QS92s/bd8D03xQgie2tuFNfaV7MDVaVzkzX0zFskfpVZ5HGI+HNDXaQLm9hEt6g+4LWZ4OpG4gvaedT8tPSaU1GkDswHyKgH0GmDJMdIIKVAOe67IDjw7F2+sqtjojNq7pwet0R0pezf8caQ8uy/rZdyVbeoUltbEf4TQ6k8Ea/TJs4kDAlvM2kzgRXFH/7prtuJr75B121EQ0kVrRfDO0WB876vAGUX0PdpZru95B6LkythLR"
`endif