// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ywshV51xz4uJxB/HlcC5ejXZphoqrgcB73lOqKLEH6ckaAGeML3zxIRNDRzU
BIRzTwMLJC6DbPs+4N/WH1g+z0aZFJ5J7U8FV64l4SbVq594Q+sLJOQhpLgP
rMeTiNdpyIXufOQz0VBxGr7gUktivqUgPaUT393DlH5/4IA9narATp77hPiF
bf2j6mKhHvHO5GTxGFned8TdizcQuz9qGRU1X+/zOaqHQxARS+Siv55Bqa51
3DhmQWZP+TkjKNfq2ilMCZB0KCxmRPLNSdXa6yy5AnFfB36MpFPgweE9m2jp
keQr6vHiGVOZAyXsbnwP3HF8NvUT3WVPB+6GT2mrWQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Rvyxi4hWXCLkQRMzEQuZJuydwutrkDX7f+78mxX8CQSWj2FkDH2dR6XbhJU7
yOzKtmpnEIp3iXH6OLQPqe98QOjCfncyLYRCC4gkwG75EwvBDQys4iynbjD4
yBgSOqGowdDEX4PWnmCF3He4vY8Tcoje5kjGTpcff7iINzh/6xPx/wOkBylT
234sIiO58+E1z4jddcRYdA1WOFd3f0RiJ1N9GOsEZJF9oF6RtV0CRhSaOc7O
zn34ep4hd6ytafF+6hNEEL1iDd2y4d7gxhT6rN5JgRitjntjo4BvfqkazLNY
2pIGuJEYNSUxy/6Wm9kMVUBFeyDR0jS4yQh9ePaHlA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aj3xSBi+KXaE4rT+s4SJs5Qjh8p+JsXdR4W0XSrEhQEi47GgO4Za00YlCzQK
fiPYOAqeW69rVcKEX36dBz6GivzcVj7mIC20CLEuwrtb/JKb7pZX/i9Yvy3N
ZmLkVFXcvNCdQuHCmRWew6+ysPB3b3pxmzALp0QeJHPCoG3f6LrKmlhhHRtk
6ARYac76ZP0VpOq+qu3efHaFPwUmoh3EbQBGAzJUBCTgmGhmIF3wBRepn8Le
DYVDBKv5R6OSmzAHCUOvtQHy3jy2+Z+bObx2176iZgrr8SoDO3nrdP7iSR5V
6qu/tXRl4nwG86N9D1Y994YmoImVGyhKgZzxxwXdkQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WLI+RytJCNpwsY2ujPgFTUwFGL4V6G9mF+iEje5YpClacYl23VEaTckgIFOx
h7A2pnssEuqf6DUp2ON6kJI5+/fZVIlCG1O1Oard6QqXv5gw0nW5p+JQ+Q01
2R6UoKqBmIHcu48rf3UiB6tUCaO5JzDzmlKSEcakShwPiQOhQWxGXz5O8vFo
iZuLBjZSptQEPMKi0uF8n/gm8yT6t4oklVJRYeJcnYzGiOVEIaDCGE9TBBBx
xFpJ+iN7wxLNqPrnpdjy1aV+e4q+I46nbptx7z9DGj9VVtjH6ZrQnIFN5J6M
Hq4exRQ531yim5nfPDpARrmc++MH74L5TW3uc2BdoA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FA7yIrUF+cNvwBgUGWyLDd9xzpCIUxLfUY3N/XbGrQzOr4UkeFDtro4PaRKG
Md5RP7k5o5+kdsQtbDi2ci3uJdVAI8H6ed4EQb7P2Ws0URRDwQO/x619Jk2L
4kzzdu7GIYJU1JMiD+0LCzOvx8bSBpTwar+wX3R/5nBjNQ9f2gA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
VOPv1sVcWX+p+S4wRthTMB8zD5LWQb3T4fUGM6ZGWdkVj8cdDeL9z/beCDe+
5oeXrk1f5tYZ1ADxnRzJf3Pz8GgxXVhgwtKbdNpD9r+7pgeDhoiiVu+TlC/z
Wkhbr5GmZDYWUfRVxUmB081L40xXZMe4g2t29RUj/F+B4qzFWBKDGtZBI5ty
9JVr9pgRvBhj8W7aan0w6pprIe/ZAAMOpXGBCVQOd3Nsnxc3ljQsKN4mLRIY
9OBzvFq0FR8EdYqSv8C+L/TT7rHDEP5mjFRyxmNT7sA2BkGOpKU7ITgRB+3y
DBNdAGQM1Qh5TTt4z/uaEehEbqzvBLXXg/krJnP4qrAyrtkXeurElLrWeFBp
lWVkwVheHsL3tgLo7PI1+Sx1GWuENvEo7s/0yf+BSF2fvuMg9xk9dlfaIuWJ
ovYfYmL6//ocuF8GeJecFTB4iFc598/asC8Umn5/25dPP9LNKHv6I6220wGf
/lBbDhqp4vVfYo2IT+5fiD2Qwk6QqMkR


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jJq8qqiNFT0UKY0pd1JMHm0Vl01Rfzs8FyxVm5HnakKCpCMDuPUCUK0lqcsA
QAW8NsQIQLxlv/5/UoVWrBq5vxjiZP9V4Hnb6tn1u1/S4TK3mStT0eR7k4EA
MwxMWR4PrkNi7gRFzdfjypUG87k+CMm2XLvUrG/+DBUxFy+LBUc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rL4I/GeUv1pTDJLVQyNb4DC5oFcdsDe1yUKlXlVoElhXNHsqKnsl9vdR/w92
TouhLUp6HolAStwn3nkigt0c4sQelPwvEWKul36RVITyaKgK+ndN13jxrNvk
WelSz6d78azw+sle4YrfK8cyhaUQTELYvNlGTgj85C1eKr78wrE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7376)
`pragma protect data_block
lvWiEUBWFyLLLCZqWLEmvwOZbYlfNrgVkN+ota5O1iQZ6CER75aMdXtD8giS
TD4diAOFrJCS+jL6h/PehspFQv2c9vR88dTRw7veNe5FQuVu3d4ykCnt+Xkj
42oFfVejl9HUCd0OFM9cNOe4hltYRiw045mGLsBo84W7blz1RSDC9EXf/jnj
z9Gn6+G2SKtLj1pnsUUBEFTaotMV7bzROVQshnLEks0YnZCGKnoXDssqjOuw
H9hvb/ha8siFZgD2LwXoxzK5AZ9xhKhRcb3pcUpo9xhaN/hvd5Gvr7lL2LA8
jltNCjDqWKASvw1ivL/NvLvElXxkFl99hqGqyf5n94CTMKRoJIxsXc5Xd+NT
Eoa/nMGZNYqaFG9v/JR+7f3o/rq3o/KuHZ80TWKX1Cv+Tx69F0gyX60pMPgi
GmeamnzD3w7JtyHu3tyHvb1MEjoPGdQVD4R6ul6u/k4VOCGP1z47KOMbMnX/
sNYYLKgltIWhoixVr7HXH0SOV7zX0i8B8rqN+UcoeUOo4NXClKf5a9Db6JYW
k9TaFjhuqn2uZRiEDcDK0V1XMfCvIBN0lTuIDyT79VvyY9Nd1cjLfZhiydLH
zXxi3SjNfIGfEkC8ZEn78Aif4dEwCNQYAjexltflyewycmdqH3+x6RYjkmoB
TpFi52ukrbePZZgFdybf/VJED9i7Wy3uh2waaCwWdTr3WVWT9enb0xyUnHZK
VD4ITksagIFMJ0fVFewrXcX3R2LRKRgma+RPZHeD0S/VVkka84/Ev89oLKwq
kfRNVzWmJNuVQgcMpX9VoXAKUD+SUjatkWnBixFK8K+VBmeCbhTeJY33Zl0f
R0we8TkVE4TvAUgQRTSFBWWxCV+CClnHoIJ3lhVFZ6bIX1fb4okkNKIXieak
tzVODRatYdo7wK0XfgnCCyafz9YF6zUuCs1qytrLl8XA32f7IBsD72KnQYp+
ReHtV3LQlZfDWPyz8FYY6IqtFzM+TD93pgqOqkn3LeZCqnQAm9l/8qtEItfP
VGeIfIC0dpXBFVjVBg+w13QDXVhh3z5T+sq1r9CurZYgCftkQQtg7yjOQD+g
8qafYziZlz6H6h/85cH88UWuIVuDpiaQYIN4f1G9ZUv1Lhlp4fukqxJHWuNG
8xFldBH+uWegctivgGXqgJ6WfvNQqirT+rH1xNZyaNnJeUcns9uit7wj+2VL
w5myMPRWxGZD0QUQS6GLlYyWJJsNJ0gKCK4iAOYWIF8qH7zBOO/XSFnXRL6l
hmLJjXZk8uDk2sQOgjU4KREc3F+XaDmBK7kXyM8Mz9jt1qVOf/NaLZFU20Dn
G+wC94c5hO06/CbETcu4rFBSIBSKoOXel3IlOWrMkBmx07p+c/hypXsUwr3R
YHsg9lJHKd4JH4OtBMiOtQrMX+Ld1h6ItjX4bOrfSLycAxG5beuIGZ5hXNZe
FhCEb1aKpakP2fvh2/MMLf47LbBtzZuZDiqwsjUaZQvgfioEuP7Nh47neXRl
DAcd8lbgmETsKrS4Fk1ZgB4KTenLhOJ0Djixz2iONpqOGzVXOIbjR34z5lP7
oFoWwWtJt9SjlbaHbLhrhMneiMtd2bx9H/1W839k7B2atRprKyxYZEU8sMhh
TlxwtkWUh+XZteM5xd4XhBJwlY9njjuQkHBcHSYxxavpC8y89BJGvYubL4rp
gsNZhuwyjLBSeyzZuiDLQPZl9FazHcYmEIFbNNCDDAjDZpTBqSq8DcEE3o1f
sUJzP6mldAJ33RYVxyh7f6q+iVL5UAFv6fGTZLbfOwpcWWC7oSrhv0U9nYq1
qQdHX/Bg3UxhnRqq2Gi6hBd1aORJOuGZTPl2PSow8WruzlrI88rzNrTIfNQ5
0oKubCIX0oxFXQ+n06oCkssnDYXjGnqiX8beL4okM5rULwMM2bR0Zc1X0Z/I
BYyXT/2wSd6EetajqLAoeF2Qb6kyQ3obCR8LuklNGU2FVaXsid9KCM7XjxRD
5SXE/ydIN2CAWJeXyucYGNFQYdLGjcMWbUiwHFUtZoLTjulU1sgSBtVKZhgg
9O4BaMG3FVbqNTg+GpbRU6woVfs5AVbrbBp2aLeg1G/GIij5S3xeL/Pf0AmF
RFBevX8YRKrueK3WHauRw+xBA97v78NPAFDliPEdkcTg81VsAx61VDBGaTAY
QPneuVbrt2Vas8Bo6pztcsg1yB35Q5BqSrGCie0O5TWw35XQaiPeC3PZCfwX
fop4Y7FPbU2EB9/uYaXV8/9lo2qEjXhQTSmKLgkhwGYcIVOmw4kr8WZprJfh
tTdFLFa8XDVi/FXqekjnE4AlBA1NdWSRSw/NVpG85cqwA3xR73nYDmxsXGc7
EyWMwlQk4503QofHyhSRcTrvDLQPKU+qxWCVLNwz8kcKs3HXPzaQWGram3E1
OaSRNH5vXd/YilT0Efapv5LQqPnrvbfYxpVA6nAfhSTCvpyqhCbEu37MwNVb
WJMAJRXGPF9e0rI5B37Pv1WZmhIY1m6hv9lvuuimeo2ZQp+zSuecs2W3zYJZ
r7vCry7mjXW4u0oceEQDYO7ypZyZXuVY+zz3rqDJ4tsHpcxyX9579uCg0Lle
TFHdM9EB3EXLvcR2BZU84Tb2/ol1GpInP4JXpyd67D0TWoIjUZYRuwjMPlx1
bFZGfdVfvPtlk/VdR7AG0F8iso+rsehgkOUK4LBSjf4BgmWyuG7dli8O+svk
VIYKtmxG2O0cJuskANN41d3X7efEGM7jqg96tL5rsOPYPyr4f6a5Dp8pWdtF
ZUs/QemjEfATXMTxrgoJidb+4R4SJWwUYz0hQxfn3fAILKkDGEeUpgaN82UT
w7breMQQo6burRYXK5UQr6yeR4VbgjBCN7sw7riUzNCclJPs4yqYImbGf9/C
RFBXjJZVHuZgHL9QyCPOZ7p1ua273OcU9mAilVs8PEoECNYjR7n/X8og8Vt7
7iSTreTgfzPCpqP8vufJfOq7fMOzNmkze7A/BrYutQaIY/Ru+YqxXyNu5e9j
ZPDXd5oTkeRznEgdzA21CA810qCr6O1yEJb6+2ZLDdCcUZcXpiqUyEDAvlts
HF7NY7uacAXJ6lxK0oG2UA680rrCqRzXTMgJ+TyJBnHb3DvdHiqP3wsAGUpI
d920fQq0VpUAhjZRwBfNnRHwAGc6BBzpDl2CYStye1SfB6MW2sVtzov95DkB
Qk8YGapzRWcGItjnUDFlb2l5/t0JfHLaEYkP2BzyPl/1nihtF8UWxX7OfMry
mXUF9frpNYaNteVqHixpnj+ic659u0rao+5OwAnaCjWn0InU4uLVMUvfQn66
49lkWwoaT88GjeZ0IN+0y1yo1za6QsdZxw5EPkXQ+miYU3WVeRCNvfsvS0zv
AImE//k/jTW38wvW9gudPqcfU65H3KTd3F6ICd93MAmoccuB7IHB6j9gzxht
L+Xrp3qcuXP1lAHKOYrf3RZokkhJD/jRyeF8NWJdFXTkE4dEwuE/LrWWjK3o
7AtomOfqRq26+Nq4FO96ex8mk/jSK884JjDvhVK63GXkvu4IxXSZz9XWX0oB
YA70gQO5oYSuEQUiF+aKfYpT/7LsJBLJjl9z0Q4CahkUgvmfbfFGHp1g99MB
RqF2tuHvKf266TcOTBcZC+0aNMiuEgN38HkUq6rWsjyqSJ0YvnEqqRmeV/Zv
Dg6oq81awNPmbPx+WzAfQ4CL1/DaoRvzXoQwBkQyNmRrkDlEPABoBOvCvnP+
xOXcyO0vp+eE3ZDg+77npRduA1bA2O0DD4+0JR9aM88xkvyxs5qPpC3P3kdU
RylpveF7fX0mE8hqRiTONh0tOdHVTJDDxlM877tOi/XvD9AY+CJdy82vAVd/
Y8JIXrK0li0LZiGRnNNPexQyOKpZYrE21IqO9t+MyRqDeZQpDtLUnKKn4EYA
+IaiuGwV49zGSkLvHIwhKzOqjGWrqWQNkMqdM0AyiUfo076+qApcijH8tunv
9X7xdJZSOudZWS06SsL+ZhGJMKjp+i5bi6DWnoDUJaudSPo5CaPzPdSoI6IU
g5JBtx6f/PluHrTDfj/I4gjkHV1cS+8+mfqai6nPu7iWSP/k70W/JkJIykHh
Wo8W1IVuvAi+eX3UAjO3ABoNSIX7dwCiDFOGdlXq/lhZDBOoXaTIGACGEtsH
34cpd01vEMrHYc9hv/yVvzc6tVTuBcaBYzVEKT1DdddL9fRhDnD6qWB05Js6
qRqFCKt+A/iPCep8fes4BszKONmkRecriqUPS1tABYhwMIk292jhSFMDFRVB
0+hejMs+vwBZHXS/L9oYNK2ODraF2dywYjAorQc1kneIzRaeda/rZ0Fmp44q
j9F7ufMNVRWy+WGe+QmZ1mYOZe73bHZP88p19avhKSghSiY/ix8vdu0JzMWU
agfm5XFpffay7OfDyZIJLvjU8YFw1eGwogRBnNKYX3o0JR4JDUEhSRR+B2vg
jCd5qH7r8t4/N3lF/gC0r6OxgKIMDh0+EONgZIYWQbHxPbOhaY6v6ZUgnIzN
tT/vXb1vJqkagcoDc/4+VWU523lJz+lFawQUxmJdD03x8bi3lED5zur4CYK7
0SwSOIhqEJxhJMCAzOMGGCN28hscDZsRkKANxDx5AwCZw594+k2uKYQiWI3E
/L9fiB9grEcMEi/7hKRz3l7Iw8CjqlZ5l+Xg8j3+Y/wbO9KXnx3+qVYegf48
bg09sn0nxeGs1ytRQAqeec9qLYNDSYa1seBD+sG8k+qtY1+aiCDuWvpLuqgo
n4BdjNdBa5U7sRO1tupRKBJFPJsfwIgBSHVsamF1WcaNlOvD46u1wtI6ekx2
9Vw14jtVSPttD2eo5FhzGMtUvGKUMQXHvv7rETdDVyEcHsuCln7Y3A/WgXat
UBJhc04VpIKOe+Jn+9JX4LXKhz7xojm8KOlye1LAUhQ6T2Bt6owVwF3aeCA+
rzxMsONDyhA4BkBho7Kd2yz+CnE/7F89+TxmhjqcMtDAtY5E1U3Y9LrO2l+d
EcQLwct3VxMYNHXAk/ucgI9yrTX5SCgJiw1/mX6XUWSkNKwAtRfyh7abvqma
h9OdyFeS2Ul7o69RyFfeHTEQBMe2naR0us9sLs0OyZRQyoFtoyY8iEda4esM
tZxsZnIv9HlRqiUBkoTyrqWbFXt/caTx5Drmlx6hDLVjOJpmQ9HFmxqp9Yy0
2sydCI8RFXExm3ymr9v3qye9mX3wPp6QrJNUSsuYNqkDFJtVNb2Urzmfxy5h
f5ZKc7X1+F3dAMEe2wmInTCeQVSX/R7o5QnkAtuL4qxH6CL1Pc6oNTugmcYj
LmOZnyUoiXm1FNGEiflJ7wnwZIT2Q1YkAFMcOFf0BpPDVMME9C8S9nLyOyd8
z8K9dPNGpQiXSfzi8KTBTzcqtCwermlL8GsAH4PZfVNOrzdZVoFUHE3M/Acw
tR2f/OeGp0faqDoaFj/QCWS6N8CDuv2wUBaWpJY3ta0GoqJYJvKS+1C0cFQH
OhtbQjhbAr5gsz45SAFyhiJTAmAtqHiqVSzRq6y1a3af98BZkB/QoOjVKUEH
5jJYVfCmDvvhjUCRYahCaj3k1n5tljP3dJsUgPwjlcQnc2Y99J5ruzq+4g+4
ddYAdAYS6eoBMLn3e/5uITNLfSqic4qfWlKb48IcQ+lm4Ngb76W+CUBduvDd
5qwTWr52D1/gRsbBhha4dDKY/EeBiD+/eaiN1FD83ws7r2WeDP+FNsMiJHmq
bmIawLDo18w2fpwrxoPh7kQr1AWZbZj83SMLC5NLuuyJFg8NA5lMYzFNmSdB
+XjZ688nzN6RsqScI8c4WaQ2J1ZpZWYm8BjOdVukmmBviM+bCntkXpdu/t83
BDC8aDqzjH0GKt7bepPWByYi+chiXJa+wll3l5Qp4SvKd9I1h0gHePDqHc7I
JoisFNdnQ2nddW2tLqRorUmeYONse2+5BA4yTm8otJEE1drCKHIRBoq0O/ZW
vtsas7c/PxcNl4NBaxDZirEfzrvO209YE4KOPYuktbMk19vBFvjW6Ub8C7BD
96vC+xkEiR+s4dUkNvpjcz92JEl2LbEUpUgKSFIRU9VBi8psj+5HWm2ULdn7
Kew6JD2fczX3Eqe361zJXHQBttzAbPGhbJQtKMYm6GhkgwQxVLaZu+obT1VJ
zauV+t9/tczO3KE7VC7WG5j1de2uhKQsXSlHOHanh1ZE/YHGqwARX+MHTRz/
u+jXhhHkEF/tgaPOJ8U9H7J2aoHAJHGxf+iIWdsq01JM9H2Eqw4C84shriez
a8wEBada2QIjNsmtfeNmi9JiteJZM16gXC3fSI5U6sWW0Pz5nAOURIzJx5Gp
5CnEn5/7IFTy5Jz1XBD1S4ot0CvPV6RI+uIFxkc7t6IU7J9y0ae4lleB1tik
kBU3owFMgS9Zuo7ZecoCUUEwhk2TA5ZEy24ffi6Ayp/hBwlGSMB5PMWEZLjI
cexk85ul630crJzgMPUdoWzh4r9d26oOBtQm1fgY+359cto4Ih7srY++yVzC
PceKilfiDwPe0hNDgj75qsFNfFjyDL2p+GdilmKQWyRNVrQquPVtcxML05V/
v7tXn4Ww59KVHbZ7UVBhNbli+2EihNZQ/tDQXaW3DR7RqjDktFbPhySMlMER
H1v+bgeBkHoCUUP7156q5nieuUQGWbtdDQGIrevHvLmC8Dakz7F3mjQ28VEj
ybv9zJIqxYKIgar3854lwr9U4al9cIDJ1hIrK60JEIMAxTA8YkrGXwgXRvp7
U/o+kkoQOunolze5EixA7k435ZqDJ0j8TMvlUKoJf5gpLPgclBsxiMRT+ZNU
S0zmLortLnDW6ttkbEmcq1KWgKnwLhVoAAQAD98R+EqdXlPa0q0FDr/KOHsd
sCGIjw6/GcVVB47wNOomD17ho0pWybm27Pv25HirCb/2OuYODa7RlStsPjfL
wORNMLP8g4aMwO4cWBUgv1+IywYJbvhLqhpUktOtlIP7cPA+EN89gXWAE2ye
d2LZZpHOCQ299xjwCx46n0uugWgYZzaO6FOaLpBiPE87BXVZnRsLZXvuQbb4
VNma0rqTe3Bn6SSCPEIdgwhw4qlGX0TpZneDOPdYnTncCqV0hNeAEN0v7VtM
jyK7Kgy9BzaubhBbQPNRh8bOJDbk6X2POkJt7sCOp4bQyd+rk2IgBRW5iFp3
Z91ABW0LWFF88kIaZ7n7uslFATXududSk9CLyuwGluTCuDzYJVjSZi8qOep5
EJT6lQaX8SXtw7EGw8QtqytnmTRu4nUSyLLvJAAyhX4F5weV0YYEXwQ4VIoi
A+FoB4Z0OKHjOxUtgQR83NNQoJo5jIrZcUvfgd0W/Np8dXVdO5FOcGL08uBU
3Do/SaDhaflCHn9d+hQoHplz+peWj8GHTTLU7tCquobYPUfEi5MrQzEx7dH+
StiGvA1K0UsOqX3tkV3A1G9V/Fxj5AiC4O7LJam08bYmaDz58GtrIYRkrgOZ
LT8xehvzhYqYi4giq0Zmh09sdqvT3dL5st5UTVUBD1S0m42KP869/oQ/GOdk
8tJdRhojuu6NeWm7zaICjd+mY4ZXQ0oXmvUYidwDXGkDFqvSFeCpFOAlxILs
BJIkPgv9Eoa1Ha+HYKDXz/OQvqk6bQlzNxBgmPyKPOiTRiCclKB/0LFZDNSZ
mxvfPW5H06hB5bdEzPgA4r2STwlyoPmTCSED7JWE0EfmFJAYICXpPFDhrpHd
+ljF9NF+TblrOmNrgt/c2yKXfY8ntuXV0yOu48aJyJJz3lCRMF7YCYhi8OiF
rs+Ac11T72jGmKso4zBvjNW6kjTKCMEiGdyHa3XHKeVUyuidhlGTB6SCwFXJ
rqQwOmu8jawsnJdOeAM6+5vAQA8G3TrpECovkylMq4up5RJAxjJYuxD1dG3v
fcDTIfzlg/2qguwSl4cNriUrlBGUJflTuKcZYcQNcq7ARYeiNi0gVnZxpG2L
/i55U1DbBM8mIz10YndUpT8VWiOOMs00mt2MINUWyyjAdI/p/juVwDKtM6y6
TJksxTKriDdXtGaO74bXRClb3F29LTkRgZbXQTO7TaDsDpxtW2WXvW99aAcT
XdFT6c74A8Vbck6pCRl4QT3jlrbKEL72lhFxDoOnnuxZFw+sn6rmy8LBYtfa
QYORKRLgJJub/fUHzvN8Gy+8AbXzlG++ED71qWvnDjbAErTMdxqeffTMXowe
Q9gWyzKJRFjh8MtBJFxdiRjjG/3grzwDcMrcCLKQ0u6bcyrXLZBSkbNTWd2T
/4LAXog0VKfdhHr8qtF9HvxG/5TndTUuC5nNvzbxDWw3NpQaM2AC5BCLYR0H
XMWsqn6aTLMo2dBJBqSFHJk7N21Ow2BeamjlpYvaZimYTJmbZ1AMB8dOd/Ex
ZFcd54d1wIdh4Uz43BOGsJmkRi4tV2L/JMH5VEtS/GF4/cMW29DEios64JT8
py0bkqN22uI7AK7QwL86DWoGi+tQBGXDt9mx7GJb9ZcGIJ2aFhXOJMlcsf21
R+8gUoZ1WEKP632LjcLHXCIfruzWwZulR2TKurUKZc2vZ6cmdQB1AZAHLHD+
Ch7OnnwyLxVdDNaeeWxWWTNBASpd+6hC7tKVK6r9Sn4jdRRnZoWgeK2HCOcO
ma/P3i4smeUZM10pjbldU63Cohwznp7dE7MyrwwqTjIIFPYQRFAm30/dv5sH
DjoH1ESyoPcyDi5MjiL0Zb9ivq6YJca3HdwgrI68dMxqy6K/U4AIN2QPxS5A
TDzZWDv/wdpMwvQ+bgXRJZq2YTVi7bnahBitfMXDEU2eruUjIyPdmACuuWGV
SU6fw5TTdPRy3hecNUMVkDxcPHeIrzAgDu5HJcXjRTy094cfC9tsdDP6mqEz
g7a9peAAs1ovlasI8klGRR4sXU+nz8YOprMD+G/2Y4czQsPv7FdScmK8m/uf
Ed2Mhu81xAZt+BDbVV6tntpzl/BCS+mjHPhQy1dMsM5k9kuNSUqRjXINbPwV
l43PBztb9XI+booQok0zAo2kMzdAnAi1V4Dru24J/NkObNkJyBIa5ewZfSta
5yq/dSa0cKBkIel0bK09KDZVc5TQUTWI2BwQflDBqFaPidfpLLbPzy/1OAIc
YR1+hQq9slrkLmZxgf/5k1qMzQLfZHAgHlod69hI1ErmhvK9TRtnFQWQCfYX
qKhSSR520BvcpJg8zSP17W60uIHCDyBVUiIM0sN2byWn3mALEIbx5jiSPFh+
HK4agu4nOE8T+dNq2pnq5Ww78Y2+GrFrLp+iRgf8HdH20kM4Ki8wOZPHnYOq
CvSjcMLia5Lv5i5j1XLkxNMD8jlaQf/qfsL337IpJUqfxn2UzxQuaFsDmPfJ
gO/5QWcudiE5PII9XXd9U15Vln5ib/b7RsviZSUJld0rZoKI/4OQyBqDPw28
IY0BD/rspRa6RYP3ZhPAjI6prSZRrdNRJQP4wBAMrf81dh/TtpNd6cIDbswi
2gUGKTbl1N3zcjz4qPb8wY6n4PBebmC9/b4rb5cOJDvEm/cu2e3NEU8OwDRj
fzhaWhhT6FKJJPbaBMuI5WvD9gUPFGXoyf4KiDcH7w13iBYigMcdKc6vHcGN
YtB/U41N7d9B4fVhhooSsC8q0SC3ugrhAavFNO4uMM6izq194NwIWdBGfiPy
9Cbr3lVOUc4x12svqCPhJjOHMaQoBfpcs8pNJG2UR+4UVx5TIoDzd8vMIc+/
EM0GNjux2kiwG85pNiRqQYi9WKqfBE0V/QbUJPPW4pLrVbbjWaQgq28X8bBi
/9RyhksPhHoOjD0ZZ4BIxgSOsdhBZlCAIz1t/gdvJxOBJhD1lrzW7WG+JOYx
Djzkbt9qlri4gGsYpkhiAi8mQTFidfuFXXyCkbSe9G91FGxkKw+yxtk=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qTHi3DwXzRl0JZIyv9YzFVkgChjlAUhDnpRURKX53OAkgr0D+pPTBUm9Ri8eNE4I4i53jV+DqbxrZXNVNga1DhK5yk4XHGJb1KRT3qjx38rwYeDZqT1VLOlE8YA5v53y3OJY1OjNUTOZNFU63i3NGXFvpVYqYzZYA8sx0rgwLjTiwi+CN5zXx/ep4270i7sgW87T5KeS6nNBMgkZoW2+jdSOeeOOI6BQOeN9shADrJ2yx36emt7PVeedKS6josSSgQ0TsEe2sAjH8BJLtWosX4SGP5O2tNsfBbSogxN0TYF7hSCGVSxsfbV33D4IOhW/o5BjJAnROm3b9oFcdC8hRi490KHBxXdZJ8L5IVEsq2o561yxHY4PN5cvjktMEmlGLtvAGTscAe590ZB2niht2g4ExwyD+Zg6SgdcZbhNK7t/NrYmc6tulM6mxEsdIMr5Pv5LkU+ur4JTLYUKPq6IBERyuxpMmyLUuVUkIuSMOcgYp/p4p4bCAjmP+5HrddUuftDTtU5Uk66qURtnO24Sc2yQZlVDhSkE0si6a9DWMgiKyyOsKlQUF+IySF13agBCkSQ0XwIVtPpIzf+OPa9+hUz/oiqrwJdqteJQGFNUl6uIsW1Wyd7MbnL8SYJ5Uv6ok/ozc0dvQoKGwwH2HPKxHjbcyGSPMtg+zc+c2qxVNW2A6wFBvPn5s2XQ1CVE0gI95YgspKXapx+zDTF5roKQhI5veiXx145BTeCiKs7IpimA2lN4AUqZ/wJoCmRt8fiHcBzQsKptYtH5XV020TUwchs"
`endif