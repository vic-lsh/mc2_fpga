// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KRRkh1yQ4JsNbMWJXXve+gofzlf+RpwLQQM7ZkIVKswCJOjO3UGA9Mg5k+MV
p44iqlUhGHGkwqc/f52Lnk9D92S7XQGvKWwsM2rLCj6/mqy3TX14ICqkBHtd
l8fJBoC/zjHXOAE9HT3GRkiz8PJdE11n1P1sdT0j8Cutk199qyz3ji+QDDBX
WcxgyqPsBcMmaPg38+iDwibeYGAqwi08erY74XZF2nCJu+Kin5tGlVnp+4ij
kWQI4nH9YcQh8Vvn7aWQNLVbDeN1MnXihAV8C+J52YHSGGUCxMXUItRSCK5k
rjyGrLntFv4YUbxwRKRU2YTiDvyk5j+UcSMXgKkrOw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eiCnnf0CBBO6FnsJt30CqJBAnAl839rQumzP0DjzoVMZCE69fnKQuZ5RbCbG
Qq9FUiGpYFOoMcBt9UuUVdnISR9sfBuAk/VMpAk1DcNBsBQsGNacEugPQHSW
ePCh2EXTAStvlmtJ5N6DUp8IS9JlE0UjPATZttW6XusJnDM5LiXg042Pygn2
V2knuJI3On/L5c/OEKyo+7x+SXsPCHNIcl6/SXO523XDx30NWaKQo+uAxIz4
pePoushBFlHP8fEU9fE/gMG5F9G+xl7ZAuF9BHZBX4S1UMto4g1vGT12KPbh
SCc4p9Nqhs/ABNBMfu5KkUQEqYETxpOSkN0rJSHvxQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
X4KeTxNXMSpUi3nryM6JThHrQejxOmvWhKCZBrLzWSS8gdDSGP9Xc+IaRrNR
YRlvZT5r5sJmbEmH5mGZodoOYpJo3cNEJxwFeXS7q54a3EMqQJkq3KiwnvNv
NfvoTPhkMcJkWs7dACSxSRNA25xLrQdPjVZRFGAT2z5T0KrnByyMB3q4RLJ9
lX7WWpwwb9JOv0LQ06SCnbGTdQCZcKuKYT81u3t4JFFUWMrGr32Q8vPZqGsU
wO7wiIdkSMzZWKF1sQr9kWcVCcrKYNN89lwnLzRJiA6FgOmDVGVPZ8Qvp2XQ
2bu5Tgr6XVLdzJbg1mjhby3o8aYaMh9hVSNY16RhWA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bnR0Df8j9hKIddKkbFfCKPWV1JDdTofGQgkG5RuplnI5PhrOrf5/QAbwLcNB
uUMVtkiyD/CMcx3pBJ7Fp6B9Vs/5luwUlLJAZKI8+PgwNhlP9tlGnnNd/bOP
N1W+rbY+1WeoWWVm9xNp8JyB9+CcPdslL2sdPBZlHIOW9XQZ5fLlJatBLD+A
ackoMXh0q++5wxrW1Ev24n2zR6o2Gb/iI9AbmWK/prSlh0gL+gyjoq/uBBic
OT+9fESixW5Hj6IzIOc+1I8sFM7OZob+3/4aHKtQ0kmiNhC+TYp90tvWM5d4
uUJ0wQ3GmAjMFc74rbEjyXOBoJStEBx/PyyJ9N6Q0Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bawsfqCxE9pLYi0FtI2qwp0xBDLv4GBMY7XgWmdkKknZmlIGm0/QIvXpMAmt
bJESQZUHxsXI4Uey6Djnzf8c3gCVmHACpCgo9I68qettseY7Rfxa1y0W9Omg
NeKrhoKfLQyDCrNvT0PGTuRpv9hCh5egKxRRay1+iUauDHvYLcY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
nbCcxZgfthPr2B9KJadrFY9bxudynERs1Z2eWaVv8qOnecTM18mK6ERNN8Tg
qB9VM52WbJrBnQbtWyeB/+7f7wpPebX7FXr44BXPKwn7X6m3YcT58jxkUpBE
fW7GTamjiQEypE2hATwHZvYCWIrHc4Z+ZxOGDZEle83GqyYByV16FXY4mzHd
v8Eu6bjpL0fQq8sU3bSW6iius7s78KbuQ8BDgxjEjty7GGWrlFEdPP255iSP
AzuqBITqVvDGChEIO98CILILlCIotVuj8eUVWRSWDY7hq0eWazQQw3vOBX2R
+HJxyyzIoWIwBlKtqQY0AvthfJ8oxT0c5PUuRDFhfhJHRqoxkh066MzuyLan
GH+MeE25LsRMqQniiz05mL+QmNKmj/heJpwH8UA/KfA8eTldaB/VjWvlSRWd
sGuAVpPlfSwUnqEIbaHpFlmtKTMWmJS98SfNeR5q5+9vxM81Lo3zGRo2cbNa
S4WhTI1XXVYv9zHvUIX07hegegjUe1Fb


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XhoXhz89/kAow/IiV4SkrM4CfdPIrYyqWTRjfN9nzZRMG9732IUZXzCM9uBs
MONGSU+43UfUsAESZcohQrdC0uyDwD8g/kOhFf4FwPF8OHxHho9vfNcWM4xs
dxzokm2/w6DvT4FOC6TxIwicDyh4fMWxaC4c416oBmtQUyKipQ0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DMq7oPMYqnW56eNPOZl/XpMfKtNyWZqjVi2nkeL+KcZqkQNjki6wNxUws9tx
GO5wiQiy3WpOwqZkz/Ks8GNkBv5nI8xJDqFBJK3AHIayPHvMZm3hKXcxO4cA
2gRgqY/rYOOAV6OwzTUPtS79iOWkQEMsBUXql/USNQv6C4qWclU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2272)
`pragma protect data_block
MqszfbYSSdOmNt8oq50Dfd3IncS2ArNOsg9tqyNPvfJs7wFSqm5A4HkoxxLO
MQ1jB8o7EdIhnL9cnJ4/0XqxtcCu758QsKBE/bjeFxBB/JCTlyjFid1u5kjh
AECwqeur7ELDdNc6a9hKGpNGFeT8/0PZckENj8VDQjCsabO3xUQBoG032RLh
iGF50SwY5ZZzSxxUVlSmoY+Lgre6tc3D6a/gs6h4UmqWA6e3GDa3VoWnNzMU
z9ANIyJkCl92t239N8TP61A+vgJsjncJY0K73IRLxuWoGfdGWw7WHlilkwwQ
BC/pGbH4t6hamAI53kLIsiKslnlzADizrGVQMIaGV8eiBcYZPPbQ/gAS4pHT
DPyLW8hkZGZtU0yuvxb4Idvwvi3YSixt/sHZ5oYx/hRrEZpRhOqMmmZ62yQZ
rM3dQNWz3xfILvyjxeoKiQ/mtmyQGw4Vy+1uscLKkHgSIXqoOOmwamILOATC
1WS7Nc1dI5KKEDywABqUcKTrS+SAuSwnrgEHpIMXbVmQrnJa6ktAbPMvcdJV
A5G6SRhUy9MBWJMNbZhg3SZ76W4WAnNLpwHJshwnnziX/yfYIVPonsBTt1ff
1sQ3bqeGBtSkGYqtWp/UYjmIdmKPEGoePMZ0B3KVidqP1zvX56XI8CpLuqKa
8zvFK3T4eQlQa6Z0oqBkFD9HJWvj5Nn6hKxRylpUTeo8HoF2KML2rD6fdE00
fLCAarANtyBUpbAyhCzRLzcKnPUs216ho9n2F1BaD4PcMl/o9wSwmlCx/tIR
ZRoKSWY9NLnN7DuP9pAFHQwHcUVQO1TTHSVxc/Wp0rrCIqpUQFS29k0tuzvT
UGswncF0lSjOBw6Qgh+U97BErcZ3nK73NQtzWSR28VI72Qbaueik2HTeoJD/
2CR5sLb7QgiUy4qXa1ZoAXExXfhnLdIyXkRKLxDsRwsGpIdFvkaDZIJFuBFr
MCYEwoZLF9oNdqvEC2sXFPfCYY2jISvkVbfakrGtQGFMkQfnccdolUbELYQ/
qnJ+ZOsqlGbjKnxu56YmuFqCKUuDE+7/ur+Voo/A1bwZeemgeWIxpX0gikIT
6O8Lt17npEWq8/HQQvX7XpQBPsnZv5l40VZcCcktvHqwl5jlEcBba0FVgvnm
tB37ptP9v1K/QnujVeLpJDZgarvD3NkGJ4bnuZBhIYWs0WfQfw0QsNH6Z8xh
FIr5ypZLs4jnEF2hAXuEc5bYkkSmpLuCVR4g8g63vj0frpqBT79JwmdAjoQy
E7sk5kLLP0mUSMn68/LqFYtEw2+3KxAqs1ozJBXLt1HmvzVlkPCWh9LP5uz1
aDqakb5+kFfwqOEuzGoGIHDz59woWV7JwZsl9Vq8b9UOVTL5i3U5mRLi+IGC
ccLLuyYz/Wk3xgNPfOQuOhTrzVa1i1iBcl9+U38py3O96IoaLBn5ekPETAAx
W2ujz88hDxOS1NxQalhxVtuPahB20tVsk8R7OXA2fBPghHvqE3vubDPgGh5M
/qJXxPfKWyhPGBsb9frtK7NB/6DezbvIXJ15eqDcSeyEz7f6cDocSFVDaq3w
kNB5haeyCyvzd05ZysKIiqTTBbEdyBhB4ilPg40BGFoEQQTidJgo4zsMERmr
50YRT0+9y6UHOs53Wter4+FVhfCcy8RASJIDL/VqsmLIsSF16jlG/ZVsAWzu
h0y6+1aNNWjwZ246POkxfaxloTVL3C2dhHLFMGv+X7lbBabNtBB7Kq2iqtix
IXEO3YTCKbMNEotu4/QOkZUGqo3MYhxjZQFWrw7rpd5bJS1w63aAEd+HceEI
jDO4wg1k7hGGKgco0lveKi1wOwtlbbCVZaa45GdEa0FIylY8KGYLzT5zKgm4
MAkRLMZyIQB0+ydZuc7+nqDl8JqYHZOtuk8EIsnCDCoOahFMkGVfOPlW0lF5
yWgYOoyRyI18alHcifAGwv6wONJfbPAr37PeiubJbo3iAh5b9AT4mnVrlnk+
A6Qs//ss9bfLpHj5SzM2rF4ZUTncSoM7h7n/fX9e8hFtCjOYbxyyyU4JzrUf
DfS0EnjaBaM0blm4CJLFwUEVxYFALlyFyF5UnTPfCPUgFrgC23KxvE1JVJLp
yB3c4+ORa8osmzody8AdVgXlXzDMWWDieeEi/TPSifChnQNu5EIj3GB1HUyr
gTBXc2Ri4NQCGpa4r8JKNOrEG+Eyb/2sCPJ1Z78y5ErzGAabzwyEIU4wqfHt
mFlm2011I25vl5w6s+irCURZvJljuNjqg0a1DCNtGaxZ45HG+1QpBFtiiiOV
TKkCevVUkKp2FjYDjTwXIg+l5RYuUjeDc4dG/FJCziTTRM6H8JK9kuif8bNK
ELA3C8UBmsmvj1v4HMAgWbE6urFbj5KOZ+/v+1tmZGliikhymsFMpYqxNDe2
Aac3ABXdtVEov/Lr5vwK9sIyg9IovfPr+itw0kjLZdijktAg5e629iuJmf2A
Wmp1WsvNljqulruQ3Zf4HaiicM4mRkLyAN80Pn97sbhcxo8R92NvR0kMPlcL
i0tH5S4xW1CWLhSgeU+5Qj0bgSuPrzYuX+vvuE1p/aw9iCOTFkcNctlEbe87
bT23CBD/H64nlwt3lAaJwkZTXSHh5TTSOJkLkgshGYNTp2KEXlJWm6/ANFxA
iSbAzkgeI0O7ymGv8zD2HQwruuqn3S+iciQOLj7hoSjMjDA1xiviArEesGxE
wQJNY8fgXNZTRdD8951xqe0KH2wtV6tiJI2Y4gb1NEr6vn0OwA4OPXJp2rrB
565hFS7BUj94fFjdhtoD2sVbv+xVC4oaC3pOs0rgeN7o4VSdrbMbKeSxsS0P
Mfi1BVY6y+nbnp2GZBUNuqDIcRjD9S32cWRMyFN4nU1LKWCqTrYj+L/UxJKM
ycwrlJybo8/YZVywVHpVN+xu43OGOB32T5P7KLuC3H2vvjRH3F2+RZKqTCdy
glTYI8Qwcs2e4A71unHlTjpL7B/5lI9Qsm/iS4R4opFQsBTUAth19lcZfMCx
HADORm3Y1GoBlvJ7sBJrlcfRybyl8A==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "B40jvh7ud/ahkCWXo8CJP0S9JYnc5+J2pwOdONjrEnmjRzb1YpxBEP/gM90XdEQFf8e+9j+GJABVN1VA/EUgHmy986oXHU6n9uJJjaeBsR8h22iSaiy//95eH4kKFakRZgkZDqWp0dX7AUTwRg4vZKk0rom9cx0xsiuc1Ki6fTzxDmmuuNW+yyxk/luKJogixDl7f05H1PhFx3JTfD9y6cRFGovJ+RtyYHOBbLpk0wi97zVzc5noUApADTaANZVtqbucP+HJ0z3WXCR8ycKfG/Ma/4OhU/8EcLAdmIIGnz9uxbl0hTYF/S6qpMqN2qt/dnOhGrh+RaXKpsPkQTgU5cQqzo6eUT+BzLdkogYNq0jcri6cWb6xs6s0297Tn6RcwHVP8yS0WI0OIve/MeHsUM+H8eE0pxDW/gtNCeyJlDfTrFgXUgciJ83XWckuVMZ3rcwk8QxhtGDfVg9E+0EiKm3Sxm/MU5UDzRDgH2XKEWkCZdm1n8dR0OTSXEpX1ohgL1xW50DgLAMhBHzEuwFcrXrtm84x/YG4mepgcRFTnCGoeepbLvoFB15ki6e7XC3qjcqQJPNuPDSRqIiRL6XuLHwykuEerPBM3L96JXsvCAJDj2ljovg1xci6uIkD8FW38ZUsLeh+NBPHhc3mHhZ9bdHygPJazZHgI1FUWUvBydKIHEUEuIEspei7Of6onNzmfekgpohE2SaQn/eI2KSdP0iz91LzWrh5L5kHfn7FxepE4O30QjF4U+f+SoqcDOCGjP9n2+dxXPP7QA1ezCyqly0v40NQTp7Hj12pJ0C7wEuD8Vb4CnOBTqZYaQ4h5m6zMtMwL+30eBbBw6xh6sQSu6ErBZeOUy+Ija6nYrZsuZj3OkEzn47AO61d8CDA1gKwJo8T9AiRMpGue/gAURIwmdFp3jVZM1OOtGBBO8CnJbGW1GeLysSodgUOtFgrCXkwGrVsrlIZSY0MNgK6q2icko2WisUWsBNs8FYW448LlERW72r3Ufsv5HBszHcDXEIW"
`endif