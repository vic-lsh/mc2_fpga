// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
H4kHY8PGV+qvsZPKB238kxcw8y8GB67dLF45PCzJsd3/09eLI236kx6GHQ/u
6+XEzb2RVHwgsowSNswn50lMK7rTG7sz0s0Xv+3KI/k4IOChCb9tYrkRq/oi
4v5+QWkibDLgpvo9aZxhE2UywSyh5Rowy8g5n1bBq1oZIfw9HYG5Ts/vq1sd
uJ5zd6xoLHwsjgAP0x+/TNvd/MgIur/E81Gtudm18KX/6l/Ki1nzgrn/YFXL
+9xy3AVuvMg4NkAl+QB4DdhzXZ/z+yMI23wRxsxEEQHW6HIS8extI4cRGwnB
HamW07Xior6qAd5EguzN+M7wLHduaBnGQ+C3yPhndg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZgAkVRDEpIBIoVxzo8Wz8Dk6UrO/9GTwEZPq9EhDiRiGOiG2L5U4/cpWEFa8
skmJMkjsbADclXieKpCwyUdthsMtVdR3F69Vt7cKqM0jHMLEb4ZdhPIilfkV
hO9Zu3YIayjrpL+YSSSX1YSJwVYqq1IrPN4NBO9GBntkw4DBqfxnNUQiVOgK
8DIlhg/b+VDtXwBwowsNSl+xoHvMwgmBK7bto3DN7snNYX4y9Pbn+jwQ4VUc
MqMQVDxc+k4H774jGGDVpygqTkwGn0bBh32UIxTZtK/ZJynX4M+fq6E+0yjK
58NdqJGrJRQ7W95kmGmIRoDHOpUgVhHG0C8pgE21wg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pSxFiUwo0jN8Jy1j4mTrj3xrINo8UOh1XAaIpRp8E+m4wqoACmNxCSVOy7ID
tZ2yZGE6EyFe6+V9L9HRCQ4dF5D+loZ5ABFcwdhW0nJTymttTBurarsGJGcG
K+p7hKfXeqprjoSiSEw+fV+FhpZuiPFPa0KrGOcqcPYjD7rfxPRQPC840JLR
xvsgBiSjAAhbutdA/lyNJnPSK5WVFl3nUYsQVtejeiN9Nly9FWyzg1l6V7JJ
bH6+h0up5y/Ezsi+do7H6PPAHKl36IJSTDxOD7rW03q5Vh1lboQRDqczNn0V
8n6yLU24DlG4k2VM1Px31SRvAA0jaMY78Pn70+4pJA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
A7lVNhckxadoGgTCGi/MkIfNux4TB2DE2T9dhKA+dCJSwqX7BM4CQk5kzja7
7J5lIFCumgex2RtZBiGgG78sAFATAZCb9LLLkjJgsLiWbzIc4Oh0w8MOww2M
3gdsuKWCnLUCpaiFMGe4YpdnbAREaTDXpUvaIqaQc3MO6WoCXlZu5UTF0lhp
sp+Sj3iRI+ePZcXWFVBGkkUbxEus+zzkk6dts+S2xb1s8EjRDwrUo5VGcu6l
U/qnpuOVj+XweaXrFDyA/85VIYr5aAXyHRLrjvBRISZD8ns2FGS7gUwTSvoT
8ow888WgjAvCLYaq1A6uLGMB26+h6E/eyDCFJ13MSg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UyaZ7xP0vHi9wa5NADY/11VsWUMgA6GYOiwhGuFdZyN/fKicgI0mOcuwtHo7
xWtXMdUOCytYS2YxmO3kl6C4njX5lJawlRfCfFmcDl3ymfE91ry0DwwPAcym
0Rx9kcrAVLOy5nR+whWpJ1iMAlfCZ/H19B45UzOgvUxborXGKaI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
tnUjiLaFyGpYSjLjwnga+mGh7LtZjF6Gl5+LtALZ5yydMU94w6Gp6I0TCnVp
iQcEu14f4gclIBs2kvcCN5Vzesb54j8Gx51Npv6X/Ogin1aRn4T96VhY5JbD
2CJsTOM9iyyCo/hM4bqhxPStyfXG4fndtQeLxTy1XWp/heg7Ht6W1qGH76Tt
zRTPE1kDXJJXdnO89eZbIJlXNg2Q74ocedgNtwUxjGl/utphyoLe4D27mL7N
Zfo0cGnviKZeubyBL3kI0Gjzy3Q3bKXvociyUNndJWiSzFDwSTzGmq1smxGj
UEnD3uLwhqiaKFlr0NZuJ7foI8tgCMWWR+ah85siiD1RhlK0xvX9SbHhT8eu
GLrNlwr7K3gTQJetn/E9A/u7VRILml2KMtHy2zzCcj/8SULeE3koxOkMrXWI
LOiMh0JH9FUIzxLw3LAd0ZnF48psp9PqKPle6irFSb3RF8SwPjfrHScjBlEP
B/up8flP1s+lb54QsfycViqDmbIKaVXJ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RMfSp653oyHa1+IQpm/NzgF+XnauSHdBGcKHGTKZ8TleeEBmab2M5s7EryY2
BuEocwfkXEH0w3XdfvKAS0oENwb5bZ2JNidg/z9gY4ZgMIuNglh19wTFZ8j3
AMTgEN79Q+pAzYJgghZTUOcGPjjrCYcvnBUk4KOrcbqPNXTt9mI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JoxTdtxecvB2v384IUPEIq3Idmx6pKPrKM5bw78zEdSWiX7iD0rBZ5rpvt+C
TdNABvgYjV6tbr2CWq+4A+CxB5C3Gmmz1cLxGv8gRsSu2pZkEe47TlG8DifZ
aT9FHdAERkOe4F8/r+JgnQTWbYSkEBu18s6K74T7lZCp2+q0Y/k=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10992)
`pragma protect data_block
qAc6KX7cmFQW4Bf4FSaIzybO6yx+gQGVccIiz91R+jPPT+paptiTqBs4L0mz
qBkwi5RDTHMCX7eR9eE28tmwW5g7NaKvGhwfpSerDAS5rbJLNG1JUaNBSlRr
4ccAMRfm6DEJvi2GNKBXr43Uzky90V9gHX9ItDJd+sReSkz36cRZ1Q9vM/4o
G5UQzkjaLC7PuraiUPLJk0BRk2UdcgmHT1JuDfAG7OMA7xwxuIWN7tkiv2l2
KJaCJZ9YQWWe0MhVZSNPGTWSS2O+bgOqE1+EjvxlAwg8dsHNZ/pR149W9Qf3
e9U5RWH5zukLsKalBy0Xscgp6/XLdsPjrgzfSNTee+w8a3s6p6tF00ap5AA1
lg1PM40o0axOdATgKLkhv2wJq2Bh7jbUEw0DJON9nStPXtUiROWnTGtgRsb7
rseLM3QXHpOhhhBNLQRT63FGiPwXZsQtKsAryYgWPL36w7vFfNBYlissWy9i
3uw8gljbF/X/M3jK2aptnqPlzjWoS1o91dbz1ZRZAo1UpQGOdvz8e9DfTnCB
BuwgpU5839MM2Eabbp0t7XGIIWYMdzDQfP+5G5QfGgbto7bqTYvNN85PJ9aC
n3GH+C39eZIZB90LUV139p/EH6pqWC09LunixLX7FsplvA/IyETd01rbDSMm
3+C1WA0C2phRBRUghgGH1z32ZxdItkVCBRaQjtAIWvjLPDbENj2uldzN3hML
hbbrYAbg5uYXC7PtO33jWEG70yyeh9JsmKL1cjW2BZc7MwhQJNa+kSg+wbZ0
mlMA8wV8GRM1ARVQk8Fs3/WMa6HtT7d/MOoty46sh4XgZvDy8PniotEH7/vx
JuEAcFrM4jTr2Wb4rNU/56naPQ4vQ1MCdhaBdEahd1d2IvXPRS2t3qIGhwkk
brw6RE9X9Bcw3zdQnHMgqvQXr3A02l8KKCXOdq3DfDbiN4D9XSViKKJUMFNC
a4SnKQz08Lc5qeiMw8L4ZEGWqO0cMH50WWq2KPmI9sAwtp33A3qhCWFaqH0I
23VK/nBdPAxSD6T3L1c5VHACwzGOkcQB0GjYnPjC2CvHDDBeZTQWLizpNR9U
H7F4yPWbHhkRrYW75Ys3lFeA6QXv5q+cEhhl9dyLdPtq18bT8mWPENp9pEhR
UywjgLi5Tx99oSHbCI5A/HG7EXaaW9gJ02x8yzRaDNVLUpIk57OanlFv/K+I
mSz+75RED2OG0CI38WQTKhohxzyHv+XSgsLZmFH+aU9Gr9W628Wzkv1dwR8i
k+LuVjDTi5ltS5gmzCjI2Ui7Z6aEGGb8wuDyVhObFj9mEhu0UuFoCmsV2grK
SF3REA7px9j5ZvxFY2JdH093s15o0qxBGz2FtUHDmsMZC/jtu5O3UJvZj0a3
M1cDBelUsjoenky3X4rjaM9A3y0ItzlegfgJLv4vibREAKjOlhCE/Mf94mUd
U7/jSYVtYBKqG6khSQ8ajOy2jhvh3cFZysEnkhg96mqE1IcDjGV9ybAZ9UPK
cm6Guwrl60PNKCYRtCbVnLasuRyejrHpcXndIqxBKLmbiFNnOOjoE5TjVf7l
FHlCI8ibgM8hf4VfLSpyCxxEKGjpB+RRoSZJKT5oT2GUnDKnWrn9J+aXIY6x
uvwxhMoMqWg7ZViYh3svxd8FlA5iwBjUnG9ozT607TzaIgxpv/Kre43utGRZ
ktki7bDmPgwnOBBnpIYB353y86Rt0S8vGCJDowFF4oDVDUFtIW7vZcpAFSkt
MZj7ry6dLAxfanNBkKOW/26YbKuZ9d2UV89528UTkezLMWljS6dRHvNs7Bvw
DqpZm8HL9va4ksliKt8YXidIEhTFS8JxXds28zMgaOYZ8pvP1+kdoiNgPLxj
xzHWRpBI5XOkhnEg4fnKiexDtOyng+V6nolyie/FUXsjB3eFE3nX5yQk6fur
Yfx+joM/SMN0Ywp8IHU2tcTNtrfLSRm29OC4sotuSHUXqzZ/4vAke48RBCvL
SxwVWTBZtvl5vuq3TwSUVAViPwIHGYTn7f3tsD6EJZFP0P+oy4QepdoY0JLx
1hbL+G9B/0UdQAe3I0psNey3juxwIGOI196kT7tUcO6Z1KO+THglsHfHRvyD
Q6AqrP+2E9fDEhmELuySgdK7PedphusXE4+YU4PMWuGAmtYY9V5YiI4sNJrC
XO9liGzw+ZFAKS1jPCunDTiTDt/TD3lCztc33vOA3ziga0Ogv+/bkjeY4pQf
nnBjG5DYSlV5vl/ZCcl89moptlJY7FCjx72TyLlwI74z1qlONABvjYoOnhUf
hr1tvJYFd1zV71WoUtbc5E+TQyMpd/HyHXLz+EAOki1maw3id9mKmcFLZx8k
zsj+dRpaLff2hrJuPxujG5jD6fcx0EaM8aCOusLPOGzdi4nVboAd2CO4ipRm
7X/lzUjON+dOZWgakn8yoa6xPidf/absMew98X+ZjaoqAsCJlIT2XVe3YGoc
+K7mbN3pX32DGowNwewpLFGSO+12MBlwXOijhq1SVqmMmU/6H2c27mErN7fY
//JYf8dp1vM709m/K01F3llXBwoJa2NV+RbPuWlvXLLFr0ZrHWPaASZa2NcB
pW/Zz9l5vUXkjC005gNuSu8qqmtfMFNb43eRU6AJKS/AUdNbJ189ChGKYll0
W4Ba6X4jW8D1vzs6DJ5QLtYp5FVc1ZUA9ejUkzcQ3UG0reQ63I48P3rQ8dHE
3VoK+YU2dIEw/Q2KnugHZcTp+GMBixKFGX9iVi6wMNWSNDpjcLOjSy9cHiH2
F80Bzg6GUExgjGTB9Zf6DGf1W88pay7V6LUlevuFIaFa7GCi5EyCQxF7Hiwt
dzleDngVHG7sYzuXRB9jztZt+CpeOE0ZME2sSj8ehBrDMba4W1DDZC8H10za
WOkECQb4jnCQ/VExe2HH+k66XLswukZZEVMOpDapO2wFEkR7A7oRa5y9aDzn
RSwNm4zoXo0UDGvHd0qn8aB8M7FOF+sO3f52EqQKba6n/C9vNMpCCsqe86Is
EUbbzITuVvdnD+XFwvGvul9NO0G4/OMngXsPoEMriHO+oXEzPHgaAVbqtTZK
XbLwxg3YLGM079MV+Z7gD1IMNhd51zY82HsU+uBElhcsXbYZAYcmLi1Mrnhm
xIOfZoBZmg1PV5PyI8AuRjpvgGU7nS0e77GQzuMIBj2wIF0SxkUGRAYIYdJ7
ILmcT4mIxDUZsQxS3hVSg7ks3VAznWAF30JyM/shiPGlWd9EngZf7J9cU1w/
q70s0FA8qjz6CqlzyW26CBt7ht8wDW93gBEn696IDiXKOru/854YbhNa+Gkb
o7oIcWt7jZaN+4Q7aNmeVOk2VcFtcXfhh+RS4HIH+0Lh8SPv3rsd90LxvteZ
/ep8kumdDkvcDf4l+qBIsVdvuy26YJSxcQfzYInYDUyM/5Aka+S+dbr2qCvM
JRFA8GfN1HVGpw7MDjwYCGEixSKYpTq/CecqXhy7j0n3378xc2DNMNNV1gNA
bqO0Rv+XMlo5F6RSuuju6SF7CbMx5aaprg8bAStvY/LelbISyXVmGfjDgdZI
bv44hWQmlIbIGmxgW0C7pm4jmwbxuUrwGnT2I4IiRtd/gAPKh5Ex/xLXXqfH
zvo95wrRPzLsJSxtdXzOIHIwSE0rjZFpZwOHt2knqabLlRYqdZP6UrBq5xFs
nPe2Qc63kxOPrh+jsv+YqCK9IDalJBD5t/29iAcjrLODlSA5w/Il7RPRIrrN
/u6E5XfVk1cduHaUs6Pvydrp21ry1MQb0964YxuAwLSUi6/9Jx+JYQcFGauA
fUMasOJBE6F+ALwEwdSz212q17+zGF5iD2mjhJQmdlnmi+wRgepi39RDv/5v
8MVSIIOQGWFwA3k/ka37a2RK8wKyHX3NQ87oxkKt2a3C7BwlJBTYmsPhCy5R
9KWHdwPPe/JnrAdAOSlBXpYemtvvU7I0YXfLZntkVzAsIVg++/uJE7JAcKtO
exZe2QvUqNjvVFL6mrvJt7dpOLxUyS2e78LNtnbS2uzYntCMXioqbY1mcCdh
UzXNGfM2ib4TX+l9DBH7UtsLqhO48beT3JuPEheM3DngUWyCJoXn9mqKkeaa
Vo9TcxuzNXCMU74Y1tUA1OwAulpoHw9j/QABn6HJB31Ig4k/xvab7OOI0P99
bNGqNHc7BMG7uPwfVVWa1ka641KAjP6lXiRetvIaxYqg8MBlwAoA8ggnQXOg
absY2xJ0kSKQmnsH7NXeFcsPr3UIch0UfkTxy9U4k1m5heL8fUmcwBb7aZW/
ynLQcIxU7wJV/8H/1AdAPjaFbm5EHEx45TFwd5m1HxBUjW22m37MdL1HG0SJ
H5dNrwYDQDgTUxBKFMYHbb/eXL9cG4faCj0uoeN5K58+XIjU8rvTflQIXSwP
8DR49kqkPbO+Y1XNAezjuLqeaPeKCboqmd+W2GS0DwNh/mdbPTSFya0CrBbn
ma92DWXd7CEjAEmqpEazdZNGKmAlqvavjfLQo/GgDhKPh0ROoonT4JNBxdCm
cOo5LjTn95tjTzzAi7KCR6Yk3BX0QfIG3J+U2cLf21VDaG906NdQMEnRXg5J
TIOBlimwRZP/NPII4PRBeWZuXmL0usgF3XUgc3Y0M38azIXgBoH2UqHWmRgY
tdT42N0KizursiDxYtInW40hQ+vE8nNNjKyqyAZf0MdP9mAZF/ji2uhVHNRk
g1hRtLljszbQrsCXnn7JV0dVJk/e46Y9J8RBrOOqGrjWJT6WZ3EypYMtNcm7
enWZLxK0da42Rb5/t4YHRjqKw+PmIEKlGVoco53/aVTjP5+k5zq+79ypVDL3
VOpBaT8QN0uBnn0t9VxDOqiw4DnBeXs02TqIKmoo0B9PylKABCvdb8Gb4M2n
Dfvhk5XNiQ139gB6PcxiJ45wNZzTR6zkOZXHD5Ww8qPLJxS4IFLpMgTIwlhA
qKQl4WYJgq0ADnICuVrh8nUvU5xZBDzX9EMMr/FZbUgfF4Ins5EuQUuwvzC2
ST3DR2g786emm5e/J+h8yy9JCQ9D9ayRplOsQ+W9LTgZZrlyv17qmp94mUbc
CfwHt+QhuhRUNl3fdDGqJHNwg7Ihrif4vXePs2BSj7xQgdPA5MPE85TNXLrM
Ix8J0bGm0NsXNeBiVothy2UYG5EJw1JXqRUmvR6SYeP/ZLDUZjaNgN3N//tZ
bCJCEm4MOo/y4k5SSwO462Zpu9rjMIjPnEUbkZxqFs0L1Ggqn6BUNrxYGPWF
8Rs+RPxGW7V+8qZZAjGqOx5KF+96wra6HxSR++mOulagSsIqAXrBCFHoBKfc
seP+KKn/oCJD0r3RvukpSZYSRi9w906Njlc2zMrYROZl73JZH0exg/rjqL51
UNV7FU+KKuFMa/h2XF05IasOH8l2c/M9aXli8Gwbt2n01pRaPcZJFTTs4yWE
C/9kZtPDK7n+Wq/ahUf0ig/vHft7J9/c0VkCbHeC4KSquySof8GGSyRnJo3N
pSTisGqnrRC1TIBT5eRJfYINvA5sQWe3XFnOcObjhmUNOlswPEgFhx4BciUA
nOijT1gtFuuRZCUvg0gE/BRO/2jep7cmDuVeDLIPx1CYJMBt0+eBbhje/u9u
Hc9olSfRS3gclO5TB0Ro5ZB9vSXEI1xKs3kyjNoNQdlj+JwhFlmduANjClBF
ZOt66V/QEzsX4eP8MjjBtf9+TseGiZJlbPUtcKvekYUIaof75eC1dn3Xlilz
gckf6txaXqcjRIBkkRp2X7tAIlyC0JYFKexccAqM7FBQ7Mgrw1TMgwJ6XcIT
UOFeHDQGKOWO9/nRiD4faf2SM1FH0icbZyCYXySoUdYjtLYcjwkbGp/fotbi
YswN//umm1P+cUs/0MUlIhepAKUIE0knfcjkRVrs8Sgo+g28a10sGQZzNETe
sz+bLimR9yyml25lQiJBdAYRD22sYWuYVnAyvSRl8u6sybrGIWbI9L02ygjO
zI59e+tGVsqQ0kwQIIcAtO22XG671yhKck20oa9hQReZqFVBleszb78xscFf
OT1HNNYK+lCu56CDTwq/385oHD8hzFjmxRh4Fl8AXJw5IlpaqpExouDRomJe
R1X0O3Zgd064Zb3d4qTYNaPcwkZBipyBhLm5TtTkIrR39qY1BF95FZN1ynkD
yOxy7zrN58jt/bcnBAya7afnlEDpZ6gEiKvlnTjQjHIFJzozynAHZZAePVf/
ZcYBg6D74PlIMhbssqGml4ounF9vvsPmkJdu8ycR4r2Hskn39UWbn16bA5EV
NCRP402WXlbZDEd14R4sBXzAf3w2rnPTa/0AOGzuywvwqGqn/MG5d43C6h3E
6VriKFZRUCOOz8bpvC75t8T/6VEe05Igw2xyDKE1a0qozFt5PjxGr60+FY9J
ravJsN2yGWX0P0cf1GKl0L6u0JMf9cKjWcjTRPyQHwMXxSNjEsDt4Qe0VI9y
oqzrTEjv1VuefWlyUy4W6vRf65gw1gm2yeDKh3v161X8qPaBkeGT6UJZ7hUY
akBnT/jlgFRugo2RS3oJgD1MUpz2cZCGTypfbm1Nkmn08izpz6zIXl52JaXD
9s4xq6e3xNPFvmBzrLE74tFMNU5hTikwaWhHvWQxsO9XYNeGmyBE3YSOq7o4
Z9mkhRnee/Q9BP6Pi3RILGPsYNn0ufcWuIcWoPZcllimV9RBSVlN9F6sakay
meW/UHlQlmNmUqe2LSh2M6Lh616s5qw+TeZ7FDPQ6Qf6IUUfgpz0VS7s4tFm
X/+ZKLZJxhSGUSpBIFpUHWUbGfg9nGphyETICKMXdGV2YOwPdAFa6jt5tDuf
x0igHBviloUaVWv3sc7LyGI3dbD/xirIrGwRbeLFuOWaoRpxWrorNr/fV0WB
OrCUfsH9b1QbsLQEkZ0E+5KjEIJwUxtU4hmY+6y5xV1d7OSPBNqQoTU82lio
JNFhkKmUdBuAyGeag5+SehjvF3kKlLyqmx2fZoCB/1hcyxBeDos6PKKXMsOq
py11NX8frBYeO1zKWPYtUftM+gKnkZFEPJrrqEhIlAF1KUChEjjfW9Pimpsk
hEKU7cuiVbTqiVRVF1Hh8wzARQaFqdQ2EcmzypGyCPuhfcnJ/YF5qSWhPWAN
+GBvRCwr8q8ycaMjoHF+Pu6YMicqsX7EV9pb5wdhyNjLtkm9Kq/aLhoN+3hM
TCIKlQDsDvIfZF6dpxssP+unj+zJGHzsr9UMDrSW+VyvNlhCd1yuDcwEZyK4
vGM5XWyWYhXod+xO37NKShjmvK/Y/pBZbQBsdL8mb+6raPPbGqARIQjThNW8
2KIgouJlAhV9mhJNCTFpGprUyQrOREHO9gNh36SiaZSggK5ktZERdgQlluJt
o7HPAa3NgY2sYfgvESIz0bH8ZZYgtQz3mYG3vrv/Xv50875or7cnvQU4yxIM
qw8ogfL7tXBRyxl0Mxl9v94FZgswX5JX6CSDQm1npouTyhHnSu4JLMPq4adv
d1kd9W7fKy6x2cR2eQwnS/5UcNim0/EVW4rJpu0ilM0xRAfITTJsdpnXn1qG
XfGaoWRiZ/Fpqsv/vI4sNMrn3RAYyIRys4pmry+x+EyZGu27ddSh9a/u0dlP
L5cl7ah8Z8XZDVjQTffcLN/ikPp7HzXACeXdJtoTSumNtklHNJp0flYpHe4l
+eWHWvdRtOQHGhMoJ4QSTQNUkl+t4pAh0YDmESMPWtKooEvQ5No9NjxagrQg
2U2SMAYAmxK61HeI0WafMShHx7ui9DNi2TlrEKQj2vGZS7ey+PYnR68g42pw
7WQv0a2wLqYyM/PsFOgRXpUzY1aSoOCx88m/k18CHP7UQRhMrMUGGbqd6dg/
g1Tzhxx0LfNndnfFNhZrLTqiTbBFfDidW7kM1frJoZI2dNX/lNwriKyCFD1l
VbufQZWxRBv4cmEJ2vr3S91FFvoJ4kK9FW0jrYtYXq7uV+efjeA7yQEdhvmk
zI6Tfo5StuXAXtW1HBYFKomyQvjHfxhtCykG30j0kIaofFpIwzuT72SNgsd8
xqxeQR8AsvLMYitQ7xW0OzHw34sVh6Zji11/9j2vQc4yqOK3DPDd68TJgozy
38zdyFtXN8h7a1StMQzfOSrjolGn9xABBw+8TqvLIjTJvVW7GMCpXL2zBhM2
11D224dyac9cnae+NLe/MecBK2CQ1wp+CdWEnPz7Spb3dlL7QEp5dMgVU+oU
bSAFwzHE6jTWOsv/XtUj7Eaul7970gCB4byD5lxw7vIgbMN4uY4awg8jUSas
YDT/MyTRYtJNSzUe1yfWZ7DNrRs4CXsBDCuKJm3vj9QnH8MuMHOZ01u0FrTP
ZxLkFNVRJScOfLibGxotrh2FdRtD01au1kc45fC27uc9VIEmfS9/HK4g8ixq
N9wkGXsDysZsuiEANjJGOXSSxzZXLkZBPBxpSZrfbVTrpYKAqDht/+nfrMPW
KUdF5MxTlZfV5MlHnpZe0dDcKOK/xH4LSQlM6aqfZrQNLGESVJ0h5xEKEWvq
8/nM4JUvH0R7wUIpLoRlVo0gjxeO9th9UoXD7Nmc57ufCUnMnZECKT6LIJVG
b9rf5d3tiLxbgMg9OLcD5V/eNFC3p25QyFTEsWFjZF5xiSeuBvHvJRNXXgXi
6jRLKDTTc5eCoHKrWSDxSGSr+TQ+bYR3JCeVlYY82AUxZQ4rb7BCuyb+DuIT
OUH7ZIbuoh6dYTfXJioSLP1eXl4MX16uFZ7Pvo9ll7ZmnT1ARsRrFy3p+9Es
ApJSdcSqUAvUBpEfmo+e7g/9Kkvw+6EszXR4VXQfT0iG7I2y2NNj38mypFh8
3rrYeW0TeM27Z4yrTx64Hp81u2j3gZghdG7eGdH0c8c6gz3BhgyYGTd8T8Xt
XYa+1NqiFXgZ40CbWXe6rR60nug624b3yUkEWtzg9T2U5bJRfigzFBj4pBNq
+ElCDHheKCkJ5eB9W5RrxlbHgo4QH/6V4LL2rMFbFpsd3PZ7pAhhqtiiDjvR
9lv3t/JKYXbyXxRwkK5MNVLM0MBd3bMXGKtspLWGyiBR+nu+4N3jz4VnGea3
ENDIqY5UxGLS6Fx8vNSkq9ga5M1mHjJ+/h9UCAne4D3X+7cNg8AhuBmErOC/
b54jmaWjf2qsxynF3ybjXY3VGgZq7OdshGfkvE6mnl3UcrNcpHEI9j9/VBnr
hPtA5WDBrNMGBOtendPiE4YcqN7qXvew89uWZbqMxsr30yF1n6BtKiKeLunW
H1OizOvB1S7mCJreHWsGwebEdpxaSi4twhHMCXVWLOZB11QGrwk+zYfeR0Rj
kXBP28zRxbBdzZ04buMpFlmvJX4JIi3CMPx+HrdzZcNMBp1HLKeb+i5QF+g4
MF8Cj34ktmsnIFlMP8XA4xPkQVCSevP5lK7zkcKCephRMyKJkGAzn9jqohPM
VInn/P5/LNl1mqhOxm+wVkrvAgVImccLn2cnFBxhtKcmgsECHAIYTbAeYyT6
MNMnYtFa5n9YVN1k53M1kcBBMXiGPhimgvowXCpWhspuebj/k+eHXBftNFgp
E/UR5WcnaZGvqgkBNcD/B1zvwHnQub0g8tMKYGDWwH1s6NZUAOJRpYUc2aqH
vNWZyJF90CUv7LYOCzOB2rOiNfLW2qyxgWozlxbrNkxErDP3dfh+QwdlzkuU
8PNbXFFqBRw8hxGyN3n7Ykf40H+kVNwLILMiUJo2u/Q+xOLBxpxAjEfcO9fK
BC982Q9luedQXrktba1KNknWQsVOnfLyuICS+Me3D1gmwasG+lvhW3S+jWF6
ZQO5DiGqCX6P1Di/E7jt6znGpp6E0ou5BMHthmTVPz6mtpxxWB0X20T4FpEY
1TukZvP+kkkZCQBxDDRDmofKIFod+smI59Pyvyo9wHEZhFH1zssZ1utGhehV
xV+ycHS1LWj0/6L0WQOI9y7celep0KjvsLgfnzsdP32uV0l9a4IX4BAPkXem
Mnn98vlVeyLkcd6/w2pn8hmoQ+A9TzMz7p23kUjaZkG5oni7F8LPHjxrG9PF
mg1DRjTLpXFBEn1+um/Mq5SopW7+4AfBgh5h1kPMxu2nw3/B0zgCZ1atigpc
g9JAQyCveP6mA0GTGojzxdI3YQdwz5I45KqfJhlvCxhnPRKY+har0L8qnlUp
O7zs0Up8nGoJNSHHtMJIMAe3V59LhspT/t/h/4yRSrFdO6I5IY/NxoZiCxNm
iJTQY/s/BYvzX5hx/EmBnf1s15jEzuRQN60VrYk6pkT6bulnU+YDr3c1O2yn
nUCf9gKyJjaS9lsddcpsbBldmluuwOUmKMGYjnKCpdJv5vkkPpLFgS4sKGrL
sYogXeCZAxnKhZ/RAK7++7S4I4rzU0gu3PLC0UtqtOdBtqIEe819viSO1A7e
0/923ASKc8Q5UC7P6mdNJnZFTA15Cw/+X0/R6U8oZ4k1GWcmnLNDIVu3IwWL
bPnKiDOqMOcZeNzXzMKhDrMtcaz2YeveM5pNeTTUWOTzMKOheE0peBosQGNe
gnhFla9GtzuB33Dp6q89BPbAvl0QdS3XgqzUsI/yB064ThqWWWnsCGXlNlCU
hOdPH3S5NfgSNBzAjRyYcCsasqzjRayZMDccAX90E8IVVUNrL/T8LKWuLylQ
T4Tucru0UdJIxP2bUuJBLiKy0ghxLh5jotekLZMs2srO0rYQCjqNRAhTc77L
C3IuDLeQCUSNyzGThBDlwDLaRr5CVbi99Gu0LJqwn+8pqHthhu+uSTTLCP+B
99jYq+h3EHds/v4IkQq+zUJBrI5LzmCl5nXkjq8FqUdzQAn0rltaf9Ze3AAF
Ae8CvQ5TSpZgItcJchue/xtzRfLJOeHQ09JxSIKhQu1o9deP6/L0Mf5w9tlv
Xmj/CMee96febe+ntbh8sLpv2mYLFJcvFdrhOOXr8bUtgUTEf+qZ60FztioQ
mUqkSfLtf2Vjfqt5Z0pcUK2ght8fXSfsMISlLIwcS2zDbiGV36Yfx3ACFCek
HFZVYddRjuwHyEYv9dsxJgJX+KQNNywtFKeMrCFXMHeD4Tk7CcAiFKRp+HYV
u/QmGMrcpR+PgkG+G/ku2sVT9JpP8BFmI05Ky/XuE30FgEM+zNUjGX6L25Qe
uDTaOx3E3RFguJXTKUu3xLQ7EMV9xU6mxNRMzopT8SncCJIf2dvXtXcmpWNH
69voUJhH26ggHWM/M+vv1FxV2OAdiEDAnRpdeHiNxCGX+3Hg5vDmM0Pdnkq0
sKSaCeavDLQ+LfPgFb2jBvFFiCLLGHG1OOVxgN1bZwQm2AHfRY4/ug6a3rpv
AtgK0VfavzAewzC7trJ52bpcLojD5AFMcGj2rsNfirmicDG7IazlNa+DqIDJ
42lQHS8DwyIczgXsHQqzr9WWYLf2WAajvSL1F3eFW7IX80kSiU3/u+s2Jyv1
RIAE/iEjrlLYPjivVXLqSvSiIS/BNhrlpzSJ9mrYqapzWGk717deUiPvH/xK
eWLsBeqKIj6OOBUkYXoImlLzBQcmn9AbZkWAf+IRrva8tWmBl+dRkeKpJX4O
/QvTUhzsXAsC/dgD9EqpAfk54Wr7bY+jw9THtpUd3BrigHrQT1K1SYcLGxdr
6JA1GgiycBV1Gt34xevYwm5K5JoEcFBDMn3G7DWztMkZ3KbsS5bNJxgxp3FQ
KAG15tI17Iem1ClbcLCqYQ/0fEZ7P/eYGQYZIP1W0cgl//vvXu/ONW3OcK8/
quD2EXaHV+LDBbVmttJb1x1G8j1PZC2eef0sKGy3tGAQeD0VG7smSD+COsvW
G2SualRHWPG8g0skPkMFmg4mvEkVdVUSGKnYMvCRNAB85XOGOyl9gCOUyob4
LarXOBl1/kdQp6apGjANP7E3dOemRw4W1wyLyPEEjl5aDBPqb8eftKQjELLe
5kQi2wBJxJw19S1vdM9sOChB4Nu8HULb+l827/bxxrvRnwyGnrRkUEKR47z/
1ViSF6CHX/VNbCBMMbVX/LV4ZVZKoQfCI6pUqfBDbVK9N1pu81FscB+CeYfK
GbjxYSYR0PD/McRYYSuHrWj4Mu9HoIJgIcXtlxmpKm5Gc295kMsqP7ET5VMj
xhqIZFaNy7jyIbi5J2j21VLqtuMQv/4HCSKzWCoMX2y1g2S3Mw3oyAqgxv8J
DhahvqvuwfxoVoYwneGlLWC/gsk3TD+Jkkc1AbwmnYkU/GSoCTR5H9yCH/mm
rPpgHyfxHI+HjV6ZvzCPfO91niQAgi2AkIfiHWhKGRmP8e4RREkFabshRIfb
TL0o0EMa1aQROGS8V5qJS7lYGxQe6BhA3t20B00vRXw/ftV4sZVmaBwbFFcr
Wo5237g10cOWpy2Kdlk5vxf8UgqSxBCfT0g6snaWoGeDVEgG1IEvncQiuPS8
5Oqc4Bpqy17CCIBsF6AvZ88NVRwJPTlZEkXdVaFZZLMXfB6xUcUIrRVQ8e8Q
eBuqgzt6JXgdJ6MRewu7urCCvlLtUYt9JnNmIvO8kWsPIaT/C6alOZ0h8spA
SmestpBUJMpiZ3VPCPV2SwNtZE8Q9nGTrR1qXoMq6NwfCgiqk5iADc1rjmW0
HemkBvBcG3XQn3+aRIzqPnw7lvivzSPRPBxLxCKcsN4F0RT2BMBZgU4SUVs/
/YjtXs73P0C3C/VBwlLbSW8ffp3P6vz7rFceOXhbqIa1jAxWTmUuBaoQgRx6
u1/Yqg6iV67Q2RNEh2gAOyEZRoTi1pxl/k/MbILXlX32X1LIK7lrYfLwHAer
sodAjTQZ8eTL4eNkSSCPTPBvLeW68aAYLkzKe/5A7EJip6ggCDkT1jQNu9Y3
wekkNCq2Pk4JwVqJs3NLxKXRhH1EOQhfAeNqCHQnLh2ZW6tjQwiLsE1ilIh0
EwnZx44kRmjN5QKhTV5XaqxtB2JR6cN3uRakoYvIUEttVrMlN2WLBntG8yeJ
8bbuyyEl6t4N6ij+tKETYkJbXq5QYccn49NOBM7tvxpmle83JPytrZS6TY8S
sq0SpXQIWdfKvXlRdEkdICAU5T+nZ9kbuTfOLdigUwt0f36+Jp83oLriybtc
24bapf9A4b+0s+31DV6fo8Ajl82+TTDvLSu8nLsAqJWEt2PjT/d+wMbuQMQ4
KPM96GM/G5X8pRQS0rGy7/J5N6ddX2kGGgD8Q3eooImZ6sNgn603EgMcSO1Z
zCkTSBxIALxQEhAriUq1O8nE+t7obCHH2j7PDH+hzCww1OVmUzP+aBzn7h/2
fIAiolUIdNRgw1x6GNrUc4M2NL6BzWluLoDSrzXkGGi+bCjz6Yumplf4vc8W
diAtW67vBzIG5tnisomVIF3FnfsV6YhvMUA+ZZxL5KuXcgZYEam6H0r1CwlY
LpxuhsztrYDKvWO7jjs0GF0maaiRN+tXXeEZUFul//o0pqCnePfIFIY9zdis
8ejPWPTpvyjW3H81ij9l1A/BynCD3y48ygryRbnSwQw3Xj/uHDgzHqQSO5rx
PMxU11QAOpmQRzHDDcYsKIwhO7SsGLKWEbi3RW9NjP0xg95XmKfLOGe4cmaK
z1D3H5couJZjBv2j9OH44SBB/FRXpIOUaF/MFALr6MaLNhdhwX3amQX82XZw
ol6WM432Q6TnmYPL/SzLZ/VYdT5k8PwZwxOg/w3CY0H2idqNX892c1/Ubd6r
ZS83TdNYKbdml5yB2Mg8E3hnIK5jQhNI7aDzNYouMruN/uVWxDBJ/Y57Y2ja
etWyN5dhwpwh2JyJ0c6CRAqC17JzHkYdktH4WjryO9t0SZjYI0GpQqIJhcw6
gFTUaeP0ZfT0dWuKq08y87n6BWYNjreT9bLumzwIyFmgiMINmVKwum2WwNh+
F1C4BKGHUfmMrpX3PVzlhKe1zHisAptobWgmlA05+A+Y5i7HpDRG/A40axHt
9C2v2oUfct2e2IrgFFLmWRT/cD1vY3uVuY6UCSEYx3+Sidl/CCkRBxBBOpSH
ly1VPhLSYbzx8VOSBxh0bwnCyQSiJhNqycsdsuckc97+knZw7FwgkB0JzJdd
tZGBHEFa+zXoJ46pdTEjtmLVAd7nQRz9L3buAs3Pd60BF6/4tpZ4wflkSOhC
M02fmvrK8LmYSDO404M21xmIuc9Q45FeSY+/0VNc412BdyAUM6bE0a0H3VdB
VR2lAQAN6QKGFSEVJYrU/NAJ/3++k2pQw5j+3Rm+ccVrUtF18aoXOCTae2K+
vT53abgIGM+F8g7Gc0cELlTRzh+gfVxpw0rz96HpbH9RFgjwxh0MIHbTj5aN
+ZvKRZeb/9j50UGIQpTBUtzXLnLUAq8QirvRMjRl8dPzeRCR2FykSQnIDkFo
Hmm/vfxQelUAHjINaDwmF3tiRoRc9HpbWUADeDlJLtXK1nw1TcYtstfqZ0zz
rnt8Q/vrwzoCbmneFRLcwVCPGD8RTLPqh8sJkN5LGizVhNy4k37XoJ/G/9xw
rG/QI88e29hRuaN62auT721hpH1PMFh1SSc1OkqKs/tDFeWooVs7iOsxFLsB
rUuGvpY3xIDn40goARBOdWWmNCpZpmxGQDK7TLcBxnya+9cGE+8Qibm968Y3
cHPuYmeOihhYLLNXGYSpeqJOkk4hXOD3bPPk9/S6rgIBkx8UTLY70c4YfmX0
sJd5ao/Ar8rvVA1cytAis81ul+UYnhA8nLHYiPRmZtKmvbtieY7bEDye+skE
YnOoic12KOh8wQMg014Y0KuJhii/mC2XetAacrp0uyTAAdf54dHAA+yf3vYO
L3zAV7sYr4mDXrhw

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+ErbPe4c+JM4KAwnTW0gRHqoZ1L6gh+XgxltYM1BkoSLrdSSTEAEe5LxOhUhfh1Pu6r/VJ33wL4PRvhLH3mCnBk+1e1xN8mJwNUrsuL3L+BpVYb9quAq4svZER+d/PUaClvcNAlHcxfU12qi1Kz820C7SVBM4VVI5PWir8lXfiz76lz8gB18RJdfH1th7axxPhSRc4A1rDOTx1b6eXt/+EOCm995X4b7UbZ2mb2LmKcWREalctBV+LLZruKDy1W7Wl/Gitot17fny05WvV3ferwhcWg4NSOu0+30uueMVCFdczei/rsALCnTRAs2gHXV674RSHXZlHsKYtJjjzfgQ/co0OnfZOx+R0Y7Kkl8PhOgxbfPDwB3IAA3IlminV5oTcoLEGhMVYUsVcPySKF7FMvlr1g8T5pSjStl6ae6ufzfLcueqT62QrI0Uvb6nSgm72JkEPRenvPCzHXDCSDvqSRmCN5B91prGaZLmzJgpi50aCpxNN8K6qK/cTkjTvnIVwndgQxn8GY4K91IeEdereI51UAcVcW/LpRAJ1+VcgdkbOs+QoRNl7xR9za9MIJTwAQ2LSN+WIO2ipYHPAgSSvZEKqaIP20K5cbYssxGDU18faXhItMr3/LmvTK96mD7iXbmb8nb7gKSqCcZstjSpDw+u++PABeeDkbNZPUwK75WDZagqpmhNNfZTFvcrMCHdOwknydtu7rBr3qsqzcslsMa49J2lK/5/AXVX7bIKjyJ2oYig8YTqE8KOdsnDoR1eJWLdxptWOscpQ8HjiBu7afv"
`endif