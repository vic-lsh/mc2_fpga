// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bXTxjOO5v4oFbcT/uI+wG2r19v9TwonNtsroKWtDRq1eCipjBRjekiqJdS26
GIDMkwQYJA6PvaPrpW/MaBo3Fwc7yFBBjikO6lCAvAf5QO2j5iT7elZ1j+x3
gI7cRjV6wRxxxRpBIW3j56TxxXdburtN+n9r/o+VOGR7dFN95qfJleYXR5ya
IJtiDCMbqVXW5h2kRhOY27et6T/jrIpMgxTFLrBrggbHYtelj12qOEP+PKVP
k9B63SfqlSIH4HDizYHd7D8Qmq3fZrJbe6opdxXKBQ1+NnrQtpDpp9ydGSC8
TkD9CSSnojAFkwAbc82Ewvx/4isFoVs/KxP01EemeA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dtQA4OB1BM6g+qcXJFHRtnAweNu7yvWiiN6otBPqaXCJJ88Iyhip+KhSgzn+
niVja/VxXiMR8Xo19o70Ztc3kxvlxphomYPa4m9nmu0+J3Q8tEdWfmcWEPM8
MdliP5I5aAevJKtOxLFsd5CrbSjSNw2bSwPXDq7EsP0ZfNYFoQ4pgdYoWjYq
V9u0fU+Q0mrDUnz3str/1tESZxWJuwexsJZ/kv/9HZf5dL18tAodwUUWYcM4
znwijdbQ1ayBDKDgy3tCmkYDGk/bRL1f6GVoh411yMBUdGFLhSfmtinq+qzd
5zFJ7OlK7EOZS9uNsT6tfkeRmgnn5E0suAxnK6ESsQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lwuX5DyVDRDWI20AvRXEgPAIzPxy2LMP7Uptd72uPOqx6w6yz0AiaaT0YSEc
q26yQEqiJIl2iegFnAZMjDpOhUMuww59xJ17CNBcmw5fZ8DOe6LQ2O4xjsjD
OQAhAwGWAmmL7FmPd+LDiHD+Vwmzgmu8aSxFnaUq2+0Di7BX9osPwCYacBfb
oXYciUKK93AsKj51DVfzVYFboNu0YYgujX4VYFOj8U153LqWJsypruMfkcuJ
H4QpWXyUCOMHtN6BjXZ4u3WnPaYqNaDWPhpgM9Kpn8rU9412wB6OC98viawL
gSDqjL0MOKfo+7q9NoL8QaoqqTeMROif2aafQjJAVg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
amJw4VMW+GJ+dth9HaJs87CxkAkNv+bTMxL+7v4OPbDpd5y1prD70XFmaHdc
HBJOesRUZAtJBk+GQcMnbgX43BiBqOC16zI/jsuvbKDy7ssf5nj2xcG0dUfu
wfPs8B5/2gRHkaD94IXi9JvW9r9TbghdnxzbtzMuo37grhHY+WYbmgzY0zA+
GQrAE0P9WohVqi7ELOV30equ8aLpemZMG/KBjcP5cxMiKNKfrrQ6j6szlkbA
oHKN3L0acIto9ue8zJeiyInO2NVK1nDqQXY3QTilxjLmT14hgkeCzGNlc/LW
v3SekN4f2pmHbbSx3bPOsQrpyhLiQhN1Of54I80E2Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WE18LdlxXvotIkiY6TplpKMVmWSzkc2V9S8t9RvATRbinhzjhmWHvmY1IV3y
drks5KWtmGyolDMPuHXvJgGJeJJdgKUu9eTuXbnlRLAH1rVBMSyrOnwI+6Ij
ju2DdlmQVYza49wb2FcO7YuGD9FPkXW34PoXm3HdcZ+lSEOL9/Y=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
DDwShON95tzDNJ6H20yNg57FQ76brztshS2EPX+gb2pHBfpU1Za0MZwOwCNU
W0zh0yK1/yG+mx3l/n2LeNkAYZ+LBonpLIbb9V035M/XbfQOClz8q+IGN1vd
5MK2pk4dREW0x3rKK/6+jADIxAFWKAmTGR2ze6NohT/+W3lka87qMdSfqX5W
SYeAYPe9V+PnSDwXJ60XJGfY9C9C8Kq09Wqq5DmhZuDUHj3E+TBb2KB1bDWg
AojSO96c2w65a90HzBDN2BWvDfIPR7uAlq557hxWt9tVluG6dsnaAB7Htqi4
ersUGLoPz9NkKsXqSyJiT5PvVEDzhx2ADJ0THCj+6bPb2ZYTpEzg78T5sakC
BCTU4m0NAxUPSxDuIdcH/EH+G1C6Scx0+VDKWU7ngWt9Zq884EQrrBGVAx3S
nOF2JHhvHHdNcqnVbOfYDNpKzycZD8UxwUTcCYXauw4jT55JOj0RLcmkV6/U
juaktV8r6R7GAfqL1tM+ve2lALE5T8uS


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fp/w/PZO1CB3MYjDCVpKE1XaR/7IBPNH+vTz/C4gU0z7ZENCA6joPFXYcwXs
9Q0g1RZUEXP9sroRtXQxDag2pz9d6wcMHnYBUgeKABLvuq+LLj7vKmigFGh6
O7HpaD5zfwRGbCIaSZB9a7U/sJxoRIn6nr4UUlLPNFllxQNDnrU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Eb5Ioog6lhNqN0JCi+uXkNVY+dK4HUhNsmMVTHHJZ4yLScliZBZOxJMkCHuR
iPiBQdV44aRLACmHzU+XCoDmSi27HZOC0z+fvv/oAdr+zg3YxuEfFeKvjL1g
EUigXNcz1jKbJ/ULsuJ6iKWEn1fiMKaGUVWsmJ5Ye9GLxa+K9lM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8688)
`pragma protect data_block
5HALn2N8DkYB3usVG9xq/vJaYYzS5MQBSKlTgjcW0Kfnyg9G9+T7FSqcrqqv
tRTL1J/ymPTwCni5b1KI4ME/n1ytvkDi0rS3Tqqw+nHKnkqG/4b3dRHVp349
5nEJgDFfogf6tfivrpgZ3XmovL3NBj6P9O0S29U75ZadrRO2ZBdvPcnKODgd
tXyo0GpO3VgAzUHc4NcgBgi8q9NMt0uIZLkmdTROGF0gysu/XnfzuJHNdkaT
JI57ufdjoeuS1XExX+uTIWy3pQKpSIoeVzb6ZywVcL7mEmGzLB/VpxlxqWDH
3q5xHVjyhuh4+gHtNWnG5gAl0PXCdXp23/hRN9pb/zGHPdfRaqNHKXzt0aWW
CjgkPFhHK/zsSsWfMFKiBhQEc3csByb6qNmVHfUFE3MC/xkUgxV5+dG6M+8V
faPhG7WKeYJM3JR80tbS57Jo8KSizt2pl9xDJ3PP47mrN9/hc8pTK7Ua4rdR
Qdk4cpq7zP48LHBEi6KzedaEwqdjBBRS+nRYaDqbAAZl6ooPQDciiPIRMnXc
IPuja3zyi8xqFkk+a1y73cADOgVn8lOHpN9L+/YdEGf1t3qKOkUaX8juWrkd
vROMW5nbADYoGX6uoI65sX6foZtn/cq3PoYgqdb3MzymMZQiTTIpeS3FffN9
bljgx1whtpaAxxEwn541IYqo95T+fDRw+C1cLjvhYzHNR/PxdBNsatQXV1Xq
l51ePs68bqQoYDbc/FuQyco/DYN9dJyj6PuZTX11EwRNnIg99Mjze2XLvLK2
yhGx5XQAIIX/pEX2Kun7RNHS0FEowBpNM6R2Ld4Rtu+p0TcPyBg3/03pJIJo
Hn0K2w3vVJwIwTbIpzx1l/DhROnd4QnEuJu1zYnJ0kmsVDRrD0L9FmBwlNCo
A1sXHrqU1SlOaxJFj+GPwUzUFxNHQHkLRTrlByOTuwgxNw3Tq1Gyh4CTL/Ec
JapymflRa4OJTwrYw22HSsZ3Eg77ufnPT0qPbCyJdFN698qmWKUAalFmbpHZ
cWMxSbzC2TQeacRZTOozH4EFH4LDZGJ+3W1jc143zvCXAsTX69sFRG3KhCtT
gQqHIn8VgeIkIsWLSUI6p+KP/is9zDSla5rhVMcKZA7ef5Tnqi2jx0mryoN5
I7r0DB5mWhur54Kq/DXOwSvceXFk+dp6a2lbuaBxjAcXBGekLnsvP4m6dVN4
F/JQDlrjO7ivJ3o6F9Qd/Otfp9l+U5uGySGt4ARHHFMR69tZ04Q4N46+CP++
nf0U3Xh6Fj0jwuzAazJ5MC5llwvLGCfyJ91Xmyiwp6wNk6JClVw/IL1INnV/
PjWTjQU4xnjX5e8yYNoeb0HetxQuksXUhuCLsfINaZFjV/oMSfpGieX5ADzr
LUIepOrXVOriTyknI8mmOPysFkMr+kcrp61BszAw1fnY+pdKw6/EZCgf/lun
Mt5cJXRaf+2l+pu0qVZuPOQcBbcYNu8QxtH91/gwuEjX0VkiISoaNDR/C6Ss
F2BnfujnEdwe9zUXnTD4sIQ3uO2shC6RWDMyKr6cnM0RuRCyIwYSU3BAls0Y
snHzCOhStBijkGanJZA2b1RADZ/PtkYG++HS7mUwhPKIHBUEsN181NENIR8z
dU9tgPx/9DBG6gvXpvcW2zmvn8qaCSn0L3uVSVMwKFTs52b1I8188WfyLYXB
SdCkyLyeT8mZiEDl+A64rHBSlTRaYiJj5g1wiWdb3i8UDYXRl8JugGcPAWw6
xpjWjowxYGoIQjF2kWpTw5gm9kCSi8trDbMRhWHg6wvDvUoDWfKPFk/Ix+96
0hV41LP/cY63rlbySCekJ8E0mk4TkT5IYcYtZTbw8iO6r80GHujD2Z3q6P+B
mdiHIduSL2CZu+ZFxqfspNCe56QyFrn2aoHLRM8phVb0XGTqWkRI2iTFPAAi
5pePhjpiKjTSfhfvDwJ8KHvJ9ydU9f4j3VPViPuxatrM20kA0sEMaibewVps
MTkqoHK0jRpDL8LHPyMXYG69unBALXqOBulWxtLUImfwbMAmnDjNVqiV82W5
2N1RAIN0sYZRrn6DEul//hmYTL3el4BgmX5sRqMrvyd1pZyP1ebyAzcFRrMA
ED+z/l/+1CL93jwAUulmE1pZlqSyTDqvIiQkDjpC+jPm43YWsF43tr0G9MqX
4xdxJp71nTRDGK53pzD7Ioc6oXdsf4TT7g9XmUX0XNuWxvC73mg67FD4vK1i
qwtntv9qh0PZhqPdBpt7ZOQkQloLwTXOLCQL0ExKb151s/HE5YfARxMFM/RD
3uko3uXRnfAW5SK6U3eXWCm3gNp9xDfr0WKS70mk7PAYYJ78IpYbad+NqF/s
d1ucqNah2xqhItMb2qd7MPuPY83mKpzhbtsSneeiVRPIlxCIb44f7lITZ3Ww
D7hcbzkljRTAOyhLAHxuRHVoZBQRojAzcz4uwAhLah9dqK7mIuRtsxYPP3Nt
WDbpwcypKShNMujjOA/DHChY8gpH1vWBIyNfebWBKHJPDVbi3l0nwnp/6q6a
7FhuGXTusjR6Gb30tnb4/YwubcIRElblyTJEiIyj48vt/ocBlOmHNtCcCkQE
0WCSdSSSdii/feAIwJexEuqTXJ1oFGE0uIthpz4cR7zdaH+U/E5jGa3HP+Fi
uqSEGnUfXkFDx1fbJWB5orxo78VvElSNoVZAllDlIR18laUugSiofR9vx11J
zw4hp9/qIMMypmNyl3Ugx4L1SuMpINTb78HxxmiqPQ8Xdba84hzck8rFUmZE
JlNYXvy8OQfDHzprz2iiWyZZbLd6kTvaSwthyQjI9Oy9wgCacDag9kuoTb4x
SJYo0Wag9zze1pNebMn4R3uhrbRR0GhKvgzx+mEFhVp0Mex8Qs3kXNletDy0
qQ8XpW2hqNhcOBHREGTw3RhYhwJtcmeSadgxWIfFq7WztsS6IAxPtPgBGMFb
9WPMNKkyGZKKUiGQXtnUuJHJdFeedeWpkTOyrr/Ifs52fPp4eAKCjMvW0n6J
YIuQHmTEEewt1xEPYwwuCNXMLjWvhcgVbIxFXJA81fDzsbCqrhXWrN0K7OD2
CZQ4ceu7YlzoDzCAvXM9Vv8IM5YZjJJWfHfv3LMQ7Y/p8A2/12BDk5kaO8Z/
zoGnML98ucUKET16Zl8JC5+yIXiosaLSieE3nPbLGWMDhvQlm9a40qJdFHEG
ePZIvK6z2zSCu+txyUVoCKRg+1qmQd597J7rrFI9rgpKrwTgcq4sEaqsqIgY
r8UNazJb/mNBVjWN5jaGz9Jc9iv2qsSyTW30G8+nooU2+xr2Kw9nmsTF0EwA
pl7ZGX4UHXYigKzpsxyKMjW0p6cKFzI+yGDJrFJ2ZRODA1Dr8WRrCqzoeJf8
nADBJAsED8bvOs7630Tph88mt5qLXlLpAqoRJNBn0CarEuQtEYcuHsmRffPz
AjSfAVt3yYNefz4psqYk+66w69mdKD165Cbzwz/ySmuIPJn5CVoPC5hasprl
AnLu3pa7/XfhkWiMMsSXO4YLwofWyj29lLEN62nP3I0RfY0yYu7juzGNecG1
Lk+B8kH7iDJc4BjrLAhAhxWeugvRRz+umFrmAFdaS9GwdBm8lAQYzzpJHdWu
NCtt6wMmblQ6ByGkkEo2b+7IemWbuKBfOQuZpnA4PaRnLMLyHNhjciunEDOa
xdvCjwOLncXrLoNVL2z6gQ8p3TeCt4HqCVDQXk+k9JaTHppcQusqNDrMojz+
ET9ruItVlg8c/0Cl3kSeDirdfXtUuxzJT9r8fWa5eHN3f0aF7Qg4bheLIVVj
sefEppl0JfvtiqZ9CMzE93unTq4mKXno6WWy1GDF229I09a1ZSP10Ssdr8OU
WLkubIDyCLxu9xxOxU6LhtKJ8rkmKhjk4Nc90KSIe6EmocWlU2tNpRZZZ0CC
aZQfhhX3FqFrhNJjbqWFB79CeXJ4UduqSmd4J1CPcDyTW4P3LFQfxuRILP+x
wxJtQYbjgtbiOHl0sGVttZtoeWD21Wg8r/Ix8Z2qIxgw3R4KIqLL7zJY4vil
CnQ+2B3QJ6LQRGShIeg/nXMp/qjYeOz1hVxy2BzUpduLGh5oUlQtIDY/hCrK
129LIb7tGAGssSG/vFhzych0CLSBP9j2SsavcHblyqDEZYnkXKGwQn24uzvf
YmzdS82tfGlIhQ3tFntzpAd7fQgUWZjJL8wG/ZKQuNlwnsGZGUXL5rJuWCsd
spRQA2xYMPr/ev8i9wRRudFqBgZJXyJecFECGmVEVongwtTEW0nZDtriILJr
Lc8qGxkD66KS2FXg5K+YZ+bjT6J+ZzHutFZbJc3206YVLWbTjH5ooBluFAz5
mQ3euiQTKHnBz9B9n5ebmAEvjResTEJhP+rJ9Oa0AXwfe9JQx85k6xCGbXe3
XikQzci8Ds37GdnWcr9oo/D2rW0q6EBbTrTt6K0326zAr7vy/eogPrkxvx4O
WWtrHer+rYnL5LlEyRkNu7L0Ms7KY6JV1fFSQDtPsd+iZNxnvukYvqlwZ4AX
kUgFlikOxhSfDLy3HP6S8DZr2krN5SaHPvRwU2ldtawgJ28Rafn1enhAUfCy
D7dp8kkN28UgyEomC3xkIw7WHsnmPMiWR1sMjAIFou3uMyXXj+hTy8iESE+N
IUoqpjfNHjVpzhbICPT28yjwZMAMjHcQckRRQnBB3u59KfdJLx3frhGwdUq8
uGPBGkwnfQ7cTRFeeQI2BEM2q3QMZqmmgPZQwy7pxfDjgbbuR9OEW99DWOva
vhFNTooJOghdTPjvgOgNmQQDP7hnrNvj660ko4dA8yFPmga/gi0ep28hCBEW
FFGkP449fqbhBf6STpIGvO/M5X4jNc9RrjHfZ7wxT/e7AcRgXZ7F/AnD+DDt
eZgCx8wr2fDF+WLOT3cSAK5Vo6RWEl7eMC22WK0yAlpH+a1u2WEqT2TxWStX
LlTQYO0vQTgfhY3L1oePyvbgYfEPrRnNwybEo5QdKzXNo8SHgMpTMzxbCEcG
OA2eM4K6RGgzj3pnrWMKuCc3uYE6k0bpSicZbSABP1LJ9TkX9NTK2QA4/rZ8
gHmACDmZ+LuGTPRiQ8x6LC16rNzuaasuNggDgB7AjNaAfyfRTg7/fPLJqV81
KgySzj7c2yBOwILzERdg4Rljq3CroFwmrEkdCENkFIWkaBjrtHHiWZ9+gmXO
S7Jny6Qy8XOsfTrBEWPdx2lYaz3FHeuYVgLw0TUd2uR7s7zMeKiiCEd71xjU
FG92w6c2aIduWVBOLzvyVBxXQdxcSul16Xs2Z3DIH9Xef8aEPtna7pPZXoQ6
+927/vrmBAD/+Mirml3DjEDQTGKZ1/NEibvOfnotYJwDZsy90AgLf6hPNiNd
+KmfAnp2CF/xa+1MdG3NJ5UBkSbEpri9n9lx9PvB+4SMR1+usfv6AnTbxWh2
Ue6INGpmYzcI1HLFgqj034pxFcf0/V2jLqlATkdrzS/qwRT7c8ttFm3+w8Zb
9hc61EQpRPl/ADQjnmtHjOGzRFolc9w1aHsby21Lrx1HIkAZrqVtCckT6iZJ
SXJQmsv1WD8ifzpm4V8gRJFvFm8gJmZvS7/sgoyY78lCOltwRq7PyTZ/hqGY
frrYzpiQJfhYC1VZT4TAt8OIekP4lq1zOFAPztu7rYB9jr6rqJ9erDQfgq0T
4lXIwZUfcfLQAWcuQbldtB1GEOT4tTjx2LAzq+yUvD2ZZ4Zmt5vsai7MYaxr
fVXwxSJ3EVwqb0smsWuUpIC32rqlA3hEiOq7q/PCPvbPk3feacA+MHJRcNv0
2CPaiJ8nw4LlImlrP0XCcxQ4drZj3LZz6cyIJAtI6iucOmZI7S6vX2WJ+9pX
I7ur5cefEb+j6/7RYNwfzuSN2Na2UDwdi7WsXZY21KVglChHG1HlL63tJpYx
qOTH1xxGnpwPlEAaFb5Gj8IIokZUIE2Ske3wIOUrEN3GftFNvePN1Flhq7sZ
xf/epZCQU3XICw+wwvzXOktPLTYeJCBlOVb1dpe8JgPOjzHjsHMzRWXiUxlb
53BrL2tJhj2IUn14lXffJNptUXAQCGXWXCxNe0NHhbsQkU9qMyyOfdiBnw83
SqI4/tdilgJdH/U+7mloFVXFHAZagpq07YQzfLxX62+uZLE8IOBJQwGNsyVd
qUERa85bimAQovAYwi6V7C+11hxRWY6SaZQC7RplkjWSCuK8Mezp13X3Cung
oML47xjjtDRrHwSFihvzs8Wk+okrUk7tu/AA18GPtMqkLOVH7ve2s2vETu1l
RcsrpYSaZzlG0hlrZc7rf60Y+SEiJYc0eaJfAT/gzQ6BTWlL/qHXCSQj8BA4
gMALn2jDJlqfZGz8r0OW19aPGPUw7iORUah72rwVGkBqNBLHJrJsJHudSOee
DKuVtozp36AAVondTsUdk6u9JB6mfEiMTUD5aLmz29uZv9AvUDHgWEjtxVk/
oXvDBbZD4R9OAWsGCElHgdhU0IGnZB6JzAuy9njWlKbecGW+VtxstHlHdjAw
lewila66mNNib/o6s3PHBj1ybtD/drQuqgTOtD2Me5oe2mElDpjoPiCwO2u2
GcXkRCK4yvlwHPJ1QfyZ3Ftw8+kRsSGcPUGLjBbqopxZuWRDsoujNZJgkN8C
BLhjV/b8npcsv3Jah8ErHwgtCc5hZDe/9NngRo9lXigy6pUgkau6qpZLKC9x
19ogXJGANJa3smKQVTHcMc/anSnkfS6amaaO/dkzSwSWZXrK/vl+YbqWi9pm
oB1/JJX5bl/ohCEAC1J0m/HM11RFYtPfMGlIXJxekGa6TEWLPmEEFmDq1Z+z
wxg6dQjSoK4i4Cb7MFpwjSEjYfy4SU4xjDYO05G4FU9oFuNCQ0mPg1A1GuuI
go5i7PdJD3OVnSDyo/v4EONLV9qkAFF9oAZ4AtYdw5MvwcHC2q+1VfNzs8AR
hjPCbcJ79Todf6y5L2+85h2toeEcjkWB6vxAy2KdvX9SSUFIvFT9hGetd/mH
vCFeUfMACuPu3l233vNrbjpdMLs0glL/dJ0aZmXtCJ1TWJWqvBBjywY3ZrCX
HNI+cA0xZ3/e7xFTlcu9G5lhBe3KUfANbaBhNdZU6X2n9ACb1q7qCgkTw7w4
9plMG3mT+nd7CMRINymNrHEPbHO4USItVzI8ApWZmJX3mgsOLWOTblkCeeYq
muQVeieUZliJJhC3u8CFT9j4zhdmXV3WPBdV+KWq38aQyPeo2rNvLwGyqtda
OqngSwnACRhScaYH1yrXrhtxIAaH1CAm8UA94QKAVyd7pcM4t2Mq4qRSOKnx
h50k8bLCfWoOIUb+UMT6L6oO+J7sXSdzdV08qIPOJ/4BvZPh5N9X69HaW4es
rBIJrvibElKDBkpL7vLZj7b3w9wuJ7AvIRjG1vG6nHCY2rO9BccaCHQ6OMau
HGHF1x+n49kfdau3kK40ymid+DrRsYQxvJ7XvV5qFfVARu9Y0cmcsVjXMxVd
iz1ZdbfCdV/obKjpt014LEpD06tQ1cY/rNh/v8X3xjJ7akC7Q5ZHltmu/AR+
PKzf4+r85scDrEkRzdtgD0xnoFcNv86BvmZjPcwviRIBsGXn64kuVMZouzJN
2xpv8rTP78dnsIj8pbCZ/4ojDHgOXbfzP7LXYAN3HCzh3UxsNyzm6d22F7xT
JJQdZZ/Jn28Pe26ZV9JUnKt/9VIlvyV1nBXl1eyps6AeH0asxURGI3zCn6V6
XBqvw0k9fTFXQm5EJE07U04yeDtXLyeQ3UqdTUh//0GI+Zc3S9rxLhyYSANs
06lLKbTdbGXpSnD/h3CvOVB6p2HfI3uzh3R4bRVVnyEnr7fquzOruyM5i/0L
qwqcnWWnHFWl/n0jShS6oBGNcXZ8rigwh/aMPeCJQrsu/y64unWPnAXhH29G
EDOUL370vskH3gJr4nNolFvvkk0BrLWizCT4juHNp/6OWv4ZiTHVOXwvhLfi
fKmqll+aYCBfNs4hKwmF1ofFE5KP3OmPJd0rj0eT4LsvkxcPccKWDj2rOB7N
QKLEqOy8RyKp5txfXwDjPRU5lnNB9C7v0k5/yvPvqyd0VS4LTTDs2es1RhIX
es0DfUH6Gb/0EQ8qVHGz1QWqe7ydOhWvh/T9teLeGmALrELi0XlGa0JPbKzQ
ZkTlku8DLRLNoXVk9S/+YLO92C0v/xqXTFdrvwARGLVqWNKAztO+L3ABnaYv
9Gu6VEENiuX1pQ94GRzJUrW6Xq7j5TdJQTEjCyhpvb5f6Z0cyQw/sGlnk/jc
ELxeLzMyVGweSh1y3NABw8ZObXEJ9e+LTTUFddKOvPBq+nTKtN8UVovAszTd
Gux5VsruFDbVqKLQFz4RUSwF5PzdV7LEHuAhnp4Q+2cs0Zk6TTjTTAzT4Zzw
CoZPunlvWHNXUtc4aOKNU1VbA5UvJIlIrywGtc96MFATCC0h7plm8G31XJQ2
+teApAsJO5F4iHcOZGTUvwn5ZBD2eB9uLm32JXs1W3rhWr4sM+uF163NZYTG
/4jN+HDlKxn9x+oVJwYegL9pbhrShROffL2rq3qJQzuRUXFLzI7XzmEsXVrm
BSVFiL6rZ0ZRJezRrT0sNMUWQ8T/XJdV+ZNxdbQwVIGT/Px94zS39WsHYza5
QMOkvBjAkJTB34JLu7fFu5Wb7BWgQ78AFNZh0Vbc5U34FJfXBdxS6BApbOKF
myog6VhByVA2SJm+Kxdmjqwcl72YB/w7nM/QqfuemqwEUK8/Pr7cn2GzpVMn
Nn6wXdrBz6JiDVtTbAw3LD/wZykdbANumZwJGeKEO1q7MI7qQMrDe1w2kIYX
9Yw15EfnokNQqoJb3wQ79aaAmo70pMuSR6kRkCIzHzOEJug2ig+4c/tej7uS
mx4DJO6lcJe1mooD2cxNLCnFZAiipoL8A0RD2x0XFZ3F6IT/52HLzBNBrDik
4sFmbVN5mXyNQ820IOerwg+7bZMnQRTaNAH5q6SVFM3JO77FspNJipj+XL+M
91w36hKaTn3MGBjcgmD9tzerT1H9b5etJKqtnuO9Ti3vlJ9wtkQH3qWCLfFI
9/pfOH6ik66xBGX1Zl4oArC/IjTXTIf+5ZsCMhZyDEA9APSii7glI1dUrKLy
lcaheWd3YAh1xfUlPUhetmooAQJWgm16AOPP8aAUFrOybRn8hAHUWzSruGnu
luBO9RjJbS0JlLNkQVY8r+OHDfIz5KP0CnuTMV69HhKdPiaJ/6FPAQFfbV36
CFL8C9WngDo5NlQ6iTNje+j/2ZzXuUgUFdh99NzxRX1EYZ37WWQu/YLdzITB
OgqhFlm6bQLvD6vOnQmkpAvonws8ttl3Y8S1g0M+4W6ag/baPWy8dR+aVUoP
lK3KX6hF9Zgp8kvQeej4puXt2kv6PUYs8bgrJUzSfL8ytGdllMO7eadTNLOc
2Gk+gXLZ6jQOGwoeg3J59bnCVJbNNVIxwsEb4fipBR0FAvwo1z4I/3ac/F+o
Rz7cYOCkht1RnwpevKEtLMHZet+56VGffQt/FwgZBaR/OA/8EeSUTytcPG8c
blGrykWQ/YXMRYbJPWaRuOlHMB6aGKY3akTHQkzltA6WYqIfUwW6raSeS6TN
+LK2LnNXK82TO32k0qyML4u1U7Sm+P3ezAkDnl61zd2qnxIwfFW8K8jRaZUl
h3KV4EbzVLfJQGmDIcP1fdBolqoHswL6YBa66OrZcOsomjPV3lZV55T1s7Hf
3CkGiq2PiZO+hwbUGrt6VSELpfyTM9l3A5pscM3Fe/g/ki0eP+aXusJmn8Md
jMhCBqAlgycjuNnM7XQ0vUr8AEcCmji8GddZuYlKh+1SkbhNvuzNNBp73Qz2
Teo6N2aXkE+TtfWJUJzWg80HErwlVjshvG4wPLHJYhYz9Y4yMqBlTYI5LGkf
sJ1nB0PIBWgbJ6C61Yqk+d3VzswTe8eZpHVOtXHNaZlKwkUU/TFEs91HAuBN
nfxQmHq7iytKTxFLS3BT5g5pmiAVf+XgBEjeObth3Crj9qjmqyVPn1HKpNmw
cm4OpedvBgyUwWk5XGEceSzcEf4oF590gD7vXVeCKxN+57J+pt4colMQVs74
WdVANvyB5Mym+egBGEXgspkDDhQz8SWBcCuDkGEdBHc2LMnpPaq7awbkwe+V
iiqVeRulNypj6DoIlcV2eGYV9+ByFUNbFUnjo8BXifFxBtLherJtN2yLDnmN
PaAJTaOUtStyClM9PKLqaiM/4BlaUKsw3FFPUY/V9F7zQDJ/Y4yjdoQwZOR5
dA1a9eCmU7JioHyj2g7bVZH2JJc4LM8+KmJADcmEydpv6cdJ8LNJb9ND2ieq
U7L5EQ3hXOYR7yC7kNdupOle6dMBqb8eZE4K3oHSes3eRy8S04YQ7bPjHBKV
/AnlOf3JTZnZFbvlVlUh+0vXEvR11azS7c5GGLcdqyGxCdAaxnfl0mta0Iil
paT19t65xsatDXxXL9vOm6orHLvMUSyxNyI5A1YBkfnEXR6NPksHfA/TtCIP
mrgjU0Uu+i+oCgHAyJAZGvkaAyL6IgmLibjFeNVQBXLgtHdIRTNiU8TUw2DZ
z7cHcjV3LbKBOM9Xwi3kqmhsu0+dorcgtWf991BpPYzRUNh9WFY1UATC0qsZ
pW4MTTCP1UxSXAU1fvJjyVUZWe5NYQfkNy5eepnAT90X5E+Iwr5ciQAFGjTu
1nSV3brhAKR+sjhz9CbTC3ZC5YkgSZIy2yIrf+6RJ2+TTgaxM7+2vBkhuHQT
sWohrkPmnSKVge/NfBbzWWW50JfLPrH3/bljSzolPT/NB+guflh3y5okp9v5
b/dx2h45ZNUIFk6zhJG2nwNnfiMx0glpOs9sB5UE+L3NJQuUwGPBr4i4QOOc
7p6cZgVMzy6wOqdD1PTt4f6EI4jS3r55z5LBN/k8rQKJPA5QUzrBwfm4NBPb
vWmmBaQEYZnw7y3mjPrN3Xu3OTyp1a4AUEyzghX7d2CSftkLdNe59J3WwXBq
tOcB0pr/DrcyNo6/gzmzOggawZbtpxxxRiGcC2EYnoz4FHMxJ5Imj/kCLsrk
WLFc2c/rbuZGSw0En8BpS1oQBqSqH+uFdydVVLX30GLFCFaw9k+CHqDU10sQ
/kE2cQYiwrUHZbrnrsmYgKcMukJ7ZqgCKJXummJEhH9cqaMygQuigNN8+l/Z
MU/bctM94abir/QlLFofm5tHoqpuNsGvBIZtgKP1wjYKEWf8fqibIvlyy8nf
Mta73V1wbjlhFGx7vFOs0/xrUp3ajtTnkQ0HIivEXEXnmy6itl6iOQ9nHbm/
uXGwR6H5PA32PDF/wYIIDCeSOfmGeskz+OH0NsDU/TRO8arKg8IkWTFI02R3
pxdrTwlLEo1hd2caPHgeb1ljdxTimAV+0adP9mW/fCfviQ6SQZEGs61NTQAi
1WS50y8uDhfQNwiQ2sePkn2johhAhd+whT1bZDQIh4bklo+mHZdI35To0V9R
uGxUfTypZhawtdTKQawzgPR18Kb1ag3dgLiPK1gEI7/1NR0JugbKJBIk/k1u
BIJaqHIfQQCFJJmDrIFHHIoyk1rcl5HMt29W8mqMegtzFWsSAb0xPVNHy7jz
9ppcBifyVM5qkPhpSmwuUk0bLj1h+++tDleA4BoSCwroOC8GIDBPj40fvwso
gEcL

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1KLVkvjdObzzPb7HClZqJtxY7T30Ms7W1koLcvTqhesOSo2Cw4jgSBkYZFqESf2nhJMa8PUfnGK0h0pRPoUtVvqUI76HsQ6VOsnRh/P9w3FzqopoQeQcoII15Kvr38Zh5MSzBzceU5WH1YgD8tz+UlLKUrh9kh7eT1kRe9L9s2WjfDbfOxikvpNju2FXBT7qdwVAO33H+GyCRHYKbhy3egKt02SgXhi4qY7XNbPHkndiI+mJwpsYSapJn/WBIJWOHNwyl33DJnlEsvYMKy6cjybfjMfLcuu+y6XLiMIyUIVLMpHYXqbMf+cD6WfzoboIwwsOl0EOZJz+Iohrx3GqhpN4NWGMxKeTwDYehwa2nPZJ5TDUvWxA6/f73S6rSPjDbQuDqjV0SE1byaogAzFe0fhpPadzM8rDvcyJG2Nu2/mMZ08CoLuaUuScmzMQ6RM6ynU9/yAasy/HuYZsAcbknsA1atcZbucxhM0opVS5iTn24iR6j+B5R6OzVGgWd2wRxi6kv/89vS8RDBnvtOijsJpbHHLus3RUAE5A7cSsREjoiCRlV9SXUJ80Pi3tB5xinqncg7Oiw1hde+bzmX2++ILnOfXcs+UggI9zUq3Pdz/Dw1NKNGzeh3+Ael6px8D8afYugQNpkM+R1I0eVMek1UUptu7gjmcj5aUlC5OSUTHPLAge/A21U/toXRua9LNiG31xU7yAZV09HJvtJKphbyyxCzksXC6hp4HU7XoYYahsnhGK/6E9tk8AA7K7oYhAZBVPdh4e3KTUB4xRLYh+Ez+"
`endif