// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PA9FoBDn2hevgaGKfTTQGu8SAKcVUbbVjBpV4Rs0M791oXS/npXKw1sKMEfc
ZznEwkg0Ca7g/l7qFUqBtISTsZas0S4XCaa/gvs5Ln5stALR+CnGMRxa7QMd
4pnKK6R2hvN+7o4VEM7tKyoUxd+Ri0WpU+Uol8nKydZwBZVWbc3Y7d0k2z9F
v6ixso8f5Vs2ZXdXzAf3PPg/TPN39xrCK0w/lvIGzXdio84IsM1IpiyPr9g1
NI1q2Uowl/d4qFlfL76KUCYo4PU2UV9p8HOZzfbs0JU1hiL8/uND7q4qJ8YF
+m6G+B1mVSLeU8QbEAIO61Duzi+N2Fmz5G5/PgCHqA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lSS4iLmYirgS2Ddqv7LGzeBh95WWcsKGcMB/BLwS3A4uynBjDfSjECRBvY/N
/jSBFLUpYq7fiXMLbyOrmKUGkxnIjKoe7CBayK7qBQHNhe/wFVPS1WWfsf4m
aM0D2CJpy+oVmhZrfgi8h2X5YTOEqOcYTYjiCMn5xqQG6rk9hhjQvb1KUM4f
LLROjzQStaatyK8qbxFifUdQ6df0E8P4Au/qDtT5c4KHVLB0pHNJ12qAMLjn
XdDJV7MHg9c7AyFTLlojTw3hde1zFk/dwTZGhLMTtlKHNwmgxx3HtTmGz7Ld
BhJGxBCDY/vJlmlqKzi1HcevbViOZBq4z+pJcw1Tpw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
I1HCKFy8c7io/L0a25w/3qOYt77XjYSEshQfGwfC0GqTnK4MWYjD2CILll3h
PrXXqUmWhGKyxbIrbuITj+7YmjCbeDsDWxAMthwkC+OBHYchXDtZh1KkMAnA
cstyH25V9T3idZjoocO4KjHyYYJ0MjUFsO9WISEnifPeNSAhg9UGaQGLDnBR
f53YZMIz03U7r6PLDfGGR6SGu934GaJKLGzHIJjQ3mdnnzwHvHslyuPtB/CE
WtxCEPpSOJjLa2IUVsZ0qOnQffqGEzyCYaddLNOq+ObiHlILlJ/zw+A8LpcM
++DRO/6iN9zFR0L9gYaQQnEer7AXts8zcMiPnGc22Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
M6MbV+AfQPkrHOaW/HazPrYAlF3+BpxOnHgC1N0vuyBIDg2LNyJjhr8/dQFn
8vSuXAclPlEvb4MrgOEe1YLfotgcwbZUczl87SWYZfarxp4IFtNsqcDs/KYE
b9iI2tIRK18W3eb3ySJTSACHBq0rXPlUqrjyz+IXfIYHRL88wwoUk1jyCG3B
nHYvAN8x8eqmrNv8wWMbAWU9st0Dqifwz1ydtmEOgVWO/oL8KHTlcKdwLDAP
o3DXSKCoVsA4mBQAnu10XI1wI95uYX1lkqWbPwV4uRalwd+i281m+3dnFGH6
G0xYy9LzetmpwMnB7ol+TAGfx4UleNAYm5jR3ygaZA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
h5ezR5rzmXw6fc9+/J7tYjywdmhqFDlYXlTT8TR3Jfn1Aoh1BVLQTx2a0czu
uZ4xn7vcA2neUv+ABIk5I8hnWfVmfe5ezZj1zQ7Cy86J398vK8NwnghOdYT1
mcQnThENhlLKQQQhbKpWLurt6K/5I3as8Rjwjiwbsw01xsgeyog=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
QFg/PhNMvWYQ6DxISCa3OJzvGcfpbTNr0uPHAj0IgtmFV/HT86ewCv6b0/Kz
vGr8hfMcPSZsvcEw3N5DHct/c6yj/ugl/JO3V/DOx8i3YVFZLXfLA+CPzuSD
tBoaht9SCzFw4zzvMt+q+IjXmGj03dJyD+KWULcIfUx1ntzKfgH8cCXipT3a
zcbfxCG7hyi94D5WZNGwUgMhLCKlDGohG0XvUzxuQOT1kdflDQrNNGRoHzsG
+Pv4HXGX1uWmVY8MzNvlqg/nwsLgclTChzDF/u8EvRPHFeBvIur9+z9unIwx
TZIx5NXWGguAP2IFageJ73kT7BMtgkbeD3pk4EHDzAqS24gKjaSnmREvDfYf
v59QXUpFk8nOorpMHBCd+xhprdic+YQ2Qey4ncCJ8MalmpE9WQCmLbcc53KK
7UNc/F+YnYNrz5ilDTHPeciHAPBWBCiBYrncRaz1YSUbEt/QMVJLRhZPODZI
2EC5ZyUPdGqtcDu+SPaDyuX6QMIPvJG8


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Kj5VaUgcPutFPIQj4Te06pWyxladkJRSRlCfhDUotz/HkgnGXGcgmslUKZrm
pydwD3o+KNhjqhl9NkF+yvN35qPx1FZsHoimu0W+SppJDqNMma5vKY8HqDIj
vAExyMcNKHMYI4eVzH8R0BZz/lmYq7zPTQFnTPutvMjVDQWYmyk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mn4pNVHOCvLH3k+hkSM9b8FJy/fowyM4fCnybHdgqCUHnIKzU8y5OBOQgPtY
HBN+vwue2Rsb3nJFad1aXH7nbCXbqepKYkmj9nw9PD3xQPmlESPn1Tb95VtX
fDsdYPL2l63LvOdnzildNyXndIG/t/4AlVjWsyntC3ydydXwA1M=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 44048)
`pragma protect data_block
/zht3MEvDoFrqfFDRO1UK6gjQ8FJeJG3/qYyQI76Mf4nS8qJFwlhPefCCeXg
XuILkqY2daE3EInn8CZREU8L63cHaXlqnNxoglTQSoA643rVZbJvu2PtCW/V
Kjr0aMOGeQ5zlh8zTPKkZ7Wq82r9vLbbDQCi3FXwb+LWlxG6bO4QcSJa0Tyc
9K+gWPpxlQdrllRfM+P/HsrnLIBLeVzK/AaPtW1kshN9wtjABvi6E8lPFXv8
ypkJC/m/Nmj+pwyFoogKyLAT7fCiEsj8A4jc7l5e+9xDrTbqvR166zru3B/u
dg8taEf1jgmvIuSxw4iya6bfQSQM8U8NtyZViDSCHaNBkfFpjKl4ztMVFtfM
gpzgZLPuUA30ClJhZux7giXW3bnhncytobo87gsYCf4Dl/nfR4E20ds9Q9DH
0Wi5dbKaC/eyYsSJBGteeLS0VOSB2oz1/7wwkYeWcXkuUUyTGefbYaBwmK2r
eNwTxRiDyUus5bsGlO18WdKoTAuUwjlyBTeWy1y/jtJkzs7DFRSh+sJ9Jaer
wrP1FMmMm1dTJXtF9gD7bZQzslrBgjKPr1dczn62muUiD5u10IyWjXePoefW
2JLiWddPG7AmpaT2v3Tk7nNZj5RnMi1jCxqx99hW+r+Fgf5wc3AUP7hN990M
xNPbZWYokYKYANyQVCbCs1+6HyfQR06SwfvLD+tM+2TXFez9bX+EdzTzUNzq
vTeRb4YnY/oLjiI6XyFROtkTNqbn653dJOpxLSYZ7PbdtsvXyFkRsGfcGcYb
B0tnLjAvuROqYv+Tj6Q7VL7LOAkWggMgIoSUc0w3FO/nBfbUK0c6S1uSyHzU
iE4Ac01PfWpLP19Z+7GEzN/a/uQSzzU+ooVLWMzL7bV1UEs6aAS0xLPlKwZi
sWWDNYf3b7n+RTiw5Ihk8NXWl4bu472K5nuVIgQ/uovdNBmSJrRH7WE1ooLK
f693BuoQ9Q7i973RhUp14BayWXov0+iS+rIowc3WGdEKD17TqCu1aXNVjy62
ly0OEs02qXaNSskoMrcZBnSErjNMxNn2dN0ekz1h5RYFrx4jGb6a89O1WwJC
32z37MHQbHxPGRgiCBt67rTxQvU9A4FV4JbwZvgBYiuBiAGyIj5TQhgxTQqM
rLXNMewbx+nIIhDnLppMcQH+18jT3qsL4ihbjgEfMCSgvXsKbYC+39/Ewzyf
Js2vGsOmnEfVg0kU+YPw0xFMXhDCon+PBkGTzQmTrc42qwQuTQogxDDz19jc
gebx3ElxKeE2gVEDLkK6/Y/yu9qjbb5dt2cI2kaL3MdUE0MbTJ5wf9A3+ThL
piY2v5MQlLQxNd98KGECkVwTxfoeFWeGGXPSMZud190fPHGg7glaqcn1ffoT
8h1V5aq7LqgFpgYDoqMEI0AxXwap5OhE+x1psVA3yMYOn9DL6Wp7GyQ4zwFs
roIjoYgxseCStMYd72m5kOKVS85oxbw6Ejneij++2k+OAAXDcyMWsjltPbmz
t07aZcx2kxP21jYSdiF48pdj+gDfAHXJAs2KA/JEgCNAQB5zdpoIEl4bHOCZ
FmDBXXi36GHVsJxidB0bTSo33RpYsiC/Eft0vEWFQYO/9v23dHbnK/MG3qmQ
Bon2I+gaNXGJTIZJMSytIwTVXiN7b5XKNu+99v05lg+J/BtF/DxYeXSYDyqL
7DlhBfmqREWWJ9Ujdnec398PWum1JIMfKG0Kyw06ni/m+CM980HxTiIQEYnj
+doPTvhQNa5mW84Tm4t/QuS4xhbhwntfiK6VNtCM/kdRXdfP3nzxw0ukNT28
4E98U9CoX7PwMmafX6Ml/dJEC3gjrf9687Ym9a6SmvwoA90eYRxyFe2a/gOP
HZyAWc7vxw0e2+W28/kwM2g1cR/H72fyrRUk+VRxi2D//w4spZg+BodbrM0S
O6fdzO40rZgpl60v4wv2R5IAutGkM5WOJvYMpV90+p5zxfp+x2TuuQmAVCot
wcqq9cwDT+ZBWjuF5C0R2i63V42mNf2oZlfJA6W+Q2OTFfYEiLSzbWTNAZ1H
eAePqhq2ykyMySnj0+QBbM09uynxpDEECFqekIWpZpqw/SQfWp5IWSZheZT7
Joo0NyCnNu5Pdb7+y4QRHpUg+YCp2B1WZXNhOZBiBMd5cQ0L+m/VZOlBmKst
4Q21TeNAculRdG4DAv3SuudvY4oVOuet6VLEapK7Irji8dLfLLeRfvDtASEs
A/45+BDxRjOLD57i582BOTcJNPhjGZXFtoeGiIJlIzgBFdEzQcdbPeHIN3zL
/M5RzxLP2YlWZ8FTMJqpHWvlNXz24TCcgtN/+KIH+yNsdDGhhDDQaUs2QrVw
/bGAmfmxhnOEMY29BGzPV4RrFCjYxn03GH7hZmlH2FlYlDsnTcjdej5HJcBS
teSvfCzJ/FIPF0ID+bK3atvZuQh45W24Y+7iWikjmPo1GRvz9dTKnRRoR0kn
ClbPPaH+s1TS+A8zsfQvnZkB9Dreets19LkoO+El0stebrOpD+kTLSjUmEHt
WIrVplUEEyGLcXnBYhtkozhtwCZMkmNywHETkv+MckhjJYvfVjUQq/uJzT8X
THjpqkGYbM/J9Sg1XERVD9EupTjaWPJ1QGnG1HGqCXzGnXk7edfjqBjNmDVF
WU3VC9IYGUSIEPefyQV1cjSkWYAN+ch3cbCpnpRZA+uVRv8pbQZse/9sWm93
GEITQm7avR+v0ZFz06ROyaofOcJARcBsdukeAAZ/auG+DiFLgm3ghNeJ2uQk
6DzSrimXvsEn0EmJ8j6r1lIU+ovddx8nHjdL48OQUmGT7TRmcAlaaOjWLSu3
ymRTpyCdAnXtszVH7qNw976cVHVa/xDo/aRhSl3MFhTgFshh6pQE5cERtdzF
yGVLYzrX2g17z4QxcMfMmxT6bFO+L4oMoQdP13VeMeknj1B5qkYkRSTkVhmg
Q6xKFaERwJ5j1edseOQyztwKrEgpjqz5GmZIyoNu/RNbvjo19nWcQx4BPbU/
xr+t8n4xF78OT4EPqxiCZf8WXNUy+RxFv9D2S8QA28KhrcFoKei62WEhykDY
MBqUr8Glff3xQEc9/UUW1lASStuL+W+4rtZe5ONiltKhIDi0e2tFy+OWW7gn
u3nekoMtxh9Me4VyM/6mN+r2llnyfhyRF3ix4lLP60jIvy2h78hnPHWkeTgc
Wl14FQEOIDvPRIxzbLsz2FChPkhliIMrvv6P6TKCs0PJnRqvFQOJs2OnWmMk
a2i4ZYuvBJMd+I5oONNen+0KvUfY2dYlU9SvGoJ1QaCmspLeX8igDAGDIfRf
6rYU9QucL41aEH80E8fDaWJM9HtvKYn3TP7Y6BslyI0pOcyHUX7fly7/Zx9y
HK+T0t6kvDxIqvPAUh7m78fsWsMeKjUP5DTyJfGc1sJp3VFv0jOPoUQTrfYJ
WzHopz1a4ZyjiJWiTPmBRmFkLAxvSELpy9c2gTiWcbDbwZJGtSB6wOricLv9
XsL4U3xRgA9cTE5uZj7EOxMRxAZLgsMnPlEfXQBtAKaRFK/Svq2Joeo5qgr4
Etvojh/UyTqKX6QSP93ekV0m29JqcC5HK5XJQxIWE9RHHXF2WPVzj3nN6d33
KKVQTuUfa0vyT8VDq/gpcAcCBx+5q9rFX9regsivVc5ZQqANqiXVUYmxsT3W
AszIS21Kk/OPn2CgQkI0O4KmQRqtHcWuSZEV+A5wXZaEs9+EGBpP/BhpfUlc
9O4Lnf/tObi3GebzqB12qi4HF0MW3eIWlE92cIEINGYMGQYMNsoJOM9HGaZV
RKx5VV4VlKe2+W0scTmFnpFMHSiJNdJHjZMJMorV25xv+ImPX5dkUJ3xTFNi
gjumoup8LAc23dahAaG+GNbWslZ2do21AKIkgXjcdN93q+mm3HRixhpOTOlN
nRqIs2DTrrFUoOdF7kF2CvluRhbdRomzE0S4W6e+syl8B4DZBhPAkUcFi4rx
2NUanfivqwoufOgij5/tZkgx+3urDKBQrvRBsApbC36QtlbBVov8fl4pdRGo
GZBMXBjsjoUUZVek0DgUuPYaXI6uEm5K32r86RFQ+MysBuIW9o1dxVS5yVmT
edBQ13RMv79Y3EnMOKmV5A4rvCJDVwOFIdjWb/+FRSxX5NFvH/bxc+c3nyiN
ysvO7/YliA62D7VABnB3WT7J0ZIMWpOFcdHVv5Ayg/kBs4oJsKdHLXMTpXBG
vPUkrDYKnfAVO3EMhiNZHQ8Z4D2KnI8dM2GZuClYV03bKhFoJxA+Q4ee56rb
XkVZGEJwUT9HxliMo5N/5t+BonZ8jKSmjoj+0bHYHVdp1ZeaVVdlNp9MAB1Y
jI2vSK8KlTqRyDiIHLsJoRukC4XlJ7s4ighHxSusSt87mihtke+OK9r2Elze
8C9RPGHbVnPATsT0d1HtlON/ZRPgvhDgR9tb4F7OXjT3UzLMeVK9r8cM+zYF
NQFZ2G6AQcsnMhtc185wafSE3L+kqUBobbKTp6F5mh1XGnZQcswhWSNrW4s9
SKZ8PE2+r1ca9Khy1QcG/KaSrkUOz9VekLnM/GKkwn98Hn+kpzJLERas7G6i
/ZVKCs/VderRgkA/kdeq88YPQjDBQ9p24jHy/Nse2Yznazq2gAKoiG8yCire
Y55oY1o8iagBgTTF1rI020J5+bwzF+Wu5KGrst+ca4mlVQ+j0Dj9b5aTA1MJ
kDv6EDGgraw+og9CePtyi3IuhRnRX9U1D16T9i6w4otalLuFyzqr4OsV4nkC
7tNRKmteTyN3EtXETv4mT9JGvU2Gxd2cPwhquW7tZGmSCXXZEaG72lJVANR7
05bUQoebIg5XmVLMnTewPMsQiLMUtLVG4EdZDchj4tkHuAYFgYYYwbKTzgRj
ETJNfbxk7yqQf74Z+H88wVO2QkX/GIwPn4HzYZdZ1TF/JreSvS7OIVPTBd4x
B7ApQZQoZj0ycSEZH9jzULa76EWinXESXYIGBPpPrTqzrmz74ycaIaEcNPAK
8gscQWZQQ/tJyt5mhoNpeIn/5Zn50yf3yZa4gZLwXy86rnJMTFeHs8jFfML1
6LgF3nVLBUBPiGYmuw8UxZlevUsyqRwHpqutzr/Bfy6S+mnCNBpJakDk0eni
X6GJBHhldJ6q2O6nygP2D4HdVfOL/b66oIveyTy1yGi7Nqf+DG/KWJ67jrlS
WKpTFLeKF7uvEuM+uFhfGc4BQxfjN2aOb0kCM/dI/japUzuYsJOkpgW7GpcO
G4ME9Yk4/bkXfofZmdNfRjivVJ5lAKV/e0TJ6YDTDd8N9H13qKb+YtSVd/Yk
GO4tSv1Y1UjBN4FqSbT6caVwvr83BxABs0QLteiF0YTdWDj8KlHRnqvk5vIY
xliqmN5DwsililJDSXVnpAuNK2f2QPZzD6ruqUAlqxoT/NjseZ76VaDv4gAi
dVXHcViHLwIOEJx6Qt3/KrwP6ULP6dB2GPQG9U4Q+fYxDxfD7D349mMBgVXI
Tn6amZ6EhY/fTjuyy+JrY+k2MRtsUks4ha/AJAqJkxyxmI67hf2ECh0M1VFS
dIbu3yzO5UtGQ/WxaPv7GRzLOjtQfMzeqpu8v2Mg7KayWy+zwA7by9hChwnT
vkBValVyRoALU9bw1GuYuMQlmdZSDzDqmmvFWBpagtPuqzj4VcpWerVgf4c/
U+iCN5bROqlDX6onl5XNtBQGWbQTTQ7NtGmdk8QUqHbhwodsISRPVv/S5UFJ
n0VO5dzsITWMSyPh4Y0f7ZXZtBznox6Hh6o8uRpGbsnkeYdZZcizxJZW26l7
9g4qIW+93HG/tlwiQ1Jrl1MvL3clkIDnOQfhi43un6hYttUUttQGwW7d8prk
DKdTPwoNOLhZL66YQSu+8i300EzJrt+mYmuQWdOULRagvLNFNvF7+QGjzxeW
TVzxAGXXAxsVUy3PzaF1fJcVaw/T4ayouqseJL26ewtzlIKnkvBmi7Kh+mmK
agXuhcyPBdY5dBtHWJB1J50ynDXv1yVFOGHA58ar/n2mdutvQAfffjrmS49K
ChKclIJxjCiNTDEzJsu9uqXmJZSchynrkRhN9Yv0Pl9bbAOISTbw/mEYqh6P
1DDNFw5MESaIF6zXgeKIDXj+5OyUaob7/+sJ2SI2qFI6k/474/ujdJMBFlbJ
CT2FKK4HugqfEe51dUqVG9oGPO8XDvsKlxpKW3OUVgfX874mVSClra1fr2gN
F6ZOfXQisTuz/F5TOSf9B7CrKJz8al2LHGTI1zebdpriQyI6sYqqzvYkwXoL
fnKOV6B4Acm/zAmFs427x01/W5edkKTxgSLJBUGYikzz9TIbOm2FIGKvwDSu
QBbO5zxFdf6BPMFJZ9JD0NS4FeoYFA4yiJpDoVw6B09803OMj/zDayxodLjt
6SgLN9c4EgE7kZ9vxfwwdJsWWlaUEgmTGG55xMzjyUDsB6CRTU5E64H3E1k0
IMTE/A3AM/ent/lnYTEc/3n+lrKQ17Pqj21ElVfuWoaIYON9i6r1GZlaEvQa
bWFYvEZmLflo3QZQaE0PPBaiZz0s6xGsVNLQ5dgdkglY55tNCtGXVIJDbrSp
SivfF2EZuOpCxGkh/5pnZ1HlMHBc47otGth9astsnjeViWhniJLWEWTByMJ4
PYUFp1K41okRev4u1IB8REkr831a2tm94ceYuNILYHjhgiQg6U5jLrxy15Ef
mpVqIj9wqFC6pKf5sujOZ3uQqpmOLD4LJLZmwj6DhPcdfK6gHpl6dK6eGq3Q
JkgInSNDI2USevMkJD+JBh2WSMLkSy/jQ1WCgJG9+OY7dxaScq23HkH7RcvB
dJ0UP9NDNFF1VNB4acaBzZsZvNHI+JefsoTdOQ5hu0LukfN2Mvte78INeUDV
JHaIx8ulp5n3+b6lPnTdOZEgQnrSvOwMDbpXsXoo3MPQ8YQzbx6n/do7TQcV
efyTmR/9t4USf+C/7Omsi6KqvmVvC2TKTwPGqNxY4OQfkdeuN4oaf6sNcGGm
UhT/LPB2B+Q/xurwPDDTUu2STgAMHRLWpQdDTENzR8khyPoSu85SMsQRkvi9
yeNeHIbFcoWqWMce4fTMUHe72sYRwpC4iCp+yeZYu7AnVt/rNfr/L9jhQND2
HHlLC3MmScSH4I3f3A+ygmI02LOu1MmjtE5750hhDwvoWR5KOYqEho/xSfjq
9h1V9RzsfBF05HOJ8Qs5UZolIro8GZ++bgl0TxrTIFO8ztAvhuXSbX91LN+a
TWsouBMj0HVCdKdA87uVTdW7yU2zrgydhKw4xxJ3bJ6e5X1Gvo5N9FSv0uJe
0FTnALrgtb2PXV2S2YSSNR2rFnfU2TplX9EVzXI7C2yGEFAH2nU6H9aW728R
psNqs5FK52KJJSBJTnlJ8hOI0rTirmv8W2unNainzSUdBr4/nmPrkZQdkySZ
/7rl9VjExwhPc7w3wkJhGtjehWRTqppAKUK34mINvsRxkRAA0i9AZ97oxerp
6GdiWfI4c8kHZ4YkB9dcN1YuQKd2iQwWDozuQ9LCkABYnh0v7HWg1CiqIfn8
VYxqJiK+7S+JIvhgKn72Usq8mjMT6aNInwuTzIvyumuECtwXFkwFEHjaYX2n
URLSDy93+doZZf30X7ewk6iHE2St0KxYNSrJS+7ffpOZYAwRGzb7Gs3/2bPy
wpDsPfllI/UfD2WrgtwXDYIgksocE0KOVsH/7OFawRGgVgFn7WNYzc9pv4l7
RnB+tVKFbsa1FkqU4uVtmAAYORCBnlkUDaaVaEA3fWpzpF+VBwtw8ZPrkmeU
AEyBECu2IVn7LqOiKZKEwFL0M5rmh7gD0cjF6BzZBrQWZVyFMH3lHocF2Gjn
wZ8VICVDoXpu/denBB7OTxPHqy7oOsCH9O40gIdfaJDx3pL3rnom27uMiPGt
BlwjfK3YBdP+thbNKNTAyae7kSUq7tAkhz6Mno5hp9MfAxkVWhz5nD0093Es
otYZMUig6u/+wIQa8h2Zr5WUkJ3yMjTQcOcrZlJ4oh+wI5q6yjg/MwpqktcT
UjuDuxmLHOqbLrpNDF3E+geiAqhLPRGnJklsCWsQbf4DdPlowtxDE7SQKEoX
SrcA3C1By7bNGMhqpvhuXQrxCh8UGVVwd1IDUD6JHhg74wYshibsfjOI+wqc
EbHRAImd8FCv9NGCe0kWM/XBhrSk9KpGpfzdwYNw4eBzsKwWtazs8orzAigH
wHPCrGwpzRpN7BX5WFuH+Qzw9NxBPKHNiW7RhzzDxfypcfL7WQo1cDDGhq0h
2IdYJinzksRUJkdsQ34EOqKDUDLGF1wjmQajbp26zwONYp3NW98OcZwy9W0C
wzCkZkF98nDyE23zCvQFmLOZbXYceBBNF69c6HY5ZO/1uCEB27ttKfV6vNnq
+POqImEuOxuxezZbIVZXD2t/1fpN1IlferBdK5XmBKAXTrp0Gqq224934Qmv
VkTzN6WIO40sOnaS/ZkAth74W6FuPBtjXHI1AJqJkhxN7WtWiDfhasSzhSVS
hbkz1PYvjuXomOmA4aAhoinP0jTbrh2owuh1x912UcAWq343641Z6awPl0rW
Ak8UoCqcl8+810A0eQx28c02soXbfHL0Jd82vopOUd4cJAYr5hY+J4n/BsIW
+8EC5nenCXQwpIzen1LnY6eY5nSp2rev5yCf0beVKVPLstU2+VpB5Qh/Oda/
RxXPg13asBQzdl0DsPbA63sXSxdCziTFJLEttAJfEYUP8dZdp25KaO3Hzt40
Ruv5X1ybIFRg54HjqEqyB8uGya536ay/+ZkNySq2TDHenk7hqcFZY8znwdP2
NYmoVWz+DUZwtMOp9zdSxNjWVthqWFUiS4S3J+WqsOxBDr7c1kGvp0r6gDc7
rlseycavKIYwkFiYWUW0B5iS44k5vQ+hJm4jvyP/bHN+8C4bwzTSGHToSdbw
TYU3fEcJZO+Qd4xczB+7sdkeXcQmaKTmvuHP+twGvwNvZkg3zTENuQTtyiua
z6lWxJ4XQlC3C1sFbReqBXpebJI1rZLt879IbR4O/EtcO5UQ0eYGLnyfHTeu
2YqXoum6/XgFLc1EOg5RLh74QpDQfhwaE9q5LkDD0Pq0mIEUTNDFEc5cL4Qz
2sSaAIuA1HkXESj9tuKS/521ky+aZSV56r6Gyk81Hz+orNGQhQ243g0bQ3Vl
dK/mo/qWoae3QTTL35bfJswbvsEe49sei2joHREJMVgHtyDR7Figb3L42PXx
3mIjjHGDK1I3PSoZEC+hsOwagOLweqzccRQyFzM4lo7AYBd9T60eJogvRbqm
DPzDoNZfJG6oeBe48Es0AiJPnZGIeX0iDnNiQV//oZZHGyqkX+t5Ilg8KD4u
Za0qcl0PWxbvs4c2zy8eabCKh9bX27uEzSi+kqWAVmGjKDHQnprKs7LXCi1N
OBIzPS5L9Zc81SwQDpDr1NdqRxgha68PXrBgV4kNFnwuzfJoIzGy08Iz0CMy
YrglAq+iI89j8rEw56a6wmg6+FfUvpsdoUf7WUFauHuietUethpV4ODm69DO
x2eH1JUsVosstmqOZ65lPQZNzcarYA4rx0+l/jDktLRW7f4GoZrAzKkg4qD6
QOg27FLgTJVIU386xwCmlnVCggrjZM1UVGnORQLKPkw9YOfEfkWOBVJgqXk9
hKrLuki+jyZ9lYiGi0b3V7y/dEKw1sJKC/eTf42kLncO33358zMBulJL/0dB
d3LNvxP3lDfK6Ovy0FFM7+PU6nncIx3LdW/nSeN/GECcfMVF7ViH43BOqRAy
9mpVGk7PzZmkZ3siJKWGkD/rW4aJD/OQroFvXy3O9v2uwxTI57lpMZzKHTxP
WZzJvGV556CPWErfFO68NrV59RTCITQjSANr5RcmAOX60c8uuFG54Yeme+ba
CX0604WAjNqw2tDpvQYUQ0rY9uXqzMO/+wlazAShA36/ldDuTgy8QzrvLEvl
xuN2k8BWcKkzq7YmWdHfbQHiflfj8Gri7PBLD9F8FyO5Hjwvp0tTU3JaV/fk
iPx27YTGdBlIVQMfKfIpVCHNCJNza8Mi/+cEecGiAJNPca8B+DA6Xw73ZBhk
ATIwAhH8Hj/DJPPFf2DqxIMHOb9Yss43s8CylEWFL4/fSgANQbN7z9bbg0lr
rvjb2QODitk12yFsZXZLSWZBs6EBmSNdPa2o6QpuOYbYRaRh6fIyTBePqCqI
EGHfdriCHJ57p89WHEDObs64/uFzUR8ROJDWAPTA0bjcLh9dBCgdzNHIatIi
+KYOb1Hl9w6tcMzD1ALy59T07uBG97uNlaIVpcQMlCT3T8Jt/+Ulnwew8umS
B2R/ZGpxhcKIMiLoX26g9A1QeKFX9yEpga4utkILmyDe/7n86HUDSSqyv7g1
9hVHbgjY56EkbkZmFcpBwLmiJR/Z0iz7SHRvh+I8eRB5vA0b5LhgN88pOI21
TQXenoDiBcPXJJZ+0eGOfGbGrGqGZDRt+6jxxO246Mwl0tbRKA1+sloSfJzZ
sAuDkBZ/aYCxfzXHYzmJH9iYXUQvFLP9kLnhFxskJSqi4ukegNabFXDs3vzc
TNj6cOpAqajy3i7hoYsTeNyJgbByCC8VcZrs/Piwai/ncqr/ap1u92MVF51F
oqSYWwucqaR7ULBdq7bPUVd82CBMozjBIc+7TXYmWtc5zJKMTiFQXpSZp6/p
YAZ+hG61aQ9Ev1XYl8FssF8JLK10uwv/veaAdB01mnKTSrHgsQSk3n2D2SBM
7MZXXjx1nbdTFIwt7qGdlo/0oWa/m4yMEAjyhYqChxlio3itW7yj6j8bbp3M
xvlSWNbX5Y+cbN34+JNYUZsvYLwDAtfie21rM3HDpmK0yZojQB/LLGxHCMuU
lo9byBW9/c7JViiP9/apVBwRPXfxB5fqd0RtoDuohXLsBQ1nQbtUZHNkrMW5
g3a0TZmBdAGmqaltF0FxQTUPilzNrKuNAajFAhRXSPeUV7dpcYrn5oe1K6XE
ci+omdZceaUdodfGRXq7MzJCfMK6BgBRx6hDLh34sSbUoRcLH+/lMlGVZI6r
Qq9O2nWiYoKnwZ/mrG/nFcwdYYbKmvjZlV4DDgJGVyGIdVwO9Zs02Zlcd6VO
Bp0lAcozx9O5xRP0BLRzgMGWTY78HZeM/QMdpNEzIwcGxpifT9VEYAUJ0fy9
nm/HdTexfRYy1aeap+RchinFDHv2yP7kUH6C6sr9FSMTjzlimHK7piiz/Wi+
UfiPbTmjCfhyVyMtbqHaNuMoxkmQksoCOmHXTkcHUKf80zHqzbYU4TUPYpdc
dvT37RYmz5f/S2Cg2qiFCYxNWw1cVtc3pyR/A6YsjcF5uOgOf/JkZqpMpcDT
Ub3zHjffwUE1Hjy8PjWRDQqTU2EHqM8HMtL1E06zNylHB38ObvzvD/jaOM/j
xD/JquFuslQxHmHQYV9LnYYR8R787x2glTStrOSJ6e6muvp/feaFiZCzaLGF
nri4DPnVegoz0f3tRty1aHzvCwfoApYEmK3z4NUt2SGeL7WhY33YJgisSvzQ
4hQIglP7gEHvQWz7xamcSzDGTUITg2uIYWOC9+TF7VVQULttsOLHfv0QENjF
2v7wF0zCJ0BGytsISNfYo/xBYEKBRKEBOkd5FeyVu0Hr9rmNO0ODIQEzGTsl
TN4s+h7vuzpKvgDgMmjcYsbZDDD6780jceu3xWkqDJgSj9CI0AoZ5tY6cYk8
PvGuYVFpXtjJRRkuHPy3HsA1aIBgec9l/Qjw0k5tvA3DL/MgR25k9bzf5KHW
S4QT3zC+Y58j5d9MME0S/xr143GO5JcfDOUJ5OlaesALpDoS+7AWpV+cxK8O
MzINdPTTr3iA2C6FYgS0SvvjJmx/RiIk6BtrQVYYWvUM5gl54wqjjtHpyEZj
lbO5q2c4IHVhomuITCJLBIVVIjrnBBXIUivsKbVNk/L1yqmwmGxImoyEjnQY
NFyqi2UdT2pVqsIyG9y8fDmCJlbyb5PUTFu0WP8R7VpS8jEWDEEsEeFVwrVp
iNaYbtS7mpMg68Y44mAzxUc/XWvUD+svjB/d4xBF1JmsfzpISNG3AnOU9wdX
UTgRDhIoNygL6INN6RR2cCOVtR+gse0bTJhUKx78jdiEF6MZFTy72e8mgYgQ
EvOBRJYoThWSxKg7/TzRLHHcfJTc/TuAMlg8/XDZkwZTGq1Gn3ZMAEVFSUqP
hoAJk8agq1AgBzzLG+K/8bwEfIcPkouNSEOg/V5WA9VBqMoyq0A6GvbbMMRS
sYaj2kJSdaCV1sbwWXoNOL8gYQLjNRYgcKKgrw2htWrt63px7ivo+pqkl7tb
JIDMiz/nTQlFD11OPjdsSIWES2tO1HGe+THe2Ex3X4INAgjP7GM1vcDT+Jl7
HqX9rYykmk85yRvWszrxJbTZhySbCW8kdoUS+/vhvyl5yRI5YGTgzRymbzUt
G0GKTXYZiAd51PkC4kRCyV/lHXSwfuHg9BNuCJoAg0+j43XE2Y+xvk544TST
7k5Xbcd9SeGZ308hbhy90iYbt0lbUYlS/Kz0FzoFLHidmygOGDJadHDvWjGa
4PU9TK0zUViTO0cyvdBwhBCpDIJHsb3lVJGpcDBPKWStMmQHV448s8O+N3Di
tOugP+bS7EF+SzObJsjrzKvCUyjtbHqprgOIiUH05/slZKunD/Qv888mfW96
sKgBxZrW0opnULr5DyxviM6t0DwqyK2ATegVBuj3SpW2guQ6pLQahAMYPMHJ
x28ttYIly60XVZ57M+pGr9LkqzbtI6BJww12HKS9u9DXsf4tqEC9IPjP6Vg5
/V7GbLT5+Tm7ybKyHgfUNcWczX41ntBkSxzeeEfhzuk9CSrYJ4Crjp4l8q3Y
ede1JamNHVqBg9M6qKT7okS6zBneUOEQeyo15f1CjztZGiwb2ZLppkMzXuR9
OxF19jqF8gcetJ1bfCCAjPhb8F+DxoO34kQ6a0+uT6867M3tTywxfzu9Rebn
oWidpuiZgr2azP5rbqB46B3m4rqMuq/Jls2e/TvD42ztMS7fiy9v1dXowHbV
yozbC7l+jCVAmlJWbUIJ24s45JdV+BHkem6JydHRFF7jNiT6WdiD0UOpIa3b
Rp8mPS1zBCaVIWB/3K//RMr0IWhXglp+4ywZVkAu0uHzCHFEvpIyuVqfYrbV
GmKP3AkV+SW7Bo3SsLIpDn75kooSd+pglgJnX5yVChIY6XsW6B7MeWT/GO/C
IiSV70ECXXr7Gi7y0nNOkNDRvQrdPbrmeDBP2CSArSJQIiTkgJzrbo2fbiBQ
kCY01h6OkWV/eg8vCiHc1oZqLClitP0fuaFwlkspFGtDqs80hmd8vNj/rPmD
PUCJT/pTQ354hNj/twN0djZQ9e7CHpY0Im74ZXzW1XQcdL11gV5aHv5ByhQr
uxK7kkRnQgMicZ29ApEpv7lD/z8RopNjRKtcsUrVPAiCDwmIIsiYUH+7meWo
g5b0EogYmIjaM5Wrn9oULRlu54Zsf35ZunSkKVV4bCpEujIVwj/dSfxRFHGc
qXW0Sd5ywCd0OXxBysB6Ly8EtBYTz6CkTn62sfQxuTaAVsL+zZ77vEImyt7v
zSI+xj6HRp3m6/qYnITg7oAwT9WyfrsPzS+AYhv0zy3wYnW4/a6j+h0QlkeF
yQHm1LGzudV9BGhzADg2ClWhH0dVucnLtRQ58NJu7Zbul4xvIIMUUYPCbcNu
dSecQBZ/HS/hLOHmoa33Tc0J1VCf+3NEhEKAnQ2SipuQAEd+yPX/G46SV0TW
Jcc4DM/scBGjqWqJ+Dgl1I1Y3yE1ZYrQWXC4NmAY2qV3OSUYzfL0SylE/dk3
+ivjaZTTxCBdwXaGMDCAl+RDjXyEb61f4bpltC/In60LRxp9RC9hC2S83Oiw
z26CRh5K+vu9unAWwBaWtmHw5Jgz8bk6jAWMdwJA3g+dFKYO5XHLCECtZ2Qd
d5lc65uIoY945kqpIaJDFDa9r4Vxg2cq3vHtRNmI32vzhVe0zQz9Vg8hI327
ekxQlRK/A54MaOcxruEpDBzI1S7uJTa8RmyKWe72B2rmUgVj3x43Vg219s1S
o7ykiRxo77T5aEBvpxEp9UeFoq04czdR/0zdEJCGSTqwt2YeWRH3OK0FfgbQ
H1nBICQj5Ij8+82HsPl2OwkTNdjkv3PaKwF4GIoVbqgS40tV1JQUe+zgXBW5
NVx2jT+luoS5DPwWO2/NVBDasDNPYa8N86+54E1bQByGUcLinfsqicBjJy/s
xu/SuQIaRjgUhOSpM1qEgHRblcIPJ8Uzw08RcLS32I4XHhE/lweaUNNcAT1m
eUxkEFlWKubchUK7yq268Yp4GK8Q85Qi8kUrMUrnn/bsJ0D7WUh14GGrS+is
9+152Dx9Lf47ieI37bEXLf1oudLETuzIxdJiT94S/VmW4ypZxXhMUBZjAEmq
Votft2PqyjR4Ku34rKi1FH/rHZYfSAgLoC9fHuAkgDexIpES8nC+MQ80FUcT
DC03bVPVpHmSoAWVS/OH+edJ5WDgqJDJpyYf3Ak/0QbNX5biF8ucZA0STmRZ
Ukk9vFkdFgZJ33CqvYvyZ/CZpQTsWh3TCzgRibX+eE4vu6rey5YgUXbkTKLp
GulO+PbPzyWfvv9IJ08fiyrMKL07L4KWtShgFOox6GyqHlw1YEVRjbAk/bSF
ClZs6jpFGEX4sDT62fb0QDDdIAnRrVwGE7a8C0jv2J3cnKN01aMwCBwJM1eh
Qd9IcODcKtpDEpnagb+savQLsmWNrU8ybR/zgFOrpFTqEYF3sEZEQrtOXdh/
Jcyq6gljnNixXvJ7FT3FaHuPY/w5Vyq4LJyCYK1Ad2P5CNi6L1VFgKH2x/Ux
tuwxIMJQ2NWrvXVpuREqBJjhYWuc6ufhVFygJmMlRhh/ZBDYn/91tCD9+rgw
TQS25/9UzRwDAi1e6dX7YAYRwv2P2ftIf/JwxwcKzIertxiPq8rM3rDwYk8h
v/4ybUvfiRW8M/A5AxE44D27FL89NsTMdK5TgVJvM96DbOIg/AsFJeYHFJHq
bXCcyK3xdcoV0EO0DLfjGuG3kqqaBvlcV4UhGE8EMW77WVIsVinh6Rul3mbI
sJUxmxwxYbTtnUyDFUoqHFumCQ2Eg6rA3APj+Wq6Sal2OoUOpp6p2uHQO9Lp
OyfXuENO+ReCfqS5TOIJc6Q0RourNgz3xFCuEUyJctgaaB/MybvjWocn+dk8
MHUOoKQx3bdWj5CQW9duAfHgf34T5YG8OtmhMhsbdIxryLM6nfwajQXzg/lQ
s2DkXQZlfZc4XZOkbRXNJ7AG2PAW0wAgTZQ+cDxb+phu+0ZmJbnnayin5IAQ
KmCtYEQuQjwwwc2ZKqyIciZEF8iZCegffh6btCFsBU9weS0d/Lvsf1/v9npp
VlAd3nMvMj2ZGO6+ImjVy8I5gAvVwuMsiMuuPTinpHPUO+aCK0QvQ8cCZmnz
RdFZHG97ppiYKhFSQjyCx/Kh5ScIckqlCrWN1/CN7mqfQgcBmOcktwhQosU8
rrat0s7Ke+ljpppnGEefiAW2jErY66V3K3PDVSeTf61tqWK7x3a6mYpEa0oK
tICuGL9ODs+DpIiFJyM3A0O7ZR7I10szzC45jhsCUYA5nTfOEWvexwRp0Bf8
7ZzusdWWqt9a+s5ICKQwJ13KoPJMeV63e2X9rNRugG5M9gd4U5axKWMJolqJ
R+W2PtWBlWtjWhW8qMnyhEp11urJWoAu9k1fY8dqMoClSAqXTLOLBRjf+NT5
JSMVRojh1LmtrCBvk+o+zR+B7qfSNqwA0Na3z0ca2OU9A3UgzEWNFYDltbIR
lkYt5zro8Sk53ytQGQoqyrNtBVLfKIGSm1e2Ie1vB3872uvWraUXrceAGjPv
Z1mFiHkv9TojSVj0Smj9tDQQefio6HpO5Lj736Vcy/hR+KFixjnb2EFpyTcz
GZeSNpbr2hsLiLv7wfCGbU+Ya/DE69KKdE5h5QcVnkqglAum45GgT44QJDq+
G6uzylqKoysLWZ+8ooqsJg4/wCrPv9TA+Njb91IiIv5TAwcJq9s+/Zt5WU6K
iSMJD4Y+EicZfub1idNF0Pkh1901D8cHOLHda6UxVUwoTfk0lqJ0VhuZaESM
6Ilo1wyMSMkQIQ2oH1Egs5ZkbqUFYAigrJg7YOLXgkFa0vb8x0vVc/3W9WTB
NykXzHSPh17eXKPjk6ihtanc9GQI3HWY2/gemFU/D+sICKccadUoqP7Y8b6t
tjpAIzr4Tp0SHBbYFipSsUgXNg+eom/XUf5jtV1+nfPaE9cvXJLwJ5uPJic0
RtD6CtrGLzXTWO8RmruAZtyMpzF3BkM+iYwvnWhy7T7hZ9gkXqcLlBTytbQs
oYdayifKKtZ/DY2EoLy96qvcCcdTs+zy39HehRjdWWXMgoxXtGHXPS72/H+P
CG61/zWYh5ffNAb7m9mJY7Cn/hfU/229qqNuBIfgD2+UdA4S8PC49YdvNPAL
R291/8vjHuHsv9eSHbiaC4KC/g1k79PBkc22JBZzeQWgwoXt1T6fmtaEBzQo
IK3K7PFOK2WPK4zZrT2QBVS4i5L3CoJoBNBU27gw9wusmn+VkivRV8o7XC3M
k1YF13gGO0reoOgU7BFipUeQ1L08w20R5j+grE30zRWz6eYvjS2WtVj7S428
9KjuXVe8hZEs9/tUbaZIPKXKU/YVD0z71Dw9JVcqZbXzjDhwShjqLcazEtaq
9TOLgLCt2vY1TWADCVa1zJbCSBZ95HKkDoQlVFGQ1B/7aC+VvC9W4xYKM7gA
n3aQyamq9XYOKQMCIKAOeoHLtYGLMoBLzJsLeeA0P8fFhUkZtXd7GYdA3Bbh
2wgGyugxQGC2dPQMI4j5kL85+RcXA81KDjd4xrRva6/aSgbZIJfCqTuu7KFW
Sh5DinEGAtagK8hlAnlK+gRdGuU2RlKKmpTqUfmEARDjP4nQPRb0YSz4f/MS
6RpQ3PDBZgOaFFHj1XD35CS9qJhE3e0JlDoGS1lUfkABJ9rNFGfknTg0J/Uj
GeJ6FQ0HRr1QWgqJTz34eDzqqa49vK4G0k2XF4n1Lu7w4E+J6nHKdJBDgYie
HiGBf2sMZiaCuAsgGK5ZXQ8juFbjjgdu8WLpNnaK5B+pmjkjLlRDxu4zkvM0
LYu43xAdMdnechTx4Gpu+SzcMsU5Vsus3ecf2iXBWnYvseoV4wJHSsk5R/vX
gO4/9siN2mEOoxzVQSNJvuTiNbrX3AGwkUZuxGXm7fRspwbs13DGQmQ4GlkW
PyJNuL3bh//vIZzko+4NSs2irdLRutl3qv4esIC+JQ76W3P3FvvfjD0G+G45
z+SO8Z+4uP9iYPEwmWkirutjXrg4BEjgEbA5MifNYtOB0deliVucO1EwJxWV
WvWX5gPhLC1Efn92zdyeQBwZNXhxh8A0mvPwQit+EWRqjIQbCtCrjzxgAWD+
0JLWMfPbEh15tzv9l1vfeczqkgJhbU6wLznrB3Vw3EsVSTULWMp3lBtGcwOS
FsTRSpwuPSV0Ab/AYeQzH3HNe1LPCY3v8nKxcD7lY7Ug/44qQGZ9J39iHSbk
WuD30+3491756V9cgUzWlJjUHJ2aX6i2HkNoNClncAx5FglSNO3t+ebTBDnZ
a5Usji+y4jyRz3mzCh/Uo3wqUJyaNSYG6Zv6MT9xbW5w/wGoqfAUi/vFr7Ac
+9TIshWPP3Q653GIrfKs2GD+fyuH8Mup9sQt3tM/icW4+P9vXcjNuef/u7Ui
8KULDcpQHcHsl5ojp1T1CZAeMe1lr0NUrhJ83KZqviIEnvMY3pRLEiVh/bN3
qXv+qP3x3KAsJmFpjekHGmLO9OwZ6u/xVvoA0BYxqAUPN610soSQEqDjoZ+6
SUAzdl5z+7YoCEliKg1CnX04J4dLf/e+9mV8kUZzSh7CSM3HfvMpIieBGyYF
wtD/WJYDpomNGnaDOQzWCeI3sT6lrxwXIZCi4fkEgAZ7HrnHeS1Um+Z64xka
m+Rro17VPFHnNt5vEWf+NOsmden9LyFI87t5d/jA+b1TMcUE/IlsMsemqUbY
b7JDfX4VQGZDpIJWmul9lCfFM5r1CvgEoH9xNYKazpgye+eI3DGAAiyT98z8
sW1WzCh16kT/N2vOAADBfI3vN1irhCLmnbhgs4ACMQKh+ngKZwp+co2CiKD9
JMXOJAdGiRfmSh+rOOgIxzPrFip7N58s52j+xLYuVItSFXzyF9dkcLjqsffH
FHSDA/JT1ys9ai5hyw8+j1JPx3Ph0cBFsYtLuhetossTxVtMlOhwSFotNprZ
c/7oIUISa+1NNcUm1cS0ujwmU2L7FxUnHr7Z3m7MTyUjgOw32zT0UgrRmb77
0WiYHsPc6BbOjkaTrmpJAegI0BhGR29WFCIVJLKWvvOUF6raDzBkS8SHJnVm
Azrs5Lb1chyGt4eq0ywUSmhJJkeMTmaKuiQeoxPTqxd6r7uCap+GJ1AEqjrV
JhJKqnBBDU2hrIqHMLgwAG6ZttiS0JevUORky5WOf/X9YzbkQC/nVcuk+1z5
z3c5XVII3CPz+o6/7Q/2aF4sW/Btqt2Xo9aY8rSBBCb9LoKUvLwxT0Hzyhdb
mtKpUJx5r6XvEvR+IweqavAi8J06TFfa2x4V5IvfS5oknCMhzQSoiiuzG/YE
tjQhu4s7r8bkFFOsi4xAfEfe1sQxT4SgXcmYF6jygNdZR692vBpIolIvpsBz
OhueL3O+/Nf4ocF3KsiJZ3FPfMA9LsNwXyGy1IOSD3EQ134Eg1pLZzDKZenc
5TLTjWLJTqkXvA9gVcIHOxxlsTD1EHAXvWbVgrZE9wrmizqrO7FbSFqoSz1h
GHcZlvYPXT1eD2m2NmMs/RcQLwYAZnfdN19n28q95972cmpFWMDwBPzIiOBX
xMq+ds2oVYl91fQlIK5NWm8efxgHPAHz/KG5rZakT7yjQDbpX5hgEDVP/pFA
GjE0MnY39hxpVi/ENHLVwMZAAXPKbfN6Uj76GFuJObWP9i5/wXjplqz4rFo5
Cy9AvcmdPTwksqeKPiErMYKcUTEW2QvuTDb0eGVVcMlsZZYn6yBra3VmzsNZ
cGJJodDEkXIWhVS6kl+no1yFzgHpSEKRs/ZVOcqTqUhMbXbdL7c7M+wC9ZrL
WQZilX31rYTwyXciyZM0WWu1BNWIym/uSrJqvdoMEC8tE8IZYHpqg/ip1dAZ
qRGKh67YjYXUyqVTCaNKqfKB8PlYd6HEl811ajKNryurbmlSJuCmWkx4tkvU
u0yo5kJ/SJgUo0JFviilrfW2p1q4SV34pzTpl5S5lSj4EAs9oGR8REQLLbJS
qBe8H4YTEXL8oLKioADdjdut+zFnQlQrxDPku0oFw75nGS9xjOHKe53wPvP7
Rj8PkhZNzG482jWkAqp6KkFR6llZA2Qnm91DsAx0ysq5ombvZZJVvu9Ggti8
0DgRYIiyni1MDs2Zx7As0DwxlQFpzAOouJnh8avSkl1kBllji3H7NrAYmIQ8
ydpXC/dZdlbI9ZpVfe7/sEbQdMi75egbOIOJHr0rE5XhWq1HlvL6p5UqX8Jz
E4o7DpTxF2P7c1BmpbxDKWoy1qIb6U2pa4K2HI0gKemoOTshPlyrjdjAs9bv
ZTlqFAbev888ROiy1EV20qM9mmDuwzuHCi84aE2Uei6Gn2Hz54m8jfEH022B
b6gEnZssgGAUv3fjO+6+wz8+vt+EP85dfKmIdnGI/R2a227tEucCvRKjTBAQ
NeAWhvZujMPmRWD1R/RFbZZweSHe8ynLgzL5K+obSaLcJYbt4AfHeuu6DHF1
U0StRHwtkKCJYU83wxpk8a4eZstYXYNpZ2skumgap2rkY9ANJk79i2Lj97dJ
In7970dhGXdzFH17gBN3Wb1mfjIAaoV+C0hz/J4U3dZIstFwi2Gl/LzPDNGf
xTg0OZX4Hsh10VY093gXJq1OOWJ0TRiuAbeNAP1nzy1rBkb44jAwTYqKu81O
002aeV1IYcaTCw7Gk/zF1LWyfJleT39euy3AtfzZGjRYWGxFlvAJYw1AnQIo
N/68GmWwblvTYncwb+oY6gLeZgzBgaHCjeCwK2z3lBjuonYNKZqhNWQneG0z
z6TY7ueel7c2WWFGzFC8t6rusTCbsjCsMQ56bgruiUshWVU/izsrZs34/SGv
YkWlgm4z1GIuLvdu0YxETb3B7clkkZp3gngDQ7xAlvVELn7b7KjXOJuShxWq
ItZ8NA2mp/SoZTqzp2dzKGfz49W4Jsh1n2Qton4jWtl4xz27I324o0idMrl+
5xiekePjvtR1bKHCMRKqJkaCL0cvNTGuOZhQFb09ImxUbgkRMG0xYGKe+vkW
wN1qR8nKx3PXn5sml5qGIivRUqHXXAGr1Lw8r5aTWZNKgVX+D9lRUn195fTm
j6dW/0u4d799HskXk6w5vLPb26CMJbZ+8K013jPNnfC9fyI8WIXmXihBDint
yvxfUfEN0vZRw+3jwArgiYO93U5RsDgTmOEu5F8PPzV05GHEwDnVmkB46HMe
Y3cjXstlsKxNkCku9EATU6/2mzv7GpuISRHNoC66rNkMjEieNCNNQ1z0kYvD
kIrLCkoRKN02//xPXagDdRajaD06VhsB6lbrXH5OPTO3dHZ2msQGLgTmOmbB
FVcgvlGBKPnuLvw8g0GvwF84F5IHxbZAtxYUWPDk7Wf3O4F5B7C0bq8tnWa3
rw9hQTidx/e1SijWTWvNsvnSazUup4NAy+KpocddKU16m60bzUQMDxVQnM5U
PUn0XLcqSMMhrtmlPGcpACXSd5vxf8++DoC55Xm9NpcmdD2i4mB16HfshVot
18nob76IKOwfbsbbQ2q4ESPM3vCgCnrYM1e1HQTJhd25bxfN0R5qOjmhv09c
gPI1wNGGxu2MHfsrKcMd+9O/Uyb158GK4Eotp4JE4SExKMcwxr3z0cRyKIWZ
upOgmeoCbT73+noYkYTcdEEQxkC7xSIAXslZH+zgDm6lrS+C1dxf/mzMIEDL
HV8tI1FvN64+vlxx+Rv1yXjkY2iUecQ0AlsVTekLC8KOd8/4QZ+zK9uaegOc
WLQroJSpAjgDhhwQz8W8CS8YyfaJpv+QZASYypxaMiup7BvRLt1MxvSXDg7+
gezT3ZHqcbRWKDDcCeNrAEd+oVX7AwQjjFe08capFyO7aS9+jPkqSH0U4nFS
tg53SAoJZLUXcv6aMK3p0WLK+cDbA6hBKIlI0fXfGsvWLKYqagAPvLkQWjhp
49AesYwlF6myOSxvnBEuYyCeWOqglQFPQWNh4f1OgrFSGo8Htixp57Rr7Hr3
KQh3awrhFXB+zpz0HuatQpG+8f0rA0CVH/fQKtgLOkWUdQj8ms/GDiTVSxKb
jSL7XBpLqEUA5rNpqgEsd3MyylWzRXQOQflvfIIoH8JflUV3UssIV/ZoPV/4
VXonuem1Nqn1YV7H+0a2i9cgkcI6Zz/61eZXnwkR4glL2OcqsqWrw1vV0hC9
tL/BAuLS9PMuVQefdhJJLiri+YyvR9H4R8Toyi6MfH1g82IWQt6gwt6HkIx9
+ICx/6qeHKsikkVevKk3sKDz0JYw7OieUTpSNpNoOBarFJ91jFkexNTF8TYv
czi8f8MJcFcvkA6g8ZtDv0znpsglrcrrgKHrgF/515a8vPpt9e3uf0fzbnbj
DyxGO23QqvBFmxw4En2a4LEsDOXjfglk11GgZuODTDskQ7xltfbic+mY/tly
axxW1/NgqXr1ttU1OXnNfg/SVy5FsWlBr27pJM/Ni9Mn9tSgzSyDXkxtolIC
KNuGXNwxWwhMykKZ1Bc275RgURycKYHmR5ef4Mpsws7JlVwrdfX1LFsIsyxb
U+v39QXsdcJAEhnItmjSSKeEZWN7MeD8w2P1aiOdUvf8q/9D4jSncC5c2T9d
JHBnZRKViDnwUlhOGSIlt7qA8abpAYLqDsQT9WL3ii78un3jPGxHjmCH+yK5
M62d1utBSG08oO6bCrZKPUwWksoLquqILvEMH4oVPxvDpbuDAKnnj2PB+9Sn
spU6t5dXr2WhSnmXIHIO2Yzh9lPeXA9JHQafQ2MCB7crxqw/xbxD7ECnXENF
8cFWLxh5yMbo+TE09uTunMvAtJWdWTTLH83lz2F0OcS2fo7m+u9PwJknA+wt
kqgjyEO/v7To8y+wiNqLyfmOfTCXj76O/xt3DgcyaS2qzHfV9JWdzgU1qd1J
h7BtJsQ+Uvzg4ODsVif6FGC30pw4aF+cKl0L6cgW0ZWh1R5wTkMp1asROtVs
uToiWacnLhSeMF6KvnZDwlWuCLSdxmiAjLJloAzCcN3F6NPCyT6IaKH3q2f8
KnD+BscO6EsfdS2/dUpwvbXTO/E1d+3+3Of3l3YSdPfes5Z9jvziFFrVOFy6
iHnWVgskYJgSXR3e2yV22Y3h71RZQdRa++zgISkr2GcXl5BED9kINOImuMBn
Sn2PL4pCuX8s8wWLiECPPxKoWsglvm9NGDiqzMQyOYF3MUAb1fZChR31AjVg
/HtQ2I/fCthG1jaMTLTWth+zLX7T/83BKC1TZYMfjgVEauABf8rriHgjZtvp
wyjhErX+q8EaQtNxOrfgdT/w86oVRf5dsvEf3pgBj38nbQvtIjjPrHQi1hnC
Q70FzAqMEiH3nmzB3rDHUae+KkNan0CV6RBwkGMIKHl5qnTVLM/zYPY4xjf9
1ZY9CgtGrwfCZLA4GSjjIGJMBYQCQznANmH12E41JAzDXW7j/PBMBRS7GtHK
wI1sYQSwiyd1txhw3Zg3mFVHR5xSBSlOmg84R0haC/8g6Lce1nUrSw/unnlm
Q7QZN0wT9NiFnwaUUSF+P9ybiXFVMA4/QatbugBo1LF46/BmF9P4EFAHKh7s
u1k33BnGHyXnkxS4cOSdI0j8A3eoX1xN0DE05KphdmL/CW/tvsxTELSALp6P
l2TbyKOIPwOwrqE9IUwedyqCX5M4Pqay6vjWpk+zVrDJFGEOvhKyyUSePnnF
dJN1fLO8bzSYhuemL5THF/lzKIA8WgV7nneP/rEuvOHjCb0QsjIGswHF4poY
Uava8RhmZSFYSufBmuTT/6HzBVzTLqw8hf+uVOtajs4U0/3JrfEr9Y4qzMJ7
jUlONoDaJG6KkJIoNdG3dUMm1ML0yqW8KA+pcodYJoutDB+WWVCPiOFlWFdF
1JaSqeZPXMtAvcITM9SvxiOrW1LA9FQgOIhlo6oxxkZE2EDdJQsvw88e94QB
+VQZy24HqqYiq5u7ODsR8uTSa6XcVdl760bUDOeNWMH5/9O0/ER2HO8eK5qb
1klNgoVA4oPwBc8UxkFVAIkhe3ER4MP3WTsxy7bxWwvaxy1vGR8oiJq4iRfx
jKhfYVNQcgJ0E9OAxAphbF9DznTbQgLuG+PL6DYHbymEZHhONmkBHmUO2ITN
V2Y1I9Sm4yoa12F2o5n5O50dL2TkDvjlyDEyb0dQOLZMeVMqd+Q+B13Ca/G0
dUDDdvfBOtz1C7JyW/XVbAmDc2iWm/mD1VSMmntgrlqrlkKT4O69FLXv14oU
PzbUmCCVweCMT2vm4vVVnbw90I6dhvkdEreB/OLI+KWTPTDq5NqKKqSf0+Mv
DBNcZqvudwFzuFXj0IA5N/rTJcJW8ZUnJQu1sgU5LdzkCG6PJ8hfSkztSK92
9Mhq3mKEK9kt6ZsDTy1ft9HeWNJWpsuVySpSmof27I+4VTOtTysgUWBiT999
C9toUvd28nRczfAkuxJFMhyZ/0p9PPPIv2VRDQWaPgWnYseKwa8saj6uUxaB
A2E1lI8XIEFUYPRTKSRogMTLz/HsMVb07CSvg4B2nqw+2cDYOsG3Nt2qjIJO
gLqbFE3Bb6JJKVrbsKMtqOiESu5HDvxOaJzDxRvqkWDvxZ6J+Mb96bd8ql8f
2m82LgHWIwqcBZwku6ZgMgKxqZ2jmIA9yo7tlDEPP5h8BUJXrlk6JTDc1HKG
lnuyWbjsZoF1y8B0Z2bW7qfOkp2y9QfGIvWpviFnapiDxDzCCPHmOdedW7vg
8yBzK4KxxlC6cPrFrqb9QjDglfGRViW4QxR9FTKeH7ioYLGCN9py4p2/BZ0X
ZYOKk94S0iKx99B2XKmorI2PI/Bq8psnzJW/A4BnT/S2R8qjFJqZTP5BA9Or
V9CT1BVPMb5MKo4y/vJiHGyiq47+b8015aGRb8+qXFJUx/tvH1wZ5k0Shaiq
Fif792PnpCCtthQNTdJS7sZpwsQhlDMojnga6Qsgd63zMOVrRCsPJJpR8zMb
qqI7MHIHkKdWMBsIsExvkzIBjf8Q5zWaSHa5nRjSe1k18nodFEPtL3lbSFuC
+TIPhSc7z1ndoWjgU/ndsT7cc2bcvleXTG+Q/ZjL3V1F+KIod/ZQiRZnc+Fj
KNUUoSsEadKW1b71xN7nzkJMgc8bETQ/6XwLnp3GaJd5dFPABWfE6SNdu3ue
DaNzNhjQm8wlVE8ibsyEeeKz3gSeUEaO9TkycnBGxtzeFeoIP6+X7PaeOIr/
hM8yee8rajuj9GqpWb37WGen3yHoF7q3KTuh14zWYd8KNxl3iDVrdGtmTD78
OqzRnhMntDRnJBT9lxNt9QMtDCUaWjJR26KO4wEWfgQzzHUph+wRs0xbcJR2
FQucmNvbAUEsmST6+H2crL+6fi/4vf69uhZO7q198n1GLt80PeT9uYM69UHl
7pdzL1sD/TP8pZO+oYzu+K2E4TyM/pVM6lOlmft7DMVuoFoBUc/XX+CVB6mW
oQTSng+VuKJ8QQhp7HaSD2wzG01eoHtKu5P6XgPTC44/Ag9/7c/0aXdvs/VY
kOscBV/TLT4WrGcC5/qlNM6eMqsum0JWdCo3g2JXylyukobCnGLmM9SbZDEG
ZfIh6EWQCyeqtY/UzxmvIIaARq4VAL5HGI0LInbWThT3Syy7MtSeEYVPqvNG
4AxvQJT6NmtedZ4Eu1na0MGXwSHBZAaaT16IW8dpeNLXW3Z3UbtAXIxrIyoU
qLdVtf1gvAPiRaRH9RpVtcEVNJJ99mlrFItBJP/f3UfA7bHb+Bp4r9ekAvD3
H9hc5a10WI/btAHRVWs14gxcXSqT15MqH8o+MHPoydUbiEqfv+gEjlZWtUdc
oaxcHTiPAJVbVGlko+EH/fTbFc5y7bYiZK+U/WUYHyaSh6EQmG4lkdXn/UAD
X0Aa/XoD5gMK5pk9hR1h0XWkXEkBBlRG94GHNUS3mVGWIcI6jRENrx/QqHuU
SB2jgQvbdwVKTzNFQbKs0XX9KwYf+Dy2zmkvzsGwielc1yB1kZ0eY5349T/U
I3eMstMQZxDfUUJai18ZpZlGz7P8L+d/nzw/cByYNTQ7eyg7X6S2xH+ykcHM
EhL+lQxd44uak7jTaDodQ7RZcwyh3h5kkDCtFP/tDzvLttKf8smPOYn6LGgN
vS/EQISfHWyG9Iv+aq5DP9l9jZtjtBPmny1wswnI3mKnoKXWHJ/GKcm3jJdZ
4YNB59V0BZ79mmEucTiH1v0cU6QoXlrZW2N9J44jepTzzfOnNV5cizMMQmkc
AGDhHwVEqdgsAheelUg9ayCewZEfpKs+RYeReB2cBY9rUyTjV6/bF2Shaanq
TuuBem0G1SlE8AArv1DZ7R73/aYDEbFJ4EZ83rk7LFXJhnPapACTg+SrAbQp
mApgT+74bObgcByiJYrA9brcMF857sRoghqOlIfgouXfTmHVdYlWAzJC2ArL
i1ELUm96dxQn+76Za/7ZNFV4cKjzc1V0uk6iDE7uNFy3IlyyW4jZswYab7jC
W0MTXHnklF2SyZ3R7b4JpV1FZPq+j+s6QifJTduBzPG4IIT4DHJMMw5LmDU4
BI28ILzxqoBrlymJGBt6yde2wwLqGtzq7TArycQsIBl0Z5BDoX+sdwq/l3xq
3TJsiswK+XMgfC/u3FZdRj0gOgxSKMPW8u70mZ2kSCiET2d0blDKCy8Z4HC+
FUvkWhcT9dpsLAAh9U+DXOkBEYC8DSUiQfDklXtoMaCDAs3NV2iW9l2G8iIo
a/dCPAV9bySby1E5kxpZe8gRQ0FPiDY3idZXu+XIXSeu5l2qddRcQduO18a1
/Ceji08L51SJigvhY1PkzoF50mgkfxE4R1dPBTROS9598jlm43yF1b+hDMqJ
66IC/jDin/OWLbmXSjH736eGI96HxkC44tJcgijUV2XwkQ3AB4W3xsNGGTao
LdyygjJVOf8/OcXzM9euLByzGBL9FqLO412JoLg7FwXkOpVkH5WeiVzh6Siq
gAx1uSQ3+Iu1OFLoi4IETfY1W1xtdDmb50lmS7pLoQOryBOrZV3qAETk+FVx
hkp6spwbMVRObNYmJKQDiC+pAqyjvGYnrBKlSjg1H18sL/okZ0xr50tRyuv/
q8XOnyTjXEvweQm5XHIbKvQT0aLts9V7QQ07N+rawzfdXaiV3gYuVgo2N6GW
2v4QYQic/3MMXx/r7B/B5eq40pPqKbaTKyrzWgKXlWKTH11vpA/FJtuIc1xe
zBVVgksNuDj0ydMzXiEkOFV7mHmk625W9RB5MVORSSqLa0zfKe3m2X2cS+wn
nVFyLTr37oR+TPqjm4gp+v+j7eO5Uh2fbFHIGCEauXanHeDNZSToOPcjXQUO
1joew2yUKUOP/Q3eBYtuxLkCFJO6WAqxfvTWX2zUn46Q18x2BerZFx7h9nZn
IMAklAZv++JLSdc1sk3u3j3ssoKiqo5idKIE5SpAavnPpBDAe/54d1inHGIb
2UQ7lDcNx5SuRW4m5JJseyVpW5/Xdz2dP0eE3FNK+z0i4a7GFJEgGPq8FqBc
+C8DIeClhxJDcvdPY2y+uKGS9A+LoboxEz5pWkX5TuSp0j27BE2dYX8padGz
xf7SL5/+Uclo0g1o63fqOQAIqKHlJb5DbwIZPIJ3vU8rl+HewF9854hcJwlQ
gNRFUmAhx5Ptfre00vDC1QPrMtk0Mix0zdf1sLBHmWJ2gB96Pi1i27gvEvcm
7IhToez/83EFn37gSUhmk3G8eVRys6Vdl66PHqWPrQq2h6IdS0BJANXdgEMR
7pFTKUsvo18l4sUuxRWgP1JlMqsRIScRwvLpHAWTvYWdvbeFJkYbxMDIE7vS
ij6WlUvcCL7NEz9uiV8apUNALbx8yBdVejB+VFJN2k3PcSZMaBws4gtEMzkY
Jk+g/8P6XK1GAT15QQ5ZfmPPnHrjfFGNVZAt2qlMyG1/H1TKkeIIrMRduWDY
ZrWFppdPYkUR+Q2z54ecorbNrs4abZjkuvEKs33OTg11JnA/LdI52N+OZbxJ
As43w6nH3kHW9iwhTgKZfMlWuho4a1TsQ1gbjS5FXynIEvDaU4tgNt2gGpsW
e/1eK7BsPgzT1xqkJNKy5cr0quCE2Jf+OP57l6cwkbLao9w6n0tV310s1Axe
ryTBO2s+GMcbZRPMnEG9HD7BwfIS2/DBP/5VkZQP+0XRm8iDGdvZESE5Eqjg
BFmY5RdftfXZnWGhbd/u7MtAMko5Iypn/i550yEEw41cRzi8C9meQu2WJrgC
7kGomV5kaKTjp5K+qRAnCsXDuMn2fEsJxVtL7DHTq56VTDQFVkhZ2CLMP2qG
R1OJjAY3ymVUB52lN9nCyKzGa89mfNPiVazTciUY3c/s1URP7nKsrHHKgInJ
5RQiFWsPZpi19r5ppjp+myd5qLS2hhrB2NWQ6/QYdvHGmH6GUBhrUJA8M96j
BV3O2HDLDQNLfIz3e+wZYrUF4ScIxY+Q9Y4lvsqAxNdTIb7yWnRL0MGhDhAz
/CQ2dsuhoEzcLPSwpy6j46wF2CInmfsV4cUMT4JzohKTMyuRRq/9OOv6PQv5
StFRd51u62TB4ZSTBO66NIhrFh8Ehj4bhJkjvNyJNnhfNcHkgRu7LK19lJtR
5fqyYDrz+ks1l9HSpCNEMK80TsrERuh/efQDUzvc7zLcflAJFgBZiXvegA4v
UnAtIAdC2NN7f0+JEYplvlUq4/L+H18rxhnqqimE+ZuMindkhzrz3S8+9sVE
MUpT72ax+CYkLbJZkC3FoVJWsmwlxno3wzlBi+8wBNvLlmTRa3xYG+bkrpiU
e7YhevBxRJhd7YlFakYOtvTLPAbLLsFJibRoc58a0630bQludBsZLSME6VoU
UMy5bde19D92K6B4ZFBTPLryGXYaVLuBEUJgZxWYltjiX2Q8eNFqrlAcydOS
u08zulfpnqRJMayVAOTANeU2wv8TzUg5U26mGyJgF2eQDp1Yo9wSCmNbN/nP
r2X9BdoE3wFKJfkHhXarwDNdkaj1k4KqWZ2B9ISo3IKGhpoYosmZgTA9EcgQ
xgMakMiNaE+gVAXsXRhicJbRZnuKYrx8kTBwn6MEg7kfM/2YGPlKjnphdQOC
hCx2crP9KeCiLU2VQ4FnhiqsrQeSP5JoDel+ohOoR0kH8SWHLOo6OWRKL7zC
hAZt/5nJv9HHJZ6jS9GseFIOEzn4hMN2nQTlrDjPKYxpbCPCFi9RpY38zi4A
URPGiTbn3VJ3X3Czv+l2MYA6X/wDND184LXWd5VVhF/nFbJLSp98xZ7HXhDx
IP3gupjoXuxT/0JHXTUFNUZjA5HmzyeTkZI6xNCVa3z93mcBg28YC2ET91In
0W+zFS+qM+a4Jt3FCo7Clx7ZtWqLdRi7fhudhRvMxNsRtCPtqtj2ATvw0p/d
54zb6pEEvkOuaKS8Tj7kbVVMBEXSOMj5y9ia5u0+eC1nemzHjLqUeJba219k
P+fVPfLpsiKNvabH+N9SKZSalykx6WkZ7l6j/WMYIiK8v7utHVKI03FQCmRw
mc3PpbSb8Ts2teELLkIW8O7lbHh1CfyL0MTFTftq0o7nnMxc/lo84fP/8GvA
e5BJLKE1/sLxnWJJEPEmmk+8EJmvXw1Tj5mEPttAq/8GClnOd5wRO0BGPPL/
AlSiUubRUiQsd6IQElKoR5+0QP21dBlcFPb7RPhOF4kj4PwNGItvb6iSlfBz
IiUYUVoULZuLLr1Os6k7NjPwRTZXiDLd80rGkH+VtjZAcJj5qI+HKHN8lBIF
LKKZmLpQ7g1shvBwwftoZqR1GES5lSGOLFdsTktDzc/BDP6+MQiLsm4DNqhB
ssE2VT2l8iLFjyD0PQJiSSvXWquxJXiyCJPTxe3tv4aQp6rG4zZrv4fr+Teo
Akssn69ZrHqIL5gqDPWG9S9qUmdCBnk8RnPXSitBMzJTqxa8X84POJJrvDZ2
3RXHDgKt3xNwVn6B73C65XlOTqOaBiC7gIPvWaoXhsg5TgTIOGFKZrZrKejS
YP3qe5oxRCrajpWfQaqH9yZOcGdr+awrhdQtOiPgALl2q//n5/daK2eqWd3v
TRDwwHzYK8tRWwfmdvksU4gxenG5RLgYWn1x3o9ZqqWlif/mi252jOWrLtMU
vrwEmyixIMWYiGIEr6LgQPxXMj1u6b0KhsvZaUbxhfj1F8crgedp8FQa3kK5
UhMSEpdLLPVNFdFOVS0uKEd27H6TD1xQ9eMxqtNTGRm0zVYa84m6WKxxiumL
tw4ioPx1QSP3pJVUcW8PI80xTNwT9wtFGIRwYyf/iswRGLWEjhQxrVM1NFVJ
DNsSywvOGemJqKYIQ5gE9y2dFwInRE6puWIiY35JAvUq4QBK0YOqrofDRjC8
9HIDDLPJ1tw6YCMrQK0B46sgrCLk3ULOX/fAUKhbYhr5/02j4tPfuvyOJqds
0cu9gjSxVdyCpTEsPvfjCXFRyHJs0k2fGcblDjQeXGd+lG+I9KnsHLWFJWnI
d2LdPcWRgeyMqdRhqvRT9sbsM9fXgOy5gmFLXIerFxAgvSbxO4VAe1Xb00zv
yQ7fgBiZnIIoskR2B4KHsrmqfW5/cag2GCbR2RfydajkgNAQxMAAwhwvKhai
QsDBfOE/nWFPlbHs9vzLnLN2NAkb8mC0/rt3aINifITJzELPsiEJ3QmCUvbo
nIVDOsffT5ZMlA5yMruJtXC2pn59qfpXhAV5ecJsDaMsBTVz8LxHg5U1rWHJ
Y0Q367GnZBRAqbpAtwjRuQVE+gFVmPgTRoR8Cd5daoNTIbRIEs2TMRzZ+Stv
Bl7LBwnbNjNkGrwz0PbGRLl5z+wD/RZX+EcGc5eZwdQrF6hNpMYSTnDgEKKB
e3L4Fu9YtJwg/oakLR8VF4F9/TRayzpXWGWhv0NyeWpFrOPT7jdBGtECyNlN
ak+Oox+fICX7GvCMRSEHeMNSvsh11WuPIPV7K1n3fvkXqh6kk0m8xRt/ZPUT
ywM2E09LFSwUtQhJTHeLrHJZSzs8YmClLPF9K8SAgHnro8GsAv3SICsDPo5M
6yE1IKKJUdTm50ZtwvH5uLqZd+a88QJADwJEazCAoIIvw5beNBDkOPg09tED
7TrtRn/x1VGlGVIpMllIrTgxPWPJBAGFBfCccxG+iEWvd34v/YyIhumx0zkA
BXYk3CkTGpOQErG5nY97ziI5ZVbjnjIAfyPnHpMNghiyIP/quu0k5/Vnv4vv
UBgpSqWfEELz+SbEqPgi8XCtmChsfmnuJJ77iSe9Dn/ktAqSSsvK+5IxI5xR
T2szS9ZsgzUDy9sD8kjSCUWrB2C3tZliz7dLfOe47EFROLOGEoH+Y6gCTqIP
vZzL38FSLA5ejIYHeidv/Mv8kRjGjNUV7tGI1DhHeUc+SH9LmWfAawG4Q3YO
vRuXYkKb3WGvhFT+12eT5jfE1UEaOq3uDD4uYPkGdCKurX+NTn5NEHG4yAaq
0uqLoeG+NlxrBHKWDLC3gROBLWQaLmY2G2DwgjD+DmcUaw9JOahJFNQbt+BV
ewINIcJCfGHS8fvesMmJm7pYg/GuqLXYxbSa+DE2H+lV9AdgUU+tDkRVVQHz
iu6/JMv3Ls68wRHuUsBWu7hie/J5vjtcf/mFW/cPWxuyWjMTEE4+/yrNkcOt
hWmjwZsFjqFuiZ8pU0WBDvvYLp2hI36x1RgJD/ZlY2Y/f6ne+KiWILMuHae8
iRt4Eoiv/ZEzzTTtwIka4385kk8463lgU6CYjtgz+vDnAG8FqVFxuQJhyRO9
OggSF+b5+PuHSaD3U4SD/YrAoMBUAdgsBYwgVHassflpN+6o34D4Cnw+52a7
J0hCuRacNZTuDqFgXL67wX7oromEA96JxMvKhcm/YweCZLK0FH4LjKnYPdv8
7VGWA68WgCWYby+vTj8fGWkCObJuxHLqLQm1B8KSEZODpHzlDGOWDuaDFXfi
jDdQMbS2KzX6/iVDqVlms/oD9SedYNpzegErC2QuvCCYDta3rdClgqJYVqhS
vjVHHo034w7Ujp/ls77GpRfdab0ZwEIa0G5hWwiuIdLku8FtbTV+gvJSeLEn
z41XgTbxIuzgCNijEltwven8ETILCn4NBH5fPiwhK/+CKHq8G7CyglzV9PAd
o106KdFEg57JxvdppPXhdgScIPYfUqD4nduODyNG6CVMGrts9iZgkLtOuZ3B
wSc+XuZruV2cfNsfLg99oj6QXURw2n05+olYmI4IDd0tP2Elnhc86o3bI93I
XSwOF0Y+mgdYr+s58Yhid/dWTiSKzp+IVAjbz3cV7N9hzciKv99t3y3V6eda
/XoIQn8ZU0YWpEnX9Q5HIIglk31zhyIngGKlT/x+ESHYCYtMVXPJ5/1zPHvV
5GGg4+STcQTeXX/3CmCVUGA9aeARBfnZDVzwIQpQwchQkQVMniP1jAcILfUg
bHWBI0qkL/AQSj3ts44LH+STSH+KhW75RpbhXFy2ho5EK+1oYx3BdYCqYXan
TU00tA5Jx0fnvo+b3R5m+Vs0tzj0duCcpbPUR8Zm1PmTvQOkwAELv0xZ3YNe
t3YQeLT16UrhB7cGgTHPwiX7tzuYf4LmRoBf8o6mB5lEePH00DDfYNGEaz55
kCgzc5N9HP1uxyELFk3K/m7j530qi6JX62dxCGKY8I6hEullnYtpZFvHdOo0
IKxKK8QR3OAlkbA58RASHcovxu76FrUqu7eg0IlQIVk2A+OrFCgI1HlcUbQs
3ybffDfm7bLvTSsQy4GQk9Yv7MaUq1n3codo+zw3VZIEmgprsJQccZ+PCZC0
SVOnnfFi8d8J8Pl3ucZpaJCQ3e0R+SGyi0scW1hdQtg6DmMuAeMIYVROc1Q6
CalxLbQ2os5/xbh5w4mN3NQcHSXhUOB1hDsRuQJZYU+5jCv/SDaqNtCkMBU4
V6ED3Rhs1dHBB+IejQSa9K8W/MXlSWdsTVN1j3aY3rtZhuDWvPAvVVlNj0qp
uG9t1ZVuwJJ26bH0kNuY2S8GdJPziXqs6KRf9BXxotRSkUN8aa1phBpTvvcb
gubBw7mf275BchiuXEWjS5Go27+6Q5cV8ShVbQ6TE0BYSMXUhsEYpiBl5ZAR
MIJJx5zjBzoVvcehNlTePsMsONpI2QzHV4JY/4FhR9Hfm19S3D9ZmHIA5lOh
vuyaIPyQJNJ41+sPzbACZBTl1qAo6lCiwmJOx9OuOJicUVuozxZL3TB1Kreu
PLfGKlCoSr3nP6XAF9fOGioRPPAHauLOuR4N5Wm2D+NmlbkAyXGjvnnyH2nD
BhFm1oT40pIh4GvzrfaYCoroxU07iPdNRonFSic5Q+81TaG9L5E/eKSvw8bZ
WymExpJifkd2nTxZXtFuaFEPKf79woEnPmMa0Ou2CtYLYjq/xq+1rsRqp1dS
sO/cdgcKILOPybQSkv3hZBW9O5qWGkLyR1BG8t3kB9MVyakeFkRpWqQSz9Wj
n44WFvuPw/4y5fCrid4ioKJIG+NTqeEoQz44J5/U+zuK66WQp3kb3s3q0IvS
ARrLbqcgsw7NOSYgbjh5hXHcZCBYuIhCrQ7yf8f7kwE5axQpOxhc+KI6R2ZD
wSD2+77EZue70yJIHDl0EPKwj8/rmAf6YbnN3LovfL5GpeTNUDIS56WZZdia
zDqfbiYm0qr4/MZuUBzoHnSz9DlgkZWZEbuCfmm/kM2zd6xKlZgcVC5wscXr
6W7+pOgM/r7hlB2JHvHjy0phADTUinh3tdpQO7O9w5w1ybIPAv+SlDPuIvkG
4I1j2AHMchT3Waou+jYJ6o8QOTVqXkMI6BmdZ8SL/N54aJYnfU62jLGg+7e6
RKfwHLkf2lihnH2psKWTwBszXf4TKwkd3mpDGbP05kyVofwj7Ok2NZWH4lvb
xD4uymBN+vSZSGLzv0Q7AbQRD8cc4CrcdGzcmooGCvhB8YaebsOcsqMqt2uK
TezIHSCJvKM8XN0WCCPZV5GRwLSjsuPgjReQ+TLps/0scS9EshhTMxhG2Iyf
hAb0CJyaAI6YUF2mDviGEGAK+T+CBfwujy9U1G19jplFN0MVCP83D/dqWm6H
sC3HMdIESXA9s8e4BsNoJZjKmBXtML6q2i5MFXnsmpv3YdH+esvZzTwE0Hs0
4b8pbo/jqEXAxUAwanQJ8DuLor8ZGh6J66YYNQISI/aPfnf0jlnpwPU/k3yU
O6LDKQIhhXD+xPSwt0OSJowM40mJ6vcHhwq/zQCfw28QYT8p4vIIU+OUrSxg
vODyDH3SBmugbu5CiyrIq27Nl6qJcg56C495TeKuQmsKnMfIBz4iBl+iGzKE
6FjFVG9R7ZRZkgrOy7JMSsNNG+IRb0SDYELeHfv0BjtbG6b27cB9c96jqTBV
VCERwzaLkd3s3LriUnk/CFoMNsr6eL6x/gwMXBjqRhE8DiUl15WAfMtBsgER
GSymKdm/b/Cqz6Ei04Ix3ek772CwESTauBMIKTqTc9hHvUxYnsa1mQgaEPj1
LAVZa5U+pAVuCi2v0GZ9XVi+K6SAcADupPxnd9x7SV3hIa8hyzXPki2O4zgS
EriouHx2UcIY83mszdT7TisrUK2fOO4HgY+KukbgwCYygish8E2+JJSRhWj/
jv38GOdZdGagcWBIOpXW3uZbaPykGvSeNJlMdARjlyE9KmOgx2PX1rcaYrSH
HVPZ8uw5TclSjzDDrapyjvMIHF4Be6JXblQ3SkzP+w29XdJgWmdn+XEajISO
evN/XzHozY8xn4on4tr7VTZM3ocr5h/j4cU7dQi6OAtJCGgT3kR/NaJD/Efu
jvT4xUMWJWgSPfbnUx69L5KY5+gE0sBKtvBvey5eiOp7IpY9RJITu0+jsySX
Exxim/Q/XYO4OIUfLdvx7+LcdvgRiKvthRZoN3Vmd2nZISfI9cEPP1Uufi6E
9hOsBKGAt/i7dZGYgZGrebAx1N7FtCHnj3aSNRY1+vdB7V/LqPxcqZtOvM1m
0QaaG6nhsdBZVUFYxEvSHqIRwv4ow8RiFLxbaspKURXF/MZhFdP0JGNdgP05
akRX4lmoji8m3+aCsCKvSNE58+dtlRRLFs9oTCKtTKnG0HhAkhC1MVy6eU7N
nWqN02K/udim7kZ46HNwsG5Ps9k9jGPg2xirYZHborUtOYHGxgBVG++acg3I
vDqiOM8IY3oh1btsCCSjONEEIH2HGxInZpn58EVIqmolil66HKtYl1xTViUN
lNoQKgTAQbhT79U7nB6EL5OuhzskzpYPDrNOKynmq9aXjquC0f0CkuCqUA4S
9kY4F/ndJFEAUobZdN0A771PUouGY1or9XyCgq1flwT6g7tsAKSu/AcCdpSP
wfnJV5ke9r4GON8T2KbrxBqFoPMPEVGM1FxpI/RmWvYvwZ0dJHWbsh/fknOq
N6bMwDlvcjMSH1zC+SLlvTnXIjbZ6oZUYY2U2aaY8t/pf/nhwG+5PrsfEY+E
up1RhuN6//QHlXHyWfK/OKU98TGJ3KZXBD2MCtNmaYlZ2iVUwuXmCnPtUMeD
GtTfv6H5tigriGzewLENF09AHoHkJi8R++2poNjZYayXWpwb2t9T5cOwg5dI
iL/m3qOckbeXOtGubjQv1kjrtMR9Vz7PnEly2gXd9THIUvidHVeGxKWHpMq6
Yqo7FxR8XBvNYOKS9oFcuEFq/GPSbujcl77hOE2suKtxW4RtTenUhftY+39w
VqUY2zkjLe0AklymB8nuThGQ/ujlmVbDBv/3HcmJRJoD38MY6+yvOEq17yco
I5ViGVTiKXo++tnGrxvFEAAUQBsUTEHYNFLFtPqyF8OzNjGw9UzsdrbUjzu1
RtGpqx5NZP2RkCHBx2l/xQeMZZ6LNTXQ7fqddTY2Tg8aUGYG9FqK0PBlqxwH
odyzTphBXhX2mUzoRhJN0obkTOtl618UxnmYeysYl5XKHLqGvZ+Id1Ft/IWg
FYYhItMPuHJuzAqelR5t1yO2G373VV4VHLqg/ugPoKd2K1yse54f8kGvG4Sd
DLEllYikcMlMJ0/Ie5hQQLvtj4wCHt59fjQRvrtvSkvqBpmihXKufw/ApCRu
r9gdYL/e+AOenn2DGFWqN6HSEmDHatg0i+5fftAxFKPwUYeLUIX3R2g3qEoz
YsqeVVYVdOzYOyefOJjtHsRNmTR6Es3J0VT5YCbMossc8z63yJQf/bZ4YHYH
LkUqxb5307YBifxxNu5jqRi6+iyQx/2G11BL0iv++zK1uiVEtdErzlPzry/u
f4CLyY707L4hDlpjqmKhgLBgL3gxXvD8GgwEvjTW8UMP89Mwp/K8pepAl2K4
HRa89pBV1TvH++qdXx6qhqMPwX7vYBiBqP+NAc/GkTBpaCKZfavVENc0rN4j
SySQldMGi3xkwr9RRXbmS+xhBXHoon7cKg0GGihUdegKY4Op9KN1H1oHo2Rv
tBos1ICVQd5PxjhZnzinKF8/jF7791hlAxN8jiPz59ZVMQgdRR7SaM910ivH
oqtydwxotovjr1DSC+nUpYOcdJhNVXgUTe8GKC4RRv8to3uEsV4cB2SUqRO5
50MEdTB/dYyqdrTP7Wmq2GhnEm8Q4n4aPgxm95nqW8uXoU4LlH3baz0ZI5oj
ksgkmuTNUZZsLNyjztpoUrmRjC24E26bOLhIVSXjNv93ru3PB1920aFaj7fI
nkYUR1livQfjyMAdjD3MXJsg4LTs3rtie61iFfaRquvdzAVBjffS/d+wxNXx
MVgYCnvuZiVdBLxe+xJbzWPqd1uhFtoDYN3/XmiUYLidseLzK118MR3Hgqw2
PbeszIL3WgZEZMB6e+SneGvo3M8nC1VU6eum2p5EV4zxc0LtnD63BxmK9/S9
mhVkTKfN4fan8YULSEtTPfA2TBn/oiTCIntGMv0Jg9G0P4ttB0w4bZ20Aag0
Gwg50GZSCxS+1B4pz0FnyAgxjcXWLAB1bie3Z3yranAS3ngeqaZwMuR5huhv
EmeMeGe0LSh/tNdlVQyNzqnJwc4tuQUm0dMn/JKIssNJ6A+qB4MhV6Cah8cL
OyKECT0KXZcRKoOUBUkCxKWsu/FuJxX54KkVU+U9CePTEXXTb27sXkwtehtw
zmSYeCHONiChi4YKa8+SGOGskkqksQoz8/dyadhBp8pHQ4sjDqB3f9AWsJ3i
n0R6AOeqdeeJ601C6Wv/799HkHcs/4ZfChedxnI/4czbwAGfx/57PpYKNOiR
z/28GceCAUqyRjDP9tPyEsplZYgbWiszH/lFHVV0IGDQhPPUnY3K9rehBD9B
TODsZPMzJipv7AcXx1assdE8bukYiGwE8TSyn2HoCwYtwvTY1UC08i3P0OUR
6CBxWlgJYxnN/htBz4HM/6l4NMBvE7KODDbly2+l3PoDSLKidBt4weAi7FvJ
XZJ5s43EEOs6VIddEdo8AOCyRLyipuU9oXyyrZZctrfv5mdkrdaGL2OEoAur
aaY8fOFob3QoaDezUCaD7sndKDyUFdUW6N4l6TGQQXlkURveneBzyDs9nSU7
11BGbrmHTrKxJdQkTulj66wpodPS8ZAtr8h4scNSIcoTZY16IPB2XpX5M2Nm
Znf1/Ciqk7i5RdAUpH0wwA6dIOOMhKHX8sBzPu1ge6BwLkjBpCtImEHYLbpk
KEqLpKFU4EdebyjJeYxvLg2OKAL4KURDvdUB0f5xjPaL59DDPiBkIldIABDI
xTOUE93g3ZyFnOP+zOSsLLE7RLE89ywfOl7zHsBrrzehNE3FLhCaW7ArAS2e
BpdC8dadiRrVhRgI9G/MUJMJvJsnOcqKCF/NsAaryBBNQjkjcuZxyn0S0kRF
gac6QjB22COx23co3aiIaLIe5qOAIUr1b8+O4aqqLEIUf+GvL97NHAJg31bR
sdszl8fCpJYp7TOKD+0jKGKcJwY0pp+hWpllekOvl21dvzG+DWcDoirVF6Dl
ScdUgbaTiAN/NMVzWy3o3rlvniT0czOEIfoL/4YkaYVisdPhlwBx4kYb9RXm
vBhmC5rkUcdfMxwXZV1nmz3vr5AW3GJcHqYFrXF5f36MIRpQ3DHkoEN5OD/J
rUIYGM13gcbqQiChn9okRkppYhXQPkcZU+GlQEiZiOKnaB38M/HERi0D9oWb
0x5MZaIVvdmexoRn0BTKNosgoK3rNG1Ezxy8NaVRNZnZys74goXQzdW/dWrO
Mff77sONeIX7Pst98b5BhOqof+hzM9JzZTsfcrbPve+m0ouqhpZnb3B4QaBF
mU1OMdOWatgCdSeWaigwQ9Pw9QSXv7HpOyo6L2Glldc4U16AB4Y5Uy0zR+cw
9LSQbcB74m39W518hH/fDn374rHkkbvF069doig0RVe1+ovMmCDrJQg8Ob7G
9ESPky3iQgFVPyY84b5HnPo6VfjsIipM+9T/kI3douUoi4eU5RxC2nyBiMlC
6O423Yn7MC2PpqBflmyi1aDxZUoH6IZTd83mYa7pEv/MOUT4Cig4nZ4Uw6ZW
l0DCiSSP44z7f2KAXryEX25qONV2oYNWnojK4lNFn9AT/Do5sfSYrCvps52t
6Q/rVL2e/AOMopwWuACRgSnjzSZ0ckZcFFA1mLiX2XkKBayK5QL2LL6/Mg4w
xnoGDP1xhtbtq9KrnkfocVmCDDR9xIJUUtPaZ6ADxBVcP1rYJQWOvPVAzmmi
8CHicocBX39cSDcQyC/3AVcIo/ADYi6kMj8eIOOIKeC7Qxim2I7ACeiD4PsD
onSsLpgrckb8jXcXzNsMmLBCiRs1xUm5w9Mbkv7kE/ddpUxHxS8Zx7dZhYWy
jb1aFBvLUIvKMW39XxmPwrFcQA1NtF7bjSBSDFjCstP6EN9O0CA/H+OQ99PY
ChH+PsRWpztqCKbBzt4vtMaoEgwR/6qSZChbtLrV9sBKBFO2yV4hpjPaLyF2
/SVdZZTwnLOzFvdxgF9wWk+5GlSk/BlKBt+V5yb6l2Q3L7S0uD3tpcAU6FiH
Q9xh0PkuzFtTNlBk0L1QkOtr8qY32TR6PYuC23QJDuhcr9XSBViZRNcOmrDW
EI2SukHrCsUeAdpVQlxoMWn3YQTt2D47pRJE4CBMIGdwHU/8AcbEJUgBIoU6
+lHLCMADjpDZGjdTcK2/Dasv0N2YbdtvQ+PaxvTXXdNryNEqYhZOnnk09afa
UsS701Lj/VQ6RrI6DKuRSUyCj05pL7L53Wos1xyicLilXDM0NcpHrftpiDoz
eWZ7xfKnf2Vv1oWZAkPVMlwRVpaFmPuWTldvKPKNvQndFmxkloBe9CL9yaeb
MxCobVuH+blvqke71PFsA85YMM4TOqkbOuYd+qJwdC8N6d2IPwZHazVg3BdS
i/D/ML14r2DvLquuimx0KJ3J2inw/G+GERMaSUtbRnQkvz3mcEGyVO6yMvf2
8LRyYQDWvNdQ/wzRkJQrj0jocjUzClNR239cejZXTvYNa5lToMYj+et5uhut
Sh8ClAhKXma3JNzSYHLap3K29dBuZbWKQcktAyrKylUNSZ50UID4UPV4FWJc
GFh19qYk1zznxBUblOCPUPaagqlynf9I1yAIzLsbR/A9B+K6Jcx7iVEr9ttX
Zl6lJ01MpNdqXr9iGfCAlo+AMby3d1DEETiEwEeHGTGDp7TQp84FGUYRz9kn
S7p7m+aXoTvBM6OeWn0D2bm5p0MZG1VcBXiBvEetxKUK4Neg+z3OjOOIHuK8
6VpBzROSayUVLWiQBeN8pEsiMI87IP8uURiAjwm6Yc8toSv0ecEqywGBcL3T
wnMln2/PVDubh0R+askd1KU5FDL9ddZt8mMpbkQRRKJV/3WmK10GPURZwnKP
9pNBWG2zVr6BohmLDPICNqKEkSjB/snvAtdnJxxdFJJVLZaCDX+/DaOL/tF/
ysRSy0jhNqu9xcoBOxE9tfWA/cz8aN6CypepoptnW2iDcN4TanWxo+yrTEQx
HwOOXyL3osaat5zf96W7G26zyztGvnz944g/bB0d/oOeh4LYLggXqNk6i2+x
rb8q6uGyD33Dj7J+PBEFNLptm+d38RpQvF1KbsrN5CsCEfNnppgqD52r7xo3
bleTHZ5XRP4me3OFKF/KnAIhDvIfR6cKQS5mpdJug2y4ZOr9Nf4K0pnJ3BK9
k0CgH2D507pVcNDFrc8AwH4suPzL95F/J2o/0gCL0GDRBdKbmdrL71x7Pxmk
0PGFENz/1gTZ9NQsnoGpD5qkuOYU8Ht7HJL+qvyFgjARJhqggWs0pvN5UBi+
q8IavYJgbeUymAfbqbbIs42wwVaVPx+YHnhy5X6LfJ+k/zf5kvArtIS9tY5t
5slIJUVxoxkgFaFnGVbbbIKXl4siRBerwzrngK8ft8SWbec6idmg2GyPT8uo
2gyV+7Ke2bQUVUqei8mkNbZfvPdWIbyeSv2Sw8vfw8mnUMYfxW2oFnA2ETT/
zr5hJXSdAkc7qZtdj6AhvNdEsyBsXH5swTvlsp3eBC/HWyaUv4ckeS9Wj7D0
Et7Bh3FhwaorxXt1RNuWV9T4GADyvvU0tbFtyPH5/BO5OvR5T3jfdRCCOwWi
x4sI2AeMRofkEEVTe34jukKz5l31k4umCFopM3jOgqn6LRPFmVKZT7XWkQ2W
CP42H9EKbsj2p4id1UIoGaNh01SLvs5Oc1Nx5wXyr6lEEEGEyX+Cw9aqorxU
momrvbV9Kg7R/nwsR/Ea59OFd5nw1S4uM8RwTQ0dvtQBXj3DYIDjXEbLOiRT
cKXi6C69g4AyDCat0P9orDQT29Zx0f3DhO52bTZe6IalHfNIHaJUNgDg1FZR
4brgatbOe+u4XPnOXDDBy9T4NNlaETHtNYhF+u906z1mPk7EHNE5ZeWhBrzf
G2ymcaII8d0jSMfXkUTdiXb1D0VVEj+TDTlWQBUpLKio1z8TuzsB3kduAVMb
vCbVPbdu8KUtxbiIVUZY7+Di4pLnPuWRHjd9eMyiNJmj7fo1/0UJJOSTUiJu
OfMVvMVjQlSXZpN2fRjezjng3usY+xhAlQKjROfUa2SekVARxqQaXMsiy6iz
rDbSA3gfW9S9tsS2aln9BVNi/IX4hkPctOL6sg9KTq/INPaBqc2K5otRTTpe
Ufrc68gw48p2zs5xDIiUuG345jVKv5Du9GlrfZEkZVqn1dGcP0bWrODbJDny
HARsVpcSAeLXU2TJVvTqcLs+li+iHWE/jGC2MI0Cloa4p2+q1E483vZDiJAk
RvI7Sj2UGOwTQkbXOQuwWaiFfxzDexWmEOSuDns62GxKpKl5bJlIEPkf3skH
mkmurs626HJdE+8CjDi1llVeejPkqPHf8dxBZEg+xppBuy5ad6I5wtYRrAFA
+7KnizfgdVcROsmICmuKAy0NrU6/TJUQBDATXHu4t1g4/5nY+OznXnMUE6Yc
OG4TZICso7Pt//sXPoetX/3vSuUaP+57WcDKdBJzeJlPQgm6wJ+JSJ0BJt+O
8TdsKcMn3xAQVjCH4hwQGynEhg8U2WXdG/nyTFAzkbxI3ItWw4XnpDKBz/f9
y4D81zVcwpWmlZSaLH5R5WJa8ESv/Afyf1n54oTJN0Yfs1+F8NOq/7FJiaV7
pzkcmu89gNo9GtUiLIOPf1yy4QH7SK7r8Ed6SEE0MIJBwCixy43pqI25v3kp
G14dSyn8SP4FyKuqnNVRuNu4GzWVtLS4JZ83t8YxMuukr/mHz0ssHxfa505e
lzYMmTEpPIBkikrmv0QVOX92f6k+LmIu+U1mhLxxLCtT+26A2C7jQIccjMPZ
QPdPFGlQnxmyPJA7c6iNrQjVVro/8dl9csDYbrSLJ0AJ/gv+hIWptI+TV1Ls
yq32uZZ4+WefcF9LA3C4OxD4k5gPXdbCkPsk5JrXBZWMcCIvcptl6xKifILg
/WHmGgFmjEOzXNMNwl/RxwTnun/q7yneEu5+8U6Fx1aAdRhYmw3xOvdUVAHR
lN3SzKlAkJb3atKDDjFAcaTYKViEWc2BB9WkWFNxYLCFoUuwJ4WID7i083xw
Wh4sMgebgWgpu0aKSGoeLovQkE6hwgbden0HKPiCOFE/W0JIuHdr3T8Qf9HU
mausjTHldIYURvawr/Ovz5KteB5AMnU3k2UO9703+k4JrY87oTN5zmVMNPXF
fJehpkh7pbCjmjoyAHUVBpg3CX25L0KhE80mWErdfk/xB/QS1bpWVXUhtsY9
aPcFJMI7spm13JNJtgRbn7rNcwu75GiPuKjwWkMLKTVNrDm0KP9t3LvsVbsJ
Sq/w4nu5AAUsaXBMuBMbKqdaz0Vzuh0Avfmj/CJfozBZeaW+/bhtvG3fhVPY
U72lGlJ6XCy72ipuYAKZrP9qwPlwKzwNHX+TFno/X3jO4WNEkQrw8bTv29ub
bmKVx5oBRngMxC0An0+7GizWVA1ZFoeCsuKeUI75zJ2icZy1+IKmX694qDbp
18vzCss/gwhQ78GTX9/pnYmZRDAAAr4/1errCODnOCj7YjftyQzOjOmRK5e2
MezULFOqFuXUHGV5GcPI7EwwiL/DoOBBt5lT/imVkoqm71FcqEK4nlmSjI3c
eo+nYjVBnkDiCkI3nUgdH92cvu72WGiSWAKQW64gTOpqQbHRfoVSZNCf1Mq0
QmuWckonyt5IaT6z5Ro3XsGQrfx4e2cqRm2ACcUZfa/sDcXC7WvCJhWXzyrI
iPJFTbVjAKpYMWn7ygTu9eZNMuzc8AGm9owy+BighqTnzJ6/qExnAkMI5M1/
tAOgwx0futqWwtSDJqhITs3FyfK8y4sy4rWZeoYb7xjEQgZ8QrHlBy9iWegd
4/pqyle7jawbi+9ucopJWTW4v+hxGzUXFLRs2jPgTjKM25ybCfK4U4CvlKlc
S4xCFzZLOHHIe8Fah/kZkZEu/jXijdNfmdmg9chH8fPhogEMVkri8UiZmZVr
fCZhCn16pFpdIcX/lgcaYPO5Ewf0yO4QhqSr/jKhJat9oGWH2orIDTS9v6Mk
G/U1ILo9muBOeSitbGChjh1O3MuRUINR8vGN17lUk1+6oMvzrexeDKXgttYY
wBKsQoUz8HHiBSwuL3/T/pzsvwYhf6yA1He/uiv2Qx3sj0qF9Md1er7pK+Pv
eszefMNdrhe9zGrLSzCzcpDMnBIFVlgw9QxqakqXkD57FCX7b7XJURJnQUbu
HnWh/csRpHo4QQn/kAAYDuTeC9as3xkBPwPWpey2cFIxufS5MdyAP2HUXiWN
QrIwsAR1nc+Qi3XxUiTkXkhxbfND27hAzjIxXM8LAnaGjzWG0kPcNODZzgNE
Gk4kaqrGCDVFwEZcar8E6SE/2hhJzw+aMiOEPBVX+itTlu3glKHgAEE1eoEg
H5y+aecJO2LLJwmh4uPt5S2BsHupYnZccBG2X7BVHsFCyU30lpLRgCQeEyuq
lwFi3QyBZ848c5Cd5jolG/VKYaZr5mWVJKgomEpBq0nJN4Vq5gcsW+9Znq3R
ADZ/exCov57VceqkwwxT2X5BPcc8ySigaKN4h3ibbmRdElYfkftvd2AQ76fz
rfAH2XfsZS0RzXIY3FHDxr9Z3GGpGfcI9g6yTdhtUiBAzU8ahmXjElosLAMg
JitO2aOQ2ZMm3XuIQkZzr9Dv+NbC9ewtXE+1K7jEWy5mRnEevqcto8HhEghj
ir8G/ZPU13chSeVg8acNuWa6+J9RSot8YZSpKF//NxMzL7Q81sOzlAPakXRG
dtnJ62xV/rC8bC/VAe+iBxtIUQTVRETg1OYXZrZOetSorXTKRvSDMl+/VVFC
3+6jK18eNHdSanJbWCN24HfhybB1f5Y6Uu9pgOW5Gz0Qj7kwv9dQJYnNiw6h
FuA0q5EuOf213j/Dfuwitf78V0OCZYnWnFi0al2KnJ1pxpmMKCnp0xirKZy5
Tf6lItyINCwkrOtVwxdZpfTvInxDmwecR4LYNqMHO6RuwNkdDzXjI/8cz+oY
nconvwVQzCsVXGdZmS+sVA6m/7P43MUY/m3byTdiXWH6tTo6d+9WENpPK9Xz
ParHuyP++KroIo/pORS0ZwaBZTDg1cb9wAGfh286g7uU8keMH03qrOpw5MeX
zSfPOhUbps3jqXFZgaobKjT5ao8ksp1UZHKW6owzi86BKOqSEkZl6ABH1009
h3WER1c8nvLWuIb0VjcpSjfmd/Mp/7InwyA24TOlbx8hRZ/frDuz3yi3gKrP
o0z4oes0Y2ox2Zswgh+r5ZjDo4xAhQ9dbPbre1iWFAt+zAV9oV/3/2gZWvH3
RUJwqtNpsMEAJRFF1F3ihbVDZTo7kPt3GLafMUrQRuPeOKDyLclO6TqGy6Zs
QI9dEg2XISKrZnEXzaDbNHEe+q6U2QfEgEPNRaDqqSwfznox56XHwHMI+vuR
805GJiqhaF7Lnbs6gsiGQfUh9PaS6PYYCKxkZqXfLChl/jRbxuDk2lDq+MTq
WKYcL11UG7ERLGf2LIhCmdVa3PVXChAqnmU6YkypCydGVIVJzTkHnEq+2/a1
jJeJDb/119wW9V6EGqUmL13qjCxttygZE0fWsZXLhkjcwNN3mCqJYEFr0XtB
zZky2NhWMsSK8PCMhFe1Xc4yUAx8eB3VZnMkaLayjjsVS4G4zIv4hUkp0zqr
1Q3yT8yO8HiGqWoRvlWS32/QAv6cWo1bHD6NJP0wEHJJkhzGh80rYOwQemus
BsmeZvc+52eU0OuROEfS3EaPP7a34oOGheM9ZTrV8hhWSRPS6lqbEADNv67l
QkgS9bohb+acn16LY1pDwST+BpxF+7690Pn+Nutv7JlybSqm9RnTAP/3nkdT
JTLZ8EeTlOlB7GkwreVu9hXh5HX14Swdutjn4eH2KHqHU9Tn1M8kGyHGeZlx
68eeRtV6xneG1hUPLeYUXI/SPJJ/a2NaCbTql8MUVVzDJcOJUTnRkTuV1CWS
J91BkQLYI1p2hkOlyrxb5doIfEFiULbMK6S1o3J/DjRoEhzc/MOi5UTy2dYF
0O6kTEZku7iBtSBZqPgRX1KNEBTcDAiABz1dlIwBrNJmn5r5bQEzVXGORxhZ
4JhoOqZCXYQRmRoqRbaSHLqcDow0zukAXywJAWztmfgOakRSs20nS7KKoC/u
vg5xehFuQ9ZtmLk6gu+E5e+j03eq0dLS/WuzRaWpuIfrne0hoUdV7BSunQBW
Hw+P+4yYGIxgFGtHJqixF6Ejngctoj2khnOVnQS+tt7Oml+c8nf1gu+NNbMT
d2zSj7G8+5dzPR8P3e4nScmU3Shj2RdOX4XPuXIr+cbLvIsFz+u5EvI9EgNx
B3ednDkhOTe6M/5iilCcxNfBnLwD2xy3SeNSkSgpg64nLJ4lJxzM5/IkNGq3
NOeT4GZYc8022FzTxs/uaAC2xQTSZYoAnb2bnAnIgt+8lTBSsoAqdx/2t7gL
yCXuVqRkqzEEKcIC7b+FpGgA2lE/Xsq09MuPIrCzwEeQoFwAXYGBYnC0ts+A
2dr9O9ptl1XcZMO0rlgsrFt9qt1+xtAISP+sf7T6AV3dJbbnLthkOehlP/5d
gHq8EaNe9r2vah3XCUm4TLpCfZne7dFW7W3ojcpN6NfMtaPObPAOA4nUSU4A
DP9NzNw7FObUDIcHsxcjKUtM4ugq7H97vrjSkvPOn79NMjSy6uDeLv9N5jBb
4Iy7l69JcbncXWTLsiLUsPZpEnnpSxFfMaE2HMSduWDlbR7jee5ScJJJbOnq
L3scREmzQXHtS+i497goxteWIbrSIya6IJu3etkbwBmhlAAa6Ef284oGaKI8
nawqDk7fRXQyUQehkjb++LpBMqonvNQBcfKhZhh4PjwHR7ZyeOAywsyeTygl
I6Tm18AEArGVUyllhr8FaiosLpREd9+vqXoUHyHuNEpdCUpB5HvEF+nlbD4+
X6WW+L1Jnfitsg/rGbsuKQTvSdP5OTU0VszWaZycdMf2ixG9MOroW45TxH/D
AyWPQ3/bzCjWhV6zGmGkB3VdaTLVspcMi2EKzHQ+fLiEvkAyaDoTn+Eo8HT2
GlZPHZlY81dSU6B0YcJxy6dfTvybtg0AnCLfjm4Iu6e5HAjC1SfBwXagt6N0
ssp9EJfgNMChmu6tpj8NoIPJlJwvFCmoxWwLA9EYvhv9z7Er6SxM7U+wwexz
5KOYmCCE2JAG5EMgvuihaSYCvpvJpCSrfF+vxU43wsvDuvOVXxY+4HDGKkiX
bByd3+MtMzwT47JVb+p0Li+Cju8/lQ/3EDlBvvdS8WjarZBaoyXa18HvnstJ
s/4OxVHsFChsvXubyqXIHaEHwAB6eFlylF6R3ZncVlCXt/nB62IdGry1Vxb0
hf7hlxzXRP+dUdIvaFIvty7VF/sTiMQqwvTd4VEh1LAwGdY9+et3yD7P6m7x
/1BwtpQKNOTVsSvFAcdSrJi/4ThL9r3r5tJ8F6WmNbtzlQo6aryvH5cLcEk8
GUBbV4E3pWaiATmHBMQYI9nFLPDRWdI0X7WWFC9oph4YtHFIBJ7ZIcoDQeFl
I/yfcvP3v1MUCHqZh0IOXHVdVLDFdwnQokb+69GqnyCHC1Vfk+fyjLSXOrm/
CCjQvW9ixEXmz+F09EvZ1EXCV/N1k5AK6xdeZ+6HKnB5wAird3SB46DBjo1p
0Siv7Ew1tgawAljarTE7eKpD2xUms35M4PGFIlzKBNkH5Ao26MBhfddTHgZU
W+cuT1oZf9Xi2FkXkfzYmNC6k3KI/A+ljqfJn6gH86Y+uX/XFsExZU9wqQPU
UtKAQPfkbKT2fcKoH+fzqkMtWk44bO1ILlIAqeyTYvudTGU801CQOBNCOjZF
9/UGSG3lM5zEMk4OJ+y+uh9E4KFVq8lQpfM5fXXm/RS7ThxLxmBiGgvbwnh1
ZtTfvXPCXukKWusj3cod612TubZQFRiAI4/RYRfo7INxi/ClfYBQRV1WCeMR
SDDY+4Zd8KLwPpjYWdFRXEJ06PFr48mAd+4C4S+0I5eZQJAIKXTPVdeoi1h3
iQVei/+k8zC5EDNimbnhKfC4Lyh3XwmLMm4aVkqQ1ftucRuZZC0nFjNpCffF
HYKg7RYG9scjQlW+hgK26egB5SiZODiZlTZnqVmB4o3stPHCZ2r2VFRZXmTM
mHCPHXe/o3nrpleFgU51eAkvgPHmG071Pe5zr3UucjgS059uWVS46C0nfALd
5caeZIts/edrEAUaHqvcKcPcWdHy8p+JOClISqkbvtOuPDeD7tkfNg2RlDAJ
mzPQlfhUC763d42RWhabDZ3ump7NVAFGBw5PgYrOmihjjk/MJm8j04vxGLlW
IwJNs734oLNBnMjv5iXPksu/6a/Gidwdj0zaEomd2xlE+XAlmhAa+ucfSFvy
ppoB/Ev+frAK1su2bkqY9J3FDvbpBkJQafHMg14dacQzV8Bj2wZiuF7lRgNY
y+CMzShUa1NUQr5EsBtLO4QTBeM25mYbR26Ql2hmSgRRDrFCF/3AlqU8pwrK
w3iOYClt5WrFgZMACjbeK6bu6HO9iZ+SqtoQIVGU2bplYVLp9o/LMslUtMsh
CuOk6mCEDG31Lo4K6U4EOvpOEDbuYEzbMdRmGOpdc3GCx1odE3KDWmC6/PZM
4OQQiUZHS9Zw6VbxCx/UNF83SrSIpa+q7Jf8TROsmeEpuXGO1uVu69Jo3+p4
NgXz8ldD7Cm3KbYpY47CgQ2NrIwEw5HgcG6dNluX7NS1r6gVQrFf5cLAxyOw
4xsxvhaJ07/mn3OZpRy8P+0whQmTQOukkQ0k2hVGLueH5yiYtNAyIpSEg4Mz
x+3U9aL84ap6EpR4NoV7YxD+MifOAxWs9lgKEfn3nBlzpdMJR2KPuwQ5JG0N
agfaqwOui1h0Jv42+hkcnMSU8QGlTi1f63Y6f+j1FtPE1lW3uAzDgv+OmeFg
unYOjTD/2wJHKB0NDjuoeA6CFRTSSPjTlfU11d05/npGaMZAlC4AcH69EMPw
zsUaaUOtfU5EcMv9kc6GBG4IOMGudQYytyWY1mjnYml/AtqwPoyZW30qgLL/
LXtxI7J31CK9gtKHdUznNcVmuU44Q7Xy3H65ORlA9HyC1oEmQy2AqZplf+cf
6LQ2I5D9JaUEIJodbqQLNTuR0i/3LPNezLpkvvXB2gdtkt9uRa8rqSoHZLmI
5+dZYFD2Mn02tk0LZZiqCbixdxOWxZnCuiGEwz82deCjHQridXZBvnq0GOe1
KjgJHEIzpkuWFndqJPsxutB4aPK+d9j24i48eQc9Vvwospst8WWaeo/UOuAU
N15z+Yxy+nlUslibIrdG6iB7Wu/AdT7fCITYsk/ribpNy0YWLtfb4oesJm74
7LlrS/E+Q3dIIAQe6sMJCq0+Y5YcSuYNuTfQvGHa7dRxzgBSwSWDXhP1ZWEB
y0/G7yb8t3j7Kmjt4awlGmWbG6t9mW7XR0fUZMWTVYaTavI2p9WuEiuVNBv4
a9fSc2fvuTCHofsXct7hZ7QpwTRJU0R/tThhdZaTUDzkR1egu2PpPOTu8Q7a
BA24Xs/a44H3WWvNHoZ2gqLguYshOSzfrunsHUW4ANZ2H3KP1Os4ePCP4KEB
3Na2g+pCyZ6CDWAhcxkDbz1dqu+unKMH4/gTT/RQBIY2Has1Rhng5ikWO+I8
SWzUBlJbniEkWiaeo9Ue0S576HFnZOCwhPnrXW2PNZ6f01krpaqxNKoeUbrs
TBKHLTRr5D098azUqrzQXErPDwXepXc6X9vsq8zxvEeP21zOwQvP5024MseX
XbnNhssVWotTT3aq9TMCc2FiN1lHSIHDrFWIPUN0wGcfvY9FIc8uI3wKowD3
bxBc8ZfNcbWPkCUTNDsAVCiSnABQBZCXH8cWMWV+JcHhU6sMgf9DT1LNJOGa
egDFCOJMwfwQPaaBcI+oBOs3nEvRS53sUgzoC5De7x9eAoy7wLiKL6Aqqmsu
Ujh4r36wIxR5ZnAn72NQzX4aPA0eiK25s79OfG5mrXnXIk5HuyuJCrs6/79B
NbWkAGhwyHPFjI6iYmoVo6Fxe4Fs/yAbwFZ/ac1BncCc+aMuszIHMzjnNfjf
vDuH3XzTkLoCWHGZoV7JAQ0EGOXMDZ2G8sGI3jbS+saxKTwV9LrxlP9CYpjn
ZTZkdSxvOM/7MBE0KVKBipbvbVQG3gs/2AK3c2jsJBRXIVFrcJSXBKyo5XF6
O4f3JYm8mxVE0NG+roWLd8fZ+cBvgxY51UROaMot7w0MV7pf/coXTP7ROqW7
md4x8sthf2w8/+wvWtqSZT6W1maKuFH7i7sWC869+l06nORz0cU9GVUDa27B
lEDZLUuLYghtQggXpgw4dyqGODpPLbEcG8LW6uG45TVo89up4mTdTgx9wi1p
4iYIVRKDYVZju/2IV9uBHkwt88SNFHR4JW/PkyG+PXinokTqGNY42mbSSC+2
pOEjW2uSiiX7jBgbo8P4cNCJYFtgzAxvLbsygoAeRPP3x+9OO28jU/b6jr2H
V1qcl8iE0r3WiQJJTHtsg2LWPPwZ9gYYBbakd+VkRr1v/t7Cr2RBZuaYGQJv
oVicxa2l6SGP2TID8J7+I7pwvE98NtQMELauC1lgqA2v9fhXj11On77VMnWV
V4yf+7U4NKypZPis1sTpGL+YKxpmAk6HMZTbhwMgJXmGDLm3dDahwHbaiVfv
9TYSe3NxPQrU5d2rcnIk8D/VYHCuUZwsHLBf8ZjYeNgPFhjJCZOg5t21AY+v
uP65M8mEGx6SD4BoSDlvjmHSErAc9rPmSoRxD35XZXrA4KprpSqPivHpUvQx
fV2v4KgoBF1si7bIIIovDxKPzxzPtr++TWCixTchg9x8cydQeX4/epnaIRTe
2xMCUqCwSaQ9ve2EfBW9ViCZTcs/+GNdXUToQPIhObbBnL64L3gtYGIwrFM8
kvS7JtyfbOSw51Z1CbgauGkdATOP9W/89MFk7bs9xoyuU8ZvSN+FAeZKJFSK
j7lcpzphRg2AL5YOEuMz06qFP5ezalqwXdHnkDs+HXl6+U/8MRa+JznAgFVO
eWw7V+2BTqT9UXCX1Iizixc42bhyoxDWYdlmVCkNErwiRpgDVujdQUyjRD1R
E4Dah5G4OpbrSABotX3KbcH4tN22uJKrp/R181kGGK0MFr9DdujSmZj+dr3f
wNEbTeRFmbSHs8rDuiDi0pmQQiwujXPPxtXhH66fDWHPt0sXWALJlzlL7fDT
J/0slt4s0alb1MjP6G76nbDK6KnuiG8Mn0Rqt5LVS9XHw5dgU1i6OlsYRCMG
z6s9qbCMPwD7v8dbs6YPnLx2B0+SaaLrsgCKIwdlEkVGlY1Nbv2mry3nn/Tq
tIRRnlhpw+3tjCRYkQpQjOx87g5mRQFc0FeOraEdWF3+ClKBD5v9V6bwuIKn
r2Cx1OBbKOdo0HGhd6D6zqQrZOHLstHOxipMmG2u/8GuXv20xByiOGyOfD7K
ZHrEujmtS4q+TR6I7JU+8IFzXs+/bhoh52SA1bCruytZ3twWOTQE1VZIz4aI
rys9YP2GVf+bb6fWYJzT6AURxBaL1m/7FoSatJbNhLtwKRY0XYhct6mHGKdc
MmdKeMlGa6iPqHzb4eqslYgMealk9JVyYuw4iarSqXO2IZGJJJvZ1TSFGXUk
lTcCxtr6asFX65fHghS8zDo6AWHL05Ihwaf1yIV17BVIQDvaCUUTfQIkBx2n
GED3SjQZ+xq7vHNIR2KCjqURnungmSgYKcRCV4g3Grl0h/qY5WOYIQxWc1YX
G5qVi8xeEMXsgXMBWek6yrbYGH4Z670MJApZVi5r1hP3CHPia9aUAxeyLzjY
1kKebdEflnAZ2OEp5su5RDqFyJjUmJ3eniH02N3Oghbmkb3VQ1lyeO/jdyH1
XkgqP7mO8UxHOeTOyOgJvJbGQAzfkbFRhQew6in+4HeD72QYackS3BTdfoL3
zPe8DW4uHOxeIJtz1Zm1iR5n2Dyw9D2zGFFqFCYymMGW6lP1yGhXAe5D9OOU
bXMUispFwkcZrMnpbjRh8mL9MgLUB5NHlAjtDnxdpQ5ukVxWbaNHj9fNFoG4
ltFUl2w0/Fc3iRdfghw+v7fJu9ycRIIVsv/71GqFKHugK9cyTe8XYHwipK+F
8D0FvnOFD0CziQK0Szg9eqnUfE+x3kV5n8hdU0m/LhJbU8czUgqyukVWMBd7
OcYupn4wL3eUjpKmehY7Xzz02Kp5m1w+3DM89ztM+5hY0nJMEMQDxR93Dsbf
5qmQHqbNh3js/P6Vcrgjsg54JhzJZZXJQuO536+8TQ/pN7NpWVIE+vnHHAPe
DkfX74+t7F3YLEGNbHIOjOwNCqEFF3xpwchn/vsvXGy90X00t9eV9lq5Qm8s
m+c2FG9eEafE59uz4ONu7K0mxNm7mXzT1CoxkW4dr03Kr3XmS3KGu6cNum+B
aktyiUG1U1MrU3egVD8qGtFO2TxLJCklm3gmhsP4bu2x2AkqR/djA5ab5HzL
eYg0S1kgOZ/GF8puiNZBtWWjvYu1xIaQs7Dp5bicJd5ejbyjBUsAp0gCkc2G
WP/as34xcA4hbWyMlWPJJ1w/nyBI2qyCop351x2/SLsS22n+rgsfAb2nslAM
FZaqjT+b1pin7LAKZWNx7W2oUMpJhlkcr9I6ZTU1D/1A69fq32jS2C3lIJgm
awadBpKgjnbMGitaDOP1sUTmqdrxyLDvOT5+48k2fDMYF9iMpcjsD4Vyj66x
r4ZjOo2LRBFp/sQ+H8z2Jo2EHKGlWUw+rReAaIPeu44oJCWpfZv6SRlq6hIo
puysUR+YiSQD2RVRTMHEelztKpbPl76AkLIVGOjG+LNvjZoGlEzkHRUNOt3b
O5t/uY+sdQhYU0OSj6pLrcAwt5RUqAag5+9CeMO1t8aPhos9B8RcHStza7ca
ZNQFSmufRGBgJk+nxHQl5QTgy2t8kuOsEGh47dQpEbMJLuojv/5hVi7hjyuz
3DLZbCyFXt6kdzdzubrb+CUGzTiSLsa6ltKFosoAvtwM6sqJt87vDC9Pt+hw
ofLhqYsThM3BaDFROT29cClAh6WW0UZi9rCvya5NZvMMZNJyPr+QzWq8e0LQ
wWGi71mS3FfuTkyMfHsg7pFsowK/oNj5Voe9l6jgusCnG0KS/nKZfXHXpHxX
y8NFBbizj+wk6mNmQ4ejAlJVCJC2ZHZmnLh4i7k5zs+Fy8X/fd6ymjdriCIJ
V7fo7llNPaZBEic62lUWFlgTC6vUtHFp4x9dOSUa83lX3mI5byJybK5IqPFi
gnCdqw0MD2pyGalt0B/jnagEnwA5TXnGPRr9iaYwUeeBS3DjZo9emywKSe+H
87eCufLNETnGltx3Thd3f8AhumsRXNmvvYyms7tAmVC8T3LUi/owSWwtk/B0
mSatZrE4e0EOFvPuJh0EWgZYsntpNqNWNwR0MPBEyXQUxndeANucdTJQSZO6
PITKuE2CyAjiXeN9zgGr21ezLmEtpwAhERqa1PCSmHrJM774cFf80HjYml60
EoxdCi15c3JAlKWH+XpjpsE1A9ZC0wWVxGKKLkT/4oO7wuuU2beXoeVC6Pk4
9xD1gNQTlFvxCTN7DkKp2GVcEfzCFsAAokENGD9wlZSUp+DNN2UFcT+IJAZK
/EF4QzncJxgEw9WZP2s/Im8oj7o1LayDa9Bl7BgxP8i1HZ57QHjwcXO8AynD
Jem+Tv1hgx+1ibRE5cokttgQixxe47cn5DDFaj89uDgQ0Uii5IrXurz+sQY5
LPdl96JsruIxfSBq8smIcu/kNdAKE4Mj9CWbQuN0z7CuVoSxyf8AM1LU6Z2d
zU5aWsAzyZJDWGrRD0VB0Z0IBDbfixFezuGPLoD94FwAf+IB79LySfSnyHOt
oywhGlfU52Bl5+Z1eesBLa5BGaJeSYNOvenb5tQj+r3j5vLuBqDsq3tzkB+R
KPgb/nVqCBhu8vCy6llqmqoMifTqDS6X99SW8cF7eQgwOlKMCNFB6oypfuVo
/u3bC2E5zfWi8HoHBMqKqLyonlPygfvV6zfcaihUQGe/nUxh65R97BG1RWdU
zRgu5/00wljUgQ9IP8NevSig3gcAcAYtYoTHQJFFs41OmiKjPz2qeoCleKkx
1ouEAtmuu2s+YnVZ7tXqoOAdi5W8oZZ+psS518DEN+e+pG3Ygvu54gUQjvSE
e4YVDtbBj4zY4uo+cDdUJ/eiwkXgelseYe/FqBTsnbQNGxBoQ4F4vey6armt
9beO77oK2iHhnBYcVDssQgiQmuN8fFKNm2RrE8fsgwShhu58P3MUKV/bfVXV
F4jowdUAGQCE9o6BEMhnr7Ly0CW0YgLLV1J0WF0sCSusmhdc+qfLNn5Sfsv9
QXG5H+WYSiEw1DDQ1Krxo8IhDgUhPmxzwo26BxxAuEyQH1+ktPJGJTw1Na7f
WFig6rsWv08t6O5lpERcm8j744NPC9c2TqIeAe0SzXQH4AeYwt7V0dFX5Fyx
U/jdchav3dnTxGW5/nGLQ2T6o0mIVaq5woFblYgmn/Xuzn5uWrHaZeX5wUDI
j8S05yDdvr9hiB+6Pp9fzfwGyCk4EsSZgIe59Lb5HGxVoydpC/TTRta4Vb6e
OaD6LA/wQ2iHRGPDkHRm5+2ssArkHB5KUIvrSaclvmqT4MdZiW7aZaOa30sU
SHWZsm1PBrMjPwG722BMx+HJszE6TA+LE7l3CN2wzk5LJQeOweXC/MtdNr54
RliezdAmfT1/tDsr71A+JOB9M9nXCMuD/0Vo8Z/NP7gpVxuOxcDNaHgIxF9K
8htgAM7JsAx41v2XGiuw6S4F8FgFRX0Ssc41hdA9zJUBLXWPbOThD/ASVmJN
4ddmDT6120sxwf0deeN94i3jRtfB0lwZ1L23ytDChdu4GbcibAx2eTYvLrlr
qfElf3cLycYkWCdCiBl9tUq8ifaUwKIlY8H32rnvLHq2IhwhOyhMIKEEDH0m
AZyAMCZ/iAXVmGBoBa/xaLFga5AFr43MiNhXsOr3ya6LDeRcBWnHkxRa5IcJ
JAl1HlIfKCZV1729V4C4gHSO02jiSPpQ7mlO7+/SjS+0JP/K8z7tfqgqFZJa
vBDkIiBE4ud+zfl0pfwVFv24POPpuUJWq5uhvUeDRdHBmUnUlv9GisF52Dq4
Y6cMcS1BqUKICFzf0UErzarSgzo49lW1KX9FQNi/mvsyzi3ozpYRlDch2EhE
wxQxkcz5W4Jh2vwXmKnBWKIw2Tx633lZZ/jqhrMv05FQQ6ytJ4NH8IpUteeg
qb5jxwYdnyfxseZPZ77HpGWZdsFknoEZeox/Fn63/N+Ifn31spRBpBBSFBMb
3LJKat7fvVA4XTYljjO9TzGZbab3FW+9i58XRFpHlZ0Q6wf371RGbrIsLSFf
MLLW5tOK9rh911QQ62KWD3/DUij65H2HIisxcEKlrN1KetwmRPWg02keRjBf
j55cvSnm9ikG+jvVczoQ+giDzKiRrSydJqSGBJccVdbDx+d8PNn4gllZpsID
u3x2Acdfl3hlYjtO8qA1Y5Ub0uELFOVHE7I9ndeyjgCL3azXDMX9OZBI7FUb
Tws8rIliDjuCIpFPUzWVMWM52n+1JLkOpNXofFmK/LOdwJPP57sRVgFUCINx
wbfTnvVC6jlW9UhCK9SUyQ2+sLmalS85Vr5OQ8vvrVyybbpBWVcHWKLK/c+t
WNERAaUayK0Acsm6h/HduzNTv78Kz8OCtF8/TJMGyu4l3tJKcZGahzoxs9a+
rtBA4OEGiHcEBu8JWyER4MkOFyvLEYAXIZrj7KNOwbTR6BqYWlrnhBWx7Lha
D12sFWvJU1ldGUm2CVkpxgOfQ3vk1Q4yd+QOjEdvMgyMSKpo0v0JUKMvyrJY
/UlDC5HuVZFtIbDWtzwFSaV+P83g3bNNMxlD2z0WlAW/qVlTTBVHQFdE4f/R
U8TpcC6/AQc2zQEPLEZdYsvLoP6jA4wopuiSHA5JKN2OSVzI6hHPC0N24OiM
ADzC0TA7azR0xdRvV/l7DLXgqPRaSDhAUuzmArdzrGk4fRCPddmuQjFlX523
/xPznCTykeWgPlqhSQFiVk406hk5dqtDB6cwGJkT3wVVrRQYkoofiNEsuafg
/jI/NByISq4pV5++l1axZ/mTnujNvDlnwZ1gh0+pUOUo/18bODMs47vxm/+r
g7gAzbbtSHAzVV7qKZocZFox+sIrRMt/JNbMTwSGkKV+UoYPxYviS7adbZ9E
uA210FvtsVtTnIg3kczI2CbDTtpqdKFrGu7Msh/CHs3d3rI7QeWwnjl4V3b6
rSxve4mJvs9iaiqsk+5GFNRp9mI45Z/YJgxG1b26hap5cDfffd8FoUhJLT9/
GhekgUylXeljBWzfn763+pYHokKwecg9iRnAXuLyoeOHX/k4YlgupSgH0+5s
D2CRzpkdGTY9M36hwxpnOKV7/LEHln+v4RuMAhDFWfvC3ooY1UK0Ikh/ouPd
ZUEOWuE1lfax+NA10k1m611zulGre2/vKDelHUArJzAuzYW/NvISN8fZjwZ/
LF7OdtamZnT+jNRqPftJlXqDA5rNiY5nGQp925tyLHIQT7erbR86zGPKYLWd
AAkPYSzt98xmAH99ZkIPSamo5W5NiiaHRbzPhnU05PVyTX/Z74vd7XETqzg8
84RBxsSkQWoWDm/RFoMS04uztoqM1mIk1OQmbC6e2xqz4RFdY+3oibrR2MPX
4HI84ev7cS/qtpZfNixS/DJ1VjBFsZN49XxssiO9d61aeXHM5zQ3sZDhTJB4
Mxl/H247avI6PXOmVBW6Km/Hy+z/Ii1cV50cF7NRvjM4wEnHP17kYfvRGBzU
qjaZxmSwEAEyDsHx6N+iKljnhAYTBCXWkvq+CabN4hdaWHHNRa4wSscJnXMt
8HM+8FT1/yJgkEBH/V0zA21Kh2/vNTPxKZkXjIK6lSbX0jXvbfh+Ds8e14ty
KSWwk8G9AZnjl7/+peQo4LKlfrqIouBLBf6zWhBV4oIBbe8z2pvlpCILDH+j
zOoemX4haDuTny1FOplsVz5v8J8hclsYqWbY1aLqPkl7Xu5yfjYLjjh1GkbK
glCBbW/WIoXp2dtv3HM3MeWYSOd6u7Z6o2s+/IYhODEIpmZxcNLTvL4SRVIM
PaL9z6yoYMELrDKPa3FZ5ZojzoSyCMrKrSuURtKsOdTsr++4gI1itNNuNUU4
Hl559uwUynK0PUOCF84Y0ca288kwNbbMwnFF8yi/d2sJ7NKh1nofFsGq2lhB
ZxH83Lkf5AiYvAmV/ZJGutVlyDsWmw+/jKGmwJJVTuXoxlShhxEAU9x/fRND
o9/fSwSyfvoimW5+zfjFHnw+IFUAG23tZn+qYAsLUrbWG4Grrp6hV7ff4L/V
5ZJgm5hLXW9DuvwdJCQ1h2JS0zYaRRABDUrV9xYQgi2XH2ouUrKOe2sZJ/Df
DGoGf8hWletL7SXfyLK7os3J6MOZ5knfbQiD3eVaouB0UEzBW4XzHHPr8ddo
7QCb/+y4DCqUFQyPYZDGLNAikLwlgH4JDtbOSfau7hURD/GkNX8ruS/YVKgD
F3PEql5VHJsPdk7RQo3LKrkxyh8jX9OOzEMlZv67dd+ud72jCdYQtWzTZ/BI
MD+QBucD6CZjVP0Sd/xeQ0ywepI+BWJVV0yf/yhmtOrrxBE4lLDSlmujcxsq
8TwyACjYKkufFyncgos5yprHDdARWp39AXmbMucDA8n5m7R5SZvXugdbpYhR
ksf6TaFC8pzjM/UnAowRi5/dAaEcOFPTWFrJDPEVrePgGjYK1YCnIt/8tpiP
vkCh5GUosmDjzTYKCkOdvbQW0v/hW0HsA6h5tvcg/NV+h9a97Umuj5TDBZ19
pMZYGMtOF8Yqzo68QRghfQQc/hkpKDChtTmF/bCjKFFlISXqxkeY0zQ1CJvP
47XgGMPPe8cYHtSNuBvJa0m8HeWz8dWtUuPKxERPRZJkFr9gpTO98yaQCzpo
Q0WjvBmxGrRoQHA1wzKUZB2rq3JgGXj00tTHY0y0hKAsENKmvrpFFwJRtn6v
ChMXB6DD7QqUW3gv6OzkPAbOEFjnzxxQ7lnUv/hGuJ4srV7bI/JREtil0J6i
g3XqsCI3VYNdXbVi2FLjj/06z59lGPgRxmbgi+bSLhHWycz9G0ZCWkLVke2M
iItTosFGzYZkOwicxIx1Aew8Y2SHXCWDrmOdO+pKYo/hrAPxmnmIW9klU5yG
6UJv+hOu9gNryPgkjiZNvw4A9kcJIccV/mRV+6Sgp93jlDcTXDrrQQjqdXOU
NlWga4zG04YO0AH3vA2sKCJVUgQ+FthtEJ33RmU0Qgq3gVYAA4fWg6dO+0Nc
IEMMlz69S644GDoTranSOnVnrvSmwyfDx4lvawIeUYCwNMF3ykQPwC/GolHe
jfei206Xmx3Lnh6LDAoHDRrrOgdya2i2M0kG3vD9fHkRzOTeYn7uef0EkbLp
kP4ypi8CI5Z2JyL+GLVFIRe7OlsmjXOYC9G32xr9H4QJAXkAqk1F06GPWj3S
0pJxtnURN5Cb4Fu8Q91hOQevJCuqRjE/Zxkezzv2pLIvCSfckw14yG0QIKse
tfH+wUht1O/v1M6ewF5xjPk1OuAoWCLYeEaBAGT9TDDaxIB8FxiY5iS3LUJ4
NkjVrkGinmEeI/AUtQ6PRTfAfo6LE052xoB65L+yDYZ0mTrumA/xMYU0MtnD
WV3PUt1K9H6lxS3fI2UimpvbKehPMZC3Y/e3jQlIUa8zaTr/Dhi86MBfiXLg
wICRgYSEVou2MeQVLElt8o/uO5MKespAdsIezeH218KCYeRPQSueSv+ix1KY
r7PFNz+zX7kMbZV/7Y6mMsMkJFgGNgTWreGJj7F9WcF6FvwLJeFIG6g/2N2/
HAJCz9SNzoQm4YLzYGQ0jV//gGXRwoTww/dzCmmOBWVz1yR5EWEhrR50xsw8
F9mdfX/VhR2a3n87pS4fjItV8n9+N5ggTXlnclb8i4mUaySbbum8BXeJ0i2z
FQYTwjiM2XXul3gZDQq75dFLE8Ljyz2w1TjzV6n2hDdCIKGa6+39zh9M5DXO
4ni+p3KELuGxAr8MX3xZZELWUBYVE8wHldW1Zr5/Woag7V25tCyDijq4tdnb
XePW9snjLVlRMdIQAY/F+/WA6y8dtj7AILVTHIu8lJstr2VzQqy/gyP1HH8N
iC4SS+2S8IRGgzOMXdRMLZnaMSAqcoBvM0PmWDs9/9/W5ESHjtmKSdmKeuX6
BQWoh22NRV+qzRA65lR3BHTnDYbOINuTTtIcRWYpLjar7YSwJgI0KnwPLuOx
nQ3hFeL5bbw7cVqA00S/VwZTathzscJs9cnNN8ctL6cGEuIqGhzUO///ntQW
AEHRPsNSesICqt5qzaaVud9L2kJ7LaEI9hUncgRPXt5+OwXPC3KyeLLHoTfi
9wICIyb7QyVr3/0FYnrCSE8X2YcqeOmS6Gcl1r7RFXvL/C+fXpRLvnGXJQbC
o9iv1dFgjo/fbHQ4vZ75pBzyLDgopHyyHUeHTC7nBKH1QCDmnWqnSbDvA017
Ukfa6nOvWLX2DjAfUivZ/q12eZBwNBApq9+IVcYhJhEHK1MRX8uQgWAPbXH0
Az/92SKh+Z0DPqpNJQcMlX/BFLBa3lRzYlC9qhPfwUHcTvWgOalByhFAcV2E
4AwHOiaKzgifJnidNVramYOtH8AzQFBqplYPM8/5eiqJ0rlYiexO9GUtGZR0
wjdoqBDvDYjhVpXUUo+q4SpEs1aAigA2vTI3QmusW/sf9a9W2j+KWesj+Tuy
SJpEMK7YTTcz+Slumo6vj5CgFDiPyB4SKNhQIQGHKms7LHk8kQ81p660pkST
yj/aN0rlPfp/L9ckjAmsxenJpCnkRqeXDtga40rHYZSyh6NifxNxayTN63RO
ezGeCi+p7oeU1Of6yrowXsXcY6fVxt9XQHr+EWiYnyzP6hGw5FEh9KR4Gqxi
fdeLShEMqgAK5ENuk1W3dnyN1im7lFmQqiCtQ96nMtVofaJ//E/V7y0O92sx
Vq0t1QB9VS5Zje9jYOS8Z2YuyxV//k5ebI74DMUbwCkypcuyH2RSOGt4c+xy
xNexGRgbRxuaIfNvt1v6FJ8eVEylUK8aof1td7jpZVewRAxgxTRSo/jgK0XB
mKRRsWfUmDllUwDsrI5i6AuQ4moufkCihA+SUFyBaQ31S88k0+5+PAnuzYV+
/L74TDR6EjrWsgLonjVsWj24wPZwmf3TSACXTBHQCBFx0tuOwvsDXpF+ci3G
6qv5IJ+mBBgs7wiSHih6/TaI7pD1bBLQzWKkX9XB/0g4Y+CTLHs/xVkaN3rC
xBlKwFoRW+wcvXDSvP72jMtkKemxyM7eRLBrovlEa8jDW/vpSs9e31OlnoOC
YVSbk6wy8ozFlkKq4/KQKPIVZlyAAmJDYx0KQkeseZi/o9Pwc5/LmLoL1thg
5D1u8VH7EFDmausoR7AOsrm8c92828sJ0c6YSiKQNmCorsyDpGHA9zBHWpG/
d30Yrw0j8f54/eHoqFYS3kco72QtF+A9WQVPWafBaQ+LUQr40noCboV9x+OW
r6Wmoq8n8S9mDYbXs1WVzpNoqzSXdnO7tswSdtVLuzfaJpe8u4RpvtaPovuc
ZY83McClucyxqoOWr+en9GF8WnI0dqRjBq6AZlDFdD1N/CEVfZE0OtjBpGMJ
fLtbJc2RRTNO8iLvNZli9804p4pDh5OpkuITw25CxUMn+yon1pdzUWwZsQ2U
u9ntLFkhSc5R4+5HSZ3Hpb3roIiJgoXg+pZpZIarZFQSb7apZq64ZDXHDah9
m4sMaxKQDkD3WCUpbfhEMb5fyhURPL14SBOWGjNCmbuQJYq3oiMql7OpIvKF
TzKuqyEkmA0+pgf4SjV6W6PmoB6ePJAa73VhlhBnDV1KM+8HGJI=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1Jw/R5OPLvKnnLIZ0oyjfwM82zBtCDnn7sDGjDbvZl7685rj7eClpmC4uPtH/ls0WmaJOnhrunstVN9PO/JayFg0yKKdhWp9qYc0j5m8NCkenLRktkYtG2fOzebSQKzdOQdkkD8Cxxa8e/wLTLaDvRdCeeIeAfHBVhvqPWsA64A3I4LowOg5jO+TR03886KzLRWBKJ4fXJawnj5nCema9bzqDaVfJ5jMxtKjDiGqxR5uLsS4XXARtxi3TbUyYBiaCrDrb1v6B6AZgG5aTCHWjhY19LNOhCQS/7tRkFF6XZFoSs84/a6JD2LDo/ILXT/vshNSLhGO8zoE8byCC4IBGCFPsMpBDftTm1RDx9w4iDR+zu8EjF9f3TCBrq3ijkdQcJkEAtHgaWmAnpiV4vWdDX7X+9c2xbnQhadK5qpFzx9efguPYJI4vFTfAuQU6jW+cH0WE5c3cZ+O4VWDObmJw4498c5RP06SYRa6IXTpK7heXW0d7w7nhZLIbt0a6OcjYbEnOmCqt8vhaNlHTfrKBfyC1Y32uo283wxUMPT6va7jH3YF4Ng06qWKPhaCihVlMZ/8VNNlHd3ON06eAXy7SxDRYwSbsS6L2ECXAKhh7TRcm9NyWuQAm8owSd7u1PXrPm5jqp/A9BAUp9DfHL/4Bg0hVH4/RZ3iAM1Nu2Wv3zukH1FVAOSMlTrtO/ou8M4C4KAfQhpnXTR3iIuOcpMQJi+73AHdnmXbUWYPWDy3k0pUBy+8uqyQ2BtMSDmW88GDNPi+3v9ntuMS2xnYj8nG08U"
`endif