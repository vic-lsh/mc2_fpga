// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GN8BAFlI63XxPER5zLG1iwlOa1eygZxRwqqqNusNo/v/JwwEEsHaiypLfCo0
44U8oti7C4rYqCEiE0bXdXLcfj9w6hR21vci61pwKWfWnm3yiGlj2KptECWm
RdP9ZBBa23UKZ9QJYx9I97Z9iCvnoVjosTUUJ0X+rvB0VDUV2i2eteOTR5WN
Z+Wt8g8ACwI0WYehyXBLbTk0KRT9Ep9ssoxfN+mib7gpvMHf7pJahvGrRnPc
HaW4hx+ak6CeEWHMT1m86pK0ref7Paj0CC9nr9HGYBJ81+oNx8ZxP2cHtJH2
1GZxGcphISu1zcklOIfvjVETo9YoXIbkibDtjHTEUA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mAjDwUASPTrFSdDAPM879BTota7kgWrW2JiGnVLOU66qswB6QdOYHTQpV7m/
fKCnHiqcd6no2KsBvckXC5CpgrB5kev533mtjUPMWJFMOtv2NGiDINqqXiKF
Y1TiNnHpJjxugu3CKkb7gVYd9pJ9xVij5JwyNhTZfXTLAxVXiyEoa7q3N9n9
4YeFpXZtP3MqaS6WLTL2HJ45Acot3mgWSVU/h8XX9LGv0+DaoJyabLylZCIT
Ms7iBWJ7HROWAczxwb2KZjKYaJBphN0haJT+ymbZFkEUBfmUy1e7CO3Vl0dG
Nbfg9rtBWiGxMSZ+QUB1fLcQU1uXw0irHbbsCokcDg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
irGf8IPtqgUy7CanOWRXVuIEIOMkR86rBUVvYxz3mGLoDzyhQA1w/UCdihOb
VxhnjopjtlfgGqNJgndx0+f6HoETkaVrPNSJl91zn0LFgss1vmJFIDInn0Sb
Lqy7/iG48tDRbXaZ3LWvDdh8k3PzXCQBNK1HyuD22VrbeR5uZ975NP5t4ppy
w8z0gJ+4FfOyOtHHOTIHOSiHRmnSTBAouissZAceUjuapyFlCT7b7lqSR5mZ
MAkYcU4/7sOaAGBadYBiN5n2Ichp7aDjlPHjJNatHgqkOb1HLGDUKAVBmH4g
36bDMnN7LbQkLMfcHNgH6s9gNcl0w29CGH1+mbAwxA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KV0WASSRi6WyIk5ouY/M0jatdGmKA4A3hqDjgoSmX2r6qRgBYqy606HoIIeC
V4v2jidWwINSv8RCb+KonJIBU/TUjtBuhlfRkeohR1mVSgBtKUKm+6w8sfuu
fm8wj/E9gFdtjjr5dgi6H9R8SeMQIgYZpITT9wZQjkGJ5tBH1lvXK9HTZhgM
cdTN6lbYrnqqqoON0+2A4ZgjpCjbVGIYzrkP+Gu+4fzPDnA6qE/gioQZ707z
f/thpoIh0jJ+4DTH5LjSMpTNR1j2QQa7KBb9SsVMCR5wpgRvTCG9RIEDD+a/
wPUTf+68OgkXr/rJFHUgwaITMWV+YyZ+GSBgMUsPrg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IBDVHKq28O8xXNb5Pcdyqbg8zc5KblbfGka8DMp1kN+2wLtMpC92Lg7S4uCz
qkgxRMhtP9fTQnD4wxCBf14d/HCwnrvoFsFC2AgtLESFqIPlzZm14tIZNU6y
uCb8UEa9nwb7oRYKtBhBTlT6NVt5JPI63oBMXmuLxeizR3D16Ig=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
G3Juxr1NEKnQkACWLEll9hDVsukGi4Asoeg/TcXQ6/QX5XHbJMgIafXDl1KR
TOmu1yrvSL4GMD3jJIDaAErdy8YBaDLV5wLGd5qomE+jzMixIqm23wbMFkBk
H02eO+dvwMsi2EEQgzwOGCIEORONYtdxUq5AW6g9J5IZ2Ude0Romdjh4Fb1A
Utp7M7RZidGhAlmntcRz8z7YyTH7g4mvG7v61cC2NP1F1poleyfC09JG1S23
kGY67pWiyRY9cyXUxdpliM8OUKV99ClhF3bwNuNSye6SQJjlUhyowVpYaohK
oVUcqCdcrtx/u6BWBT+NwcKYolDCrRif2pFwGZBAjo2PfFVEGl5Bx1knbG0u
43FcdDXkYl7riBpNvjF8FacvJXouTQAGhmdi/dOAi3K2+t4SPR6r7fmz/FYC
LZXkiBGlPv78pTemSOMXPJD/tCt+PVdnruXQNT6MSf6KJspmK5IsRSbOmQY2
JoB1z4RIpNarFp4fGiPSJuwSN2ce2aFE


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
l1dwXys69/YzhFLS5WxLJKzPD0IAGYPyq9pb/ppcCd6GJa8vvaNv8TtyMMP3
nJ6wtiWxDej142f4HfVkC63+bVU1Z3rJ/hsd/V8ZcyBP8Q8THYfXmXleG1bM
aalvBmP7krvtV2bfzBlKwjdddl9IPmAxkbFgUDimb3pFGU9yCps=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hkOhCjujAJ/UbDPPwPkqZfoFMZYcng3zjg7qA8vvs1cxroX8nzbgXS3Zda06
lFiWy17t5dtN/BIuH9EgvVszGEvLgv7apqPbe/s2G5DoLdoWSm5iQG1YwcNR
pKshov9v/fjqx0SXrLLvb7VThdmnGsBEjGCAdu5SvXLkt8slH1E=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1312)
`pragma protect data_block
eH5W0096DeuWBEq12a6eLQITvEMMx9hhpFZV+qlQulBM64K4WARv1Dv80cV8
c2qhgsnSRcr0DjDzWyHLvp/582PprHJfKXmRE0k2UKWq8XEsHi7dPWoLSkrB
MyuJsapoKSoIqPiP8F7f1weagUIp/Bng4XWD5lXbabPbQ0zdAPhIAlWlRCFF
jBMmCuPwKijXum3pOeWJsvo2+mDB2JSjU9Ar5DrtQP0AgqZ7PqOEiRsWUZ/c
JZTijeunrzeCTucI+vJMr3TKYn8pB6AjL0jGCPP9uSkIOARw17Iqhh6K/Bb7
VZ1XXi8d9TW/syQuL+epMMDqmAIf/vMTtV59kQZQoUTIPYT5eKHjjZcujSZH
WGGTLCW4jqizXrMDDTRDn7WXAazcPciEzSlOzW7TZlcLl8nlaUPR744rOSjk
2BBeod/JnEGYBZ3FlEZroJisW665Et23tz17CNAmK8x7yMruKC48s6nc7KD9
d7T4A1hZRxYv1qyrJr3g6TcRSKfGf4KGR+vC89eRCOuLz/K4eFrq3aKKnDeH
zGc1s++WEhAnpY9dfdh9IoQt+7W6TMkjYSValOWwx2b+k98nC29WoTJ7vkCm
/6Pdbbxv2fphl/EkrxH88dexf4/PZErF4jGUlDT46fsQuOpfZ1GFhG+hD0hi
KxRIlw1coz4WDzJRMZ0qgo/KIe1X4u389CYo6QDd+4m2bkzgnCDjF9s0VEqC
Cdm0LeukCLL4jqWcnRJwHTwpByR/2NeGeQYQUk7P+QqWvPTpOSNg+zsJBoMd
Uz3eivM+hGLGJsm/FUh7VMbomEVBKoP3UTInJhBL8M9UB2NIIYHW+sOONGAd
fleThmXzD73VpIQb9lVKRKvvPrTEuYjZ/T1nEg/oCbEuFpHPPWAu9qksu2vS
rZuFi2Ps2hb/ne/srHg2Y82EgvlcTFtTGE7LQzvdfGMfB8XfXxny5qMAQwaE
sVYS0B6pMaYsjbw9XI54Ahdx/jI7iSz5I/9e/i0kSxDd2a2vJlz+khwiEYX+
tZCt3OxvCvvW9vY0ZJylTlXC17NbQQwgiCHOhAinmt+iFYf8ayQlLG4yOZJj
dQJ/JNnufIHeVumxky379D8r3ZVWYaiH58hW+NinHNS7cNlW1d4A7ylGprvs
lUPxqvQFiOCZ7KxELN4rcsWql4Uh7ALmlQxjY6X8I3PQZWXfMzLUb6PWM6nf
3KfLm9zAhhDXp3LtwrJonE2vQKsz8er+mVb/Od0kNu7jbN9HBdMSKkWIW5Id
PP1tOsYBqfluqfDmBlVnzfOMA1/Vslg+i1pljaGLZGIq09OkFyip2AD+ZCfb
XHmtDpTKOIFr9lT+Sv4mKjmlOUbMlt7EPe07fMN+qVNjoGS1QCqY9b0Svhh5
iw7nO1tooFcjR6wWxuvXIdsdA9YPYN+U0o6GiEW61tb8UrpcIyFJAQ/wPsxg
DfDla2RXYgroyGB49AWWwR7/Vp4VEiXEgZyiBmAK8D+TMHKm0Fmz+PafqqPO
z/YGb7RAqErWKHOw8dQBcxxrnYE6Mu5O1MvtTixLa5KA6yt8NvbRTHnwp8li
nRCGxPijwH2SdYaS4mwyo5RPLWzRoh42ONdPl9LDEkrn2rS6gCCtxRW6MHQL
Uupb5hfkV9tTn7C5MfRPUXpTmr308Gl4SkX4/WPzJkQkIJJu79t7lQW5HXWP
6p5JUJSPfVSkASubFYbWiytJvpFjb2fz/e9+xTrJOX5fNTvgPKzLei4YAvM2
QfAl0xdtQg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQoxDGZsoMBDKvzNaNzuo4RBXSPB+dRpyk3mbG85wbUXBoDYh51/okJMsPVINWkxin4GUToG8C9Bx33RUIJJLPoHKkkU2Vgy8lanEFEbkQRhEjh7Z1eBcHDPw8YE8QwDTYFu9tsnuMQfXg+y06yloeVoBnFERxzJ/hcu6xzFGElnptSylNGqrQe+CwRKu9MnpV1LR8Q/T5NRR95XGnjlaTcgwrwkT6JVKPk/SWJebWEObkdztJBzpuoP7+7de6EjB6vslSJAmggPRNP1ZMV5wV5+vUCpvAjbLCQt14T/s5/Dsq5ezVdJ0/HKU0jNMXi9eN2KBzHAAEYzpSKnd7gajIKuyhXPdixk6KVf7sv58C3fSVKHSj1d9nSquB4GyQ7783obHZhe4LSfqYu2UPs1BhZQHChNC+Zj+fBVSIqWZuon8GUQtmLTSCHKVqIdr+c4RxmzEr1PB5gRBzVkDHNFEPdwqHyEj33+NCqilMUwEyrxZJJoRKgvHqzksE+VpRRvYUj2VkZLY9ID9MDZLyIjBhbwkZ5klJ2nh68p5fPh9B2YYR1BNZXk9rIsZchNanREy2SYEitVmS7xIQLOxVh7L1raCwkeD3ZpQZmc2ytU06ofzBe6shInVvjBUI4aydu4OlJx9FFM1h0gWb9Fq0kh/7z+cpbmNkvkV+f5bcvwCTVRPtBsUlulFlkOKTtvBbwcmed0KFyRlgcjEiUKkSWD+u0WSR68B5/m6jBVEJUYiglC5+5uqVn6nuWqnF3sz7d7QNIUtiJ761jilN33AtGOLfZEa"
`endif