// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
er0iuuuh/x+X8Ai0t3Nki7f2rENIJwBXx1WjXHQBYob/vNkaApsn5CirvhV2
J1mKQpxBRoWfzmYh6rMuPMer7DjAWtOE/4TZrGXvXfsNWnPluTw5YEzrwRh6
/yZ6kNZtpIph3n2FtIpnUsQC8QuFraQCIEqrhVSK+gAPFhJHlIK40rJPqE/E
sbetTzUyOSOpQ7+Vn4EB9Wp2007r+7ARdCdQtgMMRc6TrhQyotL+9fMzkPvi
4kGae43eD7jm1N/10J+jTFzoMt/4Lw5Xq7u8B9nUCvzT4M/sxv25008xHT8O
BuPJ2AlmViTrOYP8mWIYA71odN5tY1MFq2396weRQg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
naTJKNTgmDNZi4FSdXmebUPVMWYGO8wmDijH0vmUALugHfl8+quGTt4hFJ7J
MKAEDs4nJTreexLLQe0gkXgfsMrKfOVDQYFoUjpbuT8umZhgDliFsJiod10w
QiyGxTSMSFDrM/SLRamBBHlXmdnH/gzYaTbKjDPEGfQ7J+U3pf8NhMLrOyV/
yLEVMwg37j3yJzoTnDBaR53k4T411S+mmCGlclp58gybmYddsRY8LETBfkzF
BoJaP0G6dEXpkgj8rOIGYelp2zzjhdzsri7ijH9n6iPIfHerVq4OXeZCUFHD
p+UHSgjxO7uyX5TJpUHUlAteyudSYQHtV+DlxgGs0g==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AdaT3uEnaBXXFo3LKm5PWfomu36F43OzisilusNFwTsu3i19ACoY0YCsHqaK
wmM26zO+b6lCd61WgOScqtVNOHCljMgvFlcHCBtZtNKHWw5870eK/NLA1adt
4pMcarHjoJFkuhdiuNoRT0Ja/5uEoYm+9B5Nz0IeKV9DZ2htDXCwxYtRk3ZN
OxBP2O/BIfn7dPHW21hmJneMQlGR7A4as/jIkSrfB3u5pge6vDXbUCIXh/YU
9zjGIZSOKlOBtUdFBiDab6yCZinhVpTsoQl8CpDjinSvUwwlnUUro6zKxacz
dkabjTDhav5axuJPatLmAHfonrrnEc4s/lxjCnzf7Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HpB6niesySMHbe56YfhZVcq/eO5Lifcda2QgpufTbmKAYSm1tDSBSYWMFmwI
WYOQk9mP1U6QF4MuIHrARYGhGM2ENy9/fuptCa5arPqcxSzrWZvJdr3rKxdY
DEMBoIegQLdoMIgwIMJMMbKNt2l8agL0GeBcIaKwmTesPuWrybXJCDkQTOpI
wqbBNqP/0RHT/0jqBx+iY86Ow2LDlcEjgT6H4oXzT3WwSgRAKrWJdBrlkc19
MruZgg4JsB8HRVfJ151+wB6XOoGy/clYEZkuKemi7+ejHbCLR5XFnkSZRHe1
Icui77g1lNypZ/mtLoxx7tO0qpLoLFPNsVGZWcESwQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ii9juqsGYEDoWnUKSre/oS/y/jTg3KI1bpKmadSnloSESEjKOY0vRVOMQEJY
LHzAph89X/jcZS4qW09W4sMljEy/m4zil61g1ymlOsnMhcEqiUBhSNGI18hO
RK6Wc8NtBSUBdYf8fOIh8CTF+QovkFcOQDmdY0SQzUrQjXDiFMg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ZgQktd5YD26h0zj378MEPOFOoiLgJefVCerVW6ahewWe9qMLnF7p/jAZ5S/n
7LAFIFoeN18MOahgUaYmp1gwn/2ACNocjB4ZTQ/CfSoqC5+BtjXdSmORK4dc
oE27DJF5JokUvWagAC2BeI4542c8Jwtv+UH/jWpToMp8ObAq3dQBI3wstDky
TulvYTJBZYUiqS5pRqkH75Fpdi/DvB2pxvCuFnDB+lGGIJuzr5r8+NyuiS/y
qixb+X2weEzqfUBxrbtzo+VfDBTQlkV84IavfComY1rLQn0PHMKUFwsosjQk
0fLDKFtdSLNqLhIgLlZuLC7Y2i0OTxdYZR52FPwXJaZNREf7vtD6H8+81eIh
MGjXB9Lv9lvP6t0D2SAuk4ywShrTEYS6ZTRYhhMVG3a5DXu6BDPIxuP3XDPA
jRl/02+Qj5xTncIS8i0DmuecV7LyVI4dV+1iGh1ql3pUgMQpTxe/Ze06Ubt6
ryPYfrTbkpdZ1AeReCiNvM/jd/0XmpqL


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ucIxYM9URM/5sMlRGXYHYG4/VOttEkdIF8Wzt9QWFG+03IDUtygltHutnzaz
vuYiamdl4bbCKbSQ9YKhrOIKwE38dlJhqKEnA4HUZxSHzQ3Q2IxNYOkDUZLR
LVqWaIUlhxVSMgM9X7n0Up3n7NHhAjfiYPJaG+F1ml4sNp0hHXQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cDH9JXdIE8TmFhbgJe7l7AuhosUmCMA0SFO7yiB8GqnjvlIP32xlNugI0w/8
E1A+BKggFTqgY38o4lAuygun9WvAfWU4Ww1GjCoPp5bmfZ1S7Z9pH1K2q8cx
SOU87ixrQWoVXa3jDpocKyF0/vxPCLhwHAq2FHnLg3o0yl4WmZE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1296)
`pragma protect data_block
f+xy7YBIkL+VK8YgPBt3QgIAbtC8/YdUHwweixOOLmu5n092mUhk6WgFy2Kp
nTSFeoqnPYEGBh4vBJ46dMuRrv9aIqq5gqUXCGr7KDFJhwQPM/uSYhQyp5a9
OpJHvve19WZ7S9XZZTcp7fQWeRAW+Bzcu34njr+pXz+T/wcaSZ6uNsJGmFYi
PcfoTj1WvKOQ44IExUEbcSe1iHPHrbnKZ7cOouWagnFP1T8FjEOhIiT5K15m
bH4mvkGCPi8kbTO5zZ+T1Gzie8CQjDI+Pr1NG2mnCJpgPnxaJTZxkHlHiLBo
NFWl9bYwFm2o+AHFld3kbOR9ZbE4dQeERirXWHkodGjYRCtNqs1Uw4swn93F
5YPMQ4vyIeE3/PUujbqDLl5IgNVvClqz75Y5qsFDf6rxp+K//OkFju2mLQhW
IvTlggOrKrkd94Ypjw42+30RdQWDA3AqROp1HLTBb2IIt7wx4RXXXPP7X+kS
4w6KPcaxrNJZ9MgmjqbCNZssatsJuZF5iWirqMKqocMks0UcVSaToFGHgcAu
ku7LaWXV5iwHrBk7nNMcxv/WGk/GENjOdKd2W13e6k5fRr811wvCTfU0DJml
aNwZqZkcvIz8bnjPe8Va54h/zuO8HjrPFGWj/AcnGsLkiGCWkhg6RB9CZxqW
PrPzLn9MohgqGeR6Sl28qFFDIo2dQwcsc94SX4EJYQBNtoj+Eeyo1astovKU
HSJ0tzTSjxERw/fnjeESmI544oPAZXYHqWRm3OmeC5MOQYGzs1F0McJ4Ibtn
OWXTX/LkhlBkgXCtrw4PaMn/7JIft76z2rBTHBzw1Jvezzfdb9V2kvgbYQZJ
YuCSc4AjOUE0JisLDwyqbSscXh2/EY5VYQMYopCgkm/tteF5cNxh9P9OxjqR
l8MwiT/jod2K6Jkz0ym1zK3NjWJ2GqWTIETIPfFerKs2LWgJtjxoE4rF3CAU
N+ckjlEznP3HxWzbLQaWtLc1xD8Ao1GBvNBohiFtt0cLFQy30k6tpgb9avqa
p1IXN0XAccuKbXGZAw93ucwrpyzjjvfjFxPBGtIvqjqgp/CbdSDBES07UDL3
/ui41ad0oZJGeaGAm8KLFk3C97Z9qF0F1t2PqmWbHL/mKA0krLsHtTReBAns
E/7434iesJRTRSVns1rm4JYIHICznbBQvdG6o4rwOIawKslFMv3lsGWTvO7F
N832vp/iqhCGnGbl1UoaV3CPgNCTdiX1qZecMYSBYAPkLSpJE7FKOYNA1k10
SMUgNcePIhYCcenAywZoUmTNGYJMyKiEp1RrChLA+1l3ZXzireXAJ5nP714e
R2RX4Fps5w8RYfLcUOZ9YLvi1cs773Rge9fK+Vrg6+ktbM3A99+E8FASDc9C
Dh1BGE+TOYxjTdIjGGIT2vye8hg8o+uWUNbjpRVVpUPMAFlE52J68G3u/mWf
stUwKjg3A7anMpaGijtfpv4QsvOMZrUB5+AwTZRpRDoDMGzRZYfF94T1nHJG
NSfXQNB3bDQ2l5yp1VxgSmz8cfnOXdmcaSWkO4rfkgqhHHrS728Tdn4aqCgx
Xu4XL60ZVAWGgwBEl4sMWv9soBW+QOrIxJ9gq1ttPRrm5FFdhKpO0Gr7KHzj
FRHuRp2NGbifpgf6e5nivmQLItEQnT13uHxhWEjGdBq4tXf3/WA0RqMiH5fZ
uTileB9OtZaxJVaTgf7LuyeCsJutv0f18Bbe84OGFBtYDaWi

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqdxH1y7PfRNf/68IsUPbqm7uXfWVCRPcRUeOx0xLttH8Yuc3lejKZga/bIJzxtxghwVFpWliuzKbKz8QVhLfO5AcuUQi2k8xQASSBzIl1SfyPmjnr0c3FHuivQLokbKF8Fa34tkh47uze/3Vw/D7vXlxhs0Lw6hU4HXT+Czak7CfgOTs0hVy9pdB5pGq/fMIcymKYq/nx0qrc6YTUKGy0sYiQWPOBkYzCdzgHRV9Fk+tggp/idFCwnOwmRCikEO3j6VigQihAXjfOUr9czWPltayPznpFfqRYyVWu+ydLIzXjqjqZqFVGSoS7kl0EemmgEFDI6K3rEDcy503pdIfqP89f9K9OvCTpAR7zABiZ8k3d6Xs34EyB//lN7SzLlCDfIGPmaMBO+3PPCxsGXM6CURYInftmgtEavAmgIVLfTcfExKWW+pPX+1vdHfgdpvcgXFWbzyjfKQq89B//nuhiRlekEs1H3WcPuba7byv5Tzgb12NU5XtcG+0o784s+/wcJ9qGXd1XWVskq8kAUXTpxtkgQBuOSgutzYXhPFpYxwMtDo0MP9RA2833gudGf0P0LUS2muOJwOvB3IBrBevEVQRL8p5PuAJIssaGuCQOBQR2lhqFHKUXzmVprNIfIgdVScwvKnYvvbssrXpcWo5lXmW4lOWlIchqJskyB+FaFQbte0Fu9/1EX2TfkQA0QBk8lpNb1YIiayjcJLlwIch/BbxnAQtD37/N0uwhWPKl0hW5fgUKC5FlrRMQRwtZCxHkySwMDqpDAjqQwuJdvphMKq"
`endif