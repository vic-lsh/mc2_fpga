// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Tm59kEBHHBxqsvsW04/wygo0SmLt2vubSUR9bsICSLX7DUx1f5675nvacsdE
4y4B59/BOuRZhKZrT6/WQm/IBL5vK6DIUTen36thASkn13+2crRwVu5+5bZs
IjjltxLhOA3lO7VJUlQK8/QzkA0R2O5IhLNt65lb3i9ge4HW3WNXLMqxmid3
ZZwVf9q0tI1QqD856Iqd9DJ3WLTtuDpBdqKK82P9fWBu7OSx0EMYhAZ1pX4x
THBmWLLbByeTz2+q+bccnSiC4kcYezX/FOw+nopoQ7L0FJYIefPuISfrpL9Q
UWgiDplE/G5FLe8OYfIxSDdJqvSiWPRyvBq3eM/cTg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SVTb5oYd1Q/RPnsFewYaC+QXmNgwAdEP3LHvcMS+soYs3JFkvT5D4+x3EHNH
KOa1qyBA15GlmP5taYWK7nBqg+kJZ1T2sRoyw+OiJS1vJ0QCnRKnSvZDwTFV
1NaoAc0+odau/cNQzSG/PLfkrl8JLb5EBWNVcOR4gEZQflKqiqwdhk8OniOs
nTguna1/E74ASuIoVAscCX1jvHi8FUezp4JT+A3YBehxoxeM1mKKcsPdGlTy
UlMr6drAfFLom2XstLMHlJJMWkt3+bi1dcmqPrPHPUbCAJaQ65lM7kzM+ba2
R7i0fCkUhUJ/W01eN1R/ZSanxMHV7vRunZwm7LS72g==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GtlIQdA9is2E2YVQVK/Ru8wk54t/ykhyPpc90Y5esLWLsexmUSLQJ1ygX897
mTR8zatabWxQpVQKLE7QUwmVRobABzveBf65xR0DLG1DM3ZMw7VcPvZUmZSM
yXjJ8ko1mXP+kPqz61BYeRZryRvHwnQLEzA/eyx5nKdRdhUbiOLzobV3aNig
6Y1AMGQ/jmMA1z2OMjIc+QdpJ3qBLzvAVZgfDTxsNvjAxH18XJJOKuQVw4L7
8c7Tozd2XbDcF/IqwdHkkAgjM46AOpntKsWJ/U2bIMcVRtbtMFUEPTdj/0aX
nSCm1KdsQlLzZahy6u9hV4WD2dIkWDErpIAUZbPzQw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Dn+CAnQS/SGD2IV5PCUx4m+r09IeM2+PGHenDOgrK5bXS6izYlobw1d/m5bP
V9Mjxt6T23Wzwvf1DtnodtWFFBQkHgX25QVkrdr8BmrV7xPOzw3MlIxHtutB
ee+fv/Mw3hubr0WqbyNlToPD7Z1Zbg4v4JZwtwaL++5YGwsbSIZDJecYeZmA
yIs5Avsy5fTWDH6Iz/cU2hcyDqcr1eb7aAYoXxuabIFMHagpfBcwOU+uDXim
sEdNuRbyF2fnpnB399vkM846XLfJlZ3njQGY5KeDYAGyIY83qF3fDTiuRVAV
padr2Eed4KPegThrcJBHwB0JKgL/kCT1undiwvPXCQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JRoVuyKj3q7usVw/NGdnK3W41CmEYThv0PWdRapdUJPLKT8eS3f+zgt5jm+U
ci4bqp7NiMfeeAySVVRZFG9ROwifhrzJuU6OYfCEYt8kp8A3x1x17kgt3s1G
q6Dm9rBn7lrVr9Pyo7Kx00lc5htN7U9LCXM4wji3toruQPyHoTc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
eF71d80GfDI/UIkMJgx2PVF1VjpYgRlo+0upZ0pe/sytUGR4qYxDzo0BbVsm
PANToFdDrjV2euBSrkIdgdSaNnusC6KIGw2Prb1U9E1MLUvdLiC0Ou1TqL9l
81uhAnGyDpVDn7GV6EQJD9fQ4h9iM0HFe/izqh/zDoQHWu7cM7ey0SbMiEcE
iOmP2qlQuSFnb3B8sSg69gB0TzrtdDLxhSoRZOnn5ASts2sKWs1tOxey7Nse
WZuymwGfIdDP1uYBctDTlQ/p3jh73xhWqBh7nKSABhspLPAxzfyEo0xPLqLC
0OpILAT1U1IitfBki4QTCFFFV+cG7FZXI7niQBe4rH7yWmvPCBUl163Pyf6j
FYnQW6tu6oYA666Zk0dYkTlyHRJGG3QLlOkSe51BUmHqtQpx1w0fbkAPnb0y
bnEUtYCjoNuB5MYKxvDDmHx03KXClo4NMlPP7D8j2FXdf0Y+3SnNc+r4fYD1
v4JVrRh6eOpMWL4bs+x82EpqCyE+VHoi


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jVj2XIO8Co4QbBZQPuhfz7bbX1754SoTz5SUmlQ8pvZPHuSATO/mE8UYKmeq
nK3Z1WmRYs4tRThYrsAxPKxediB/UbZQoXaBpBy+vXNlHD2HxUvDCXGD1v2a
jUSGT7mEPsPVJG1hamgfCoP/QEQXRCNLLBHEO9EeMawzRGnuzEg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Wztes0bX5w2gayzroE8fRWUncq8S1G2wBGoiOf5x5dFZrcOYUJJyTcTZaynh
ZGG3LoVjJKKZI2Wlmey25jaKx2X7pwdT/k5nmR3wunMMx5wdAu+q3ywYJBXe
rS7jv/GoQETFHNtegqlc5gW0n/QVq4wylO/aU2VHtuh7T8QXNtg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4256)
`pragma protect data_block
xGKYgPcePGSfkllOJGtlYy9xOwfc2r8Q8lpuWg4mtOZGJz2vbCqoFR3gvXxy
IGMOlfF60SPUJ3J5pGOESwohP0OYq543DtLlkSPhEQwSW3uQiWqHYSrdO+Jl
CuB7JEjHUe8HrllAUGtPem+jCvqjzX0198djR5bef+Ag3vdSXhni/MYX/j8n
9Y4zmf909+T1lBfnoADqMt9XLeT+j00eLOY8z8SErOcHmOK/9m/Is5HRtB5R
WKpXoD+oJhli9/Ct33EgIFRRcdrflucY/2o2G2yfZQr0uUb0bWzk9NxzmIRP
IgesrKVsAg/ZgszeTTeUcftLaxDZvJr+m+IDk00Ldrb8O2JX+LUGzzOA9Uca
FC2DinNWzosVHsI5Ebct8em/3jtWubsrtQ5aqeEL2f6/pmrUYZ3Rr5wpZvv+
eE0t7gNstBGFzbz2BElFIrw7ustxt381BRjLBYu53rv2WiJrQ0jC3u5kLK3b
dFXttHIW3Lc8mlQ0FAn7Et1BRWcJ/0MuVx+Pb0bkIYQIVWqtphkm6AtOmUvD
4Y7Eyue8gJwPqhM7/L0tfeCnneVwnxD+8g2FgR0Ut6j1vsb5qXNvvPJ/nEJx
MQe6d66px0rXDS5Ott9bmCEVQY2FuxKlkArcpeW+MfV8H5If3cUM12JokJL0
PiFO0NQk24GvKBFIJZwixgkoEfTsqr97KXajHOCaT7JL+W/haKnvEApj1o/X
4edDJhjbBEdM6YgjWe4xb5X7PDPFn0QBO52/sfRhGbSgEONtQm8inaxb8Emy
uataITNjTWzzxdMqC5oKkaiXBaFOiLn8d2Ow7U1LHomdOVn65HU7G7RM3fqT
ANXdIiyPWUmS/xGrln3hJsrqqukt7Ghw+HVESbPbgDehw0YviMHoBxORk4sN
e8nLMsGVQzhlXEIIbk9okZWvOObd5fIm6E7ziygHaw0mEtwXkkn3ZaOusLHb
bRH4gh8MKHOH7QuISTHp+Zgphpw7bMSnMslln2GZdWL89J/Jhj8QorU02tFe
+QZdBi1kdS5SpN4SuRq7xBLpA3rJlCej2TeTluYnjB7XVR/g4r3OcIZknoSQ
BDe9NW5qGbpKj6CnCnCdfqmYI18npvN33WQLaQRajQSRSzcFaSBBuVntHW+5
G/dhcDjPxfOWw423cmH1MixuY8l466ZQglcXSrFiC59Y/YDuku8YaQMgPehW
3Dti4XTOscUlDamb4t2tZlawEqRQI2zICVW/juRJXKCMCphVIm0uclE/kb5Y
yjDdGnyPnT6jYC7h4lkl9t7vpVbxc1Csq8OzgZWY6yf6lVwkOnqyy66JBdLB
Qw2IzScNkgPxL3pCbhgsUDlQrkQDkGnQQoD6v1W2HeZhkl40DTCHLznpRmsF
Un8d58oxE7gg1m1B8brlLA3LYxVOngOJLLs4o2zn/zegvRmQUmjiOvlGjIFw
Jgojyfx8OEX5cWu2lcaM1+wfNBOZDLTADCrjeEyycdsr6xwgrJDxqnXi5BRK
UURgQM+S6+mehGkDtKaYaf39cSl2jWHaMGsj7QJbQeWvGgFR60raKB8oyYnB
O1cNNE0VhU7y4z7YDpMU6kkvIsFdY5RkzJoXdqeTlnPknA0o017Jm1JGWQDq
X4KEPnlpKLeIcrj27ImYiOhIbckr2Qr5wylfqsfJlYAS8r6y45PNfYDm23uK
xrL3ykKJR+wxNRGzp4P7V3rtIWrCZ/Ob3nnzdwUSIWViLjPSuoR6R6uPDSEW
6abqjp0zupO1E5khjZHW8v9+J/QOaopCYN8qLK9EKkpQc5lzmse6cWoRzPRY
VHvYkDKNPNQGtQUXhes3a1xm5cwgyDDE3/UY8LrU4DoaDaGYlb2SMNAzSpm5
RBb69L2gD5mKNFyMOJOmOLWXwFynjGVnB76bjtRUga8e8mCasxsawnJh2MHP
yWVGDWQpranBJh7qWqtUXaM7j4K/DPXuEfcK36xo6Z9RT7eiXJt1CShd4ltN
YBbUMJWqdvKO5eMvZh+yMaZBUdasOLzSyAPAMVuuiK089u22e+4sx+DIcSXz
fGp4/50mj7BR1tqqfKxaAmI6aJ2dnqkimhd9px2YF8kewo4yb3Iq5J2CjQox
gg5XGv0Wz+lg4eDO9q7p+17ZigAMHfpf2rVAqZuQCO3tkJQEg4DlzCuqohUR
hc4IhU0q8zuqjkuIl+wIIWJ5KeooXD+vUfHQlHYOhIu4DZnxEwoqnb2OpLqz
FdAGYjnj4TYj6zrMaG8KZ3NukiwO6crQmgnIxi/D39MWcMntBs7PzPwOFWPK
5CSSXBJT5IN7rxYmiGXT4dLdChlYkDyVej2vT0iW9AK8EuivdMCCOnBv0gr8
C+1hTr81glUvhdiujrgwuZMULdINOY2RVQ8mfk0hwwD0iHNBGipOEdDJjxjO
B41Zev7bXlAA3QxawDjsikTmYtauD940pIYyKfSjt0rdpGR1X/uHNbHPXW0b
ssfdg1hu6gwkes0iB7jj2E32bHJ2JESRPCfCDBhh0KGUvTr3pIQcuBCEJw0f
qXOTCtOYROiYzEzmrfqtzj8KuL64Ze1KWPZ0NOAUbE7Z7huekqzciqozvxCf
dy+wELSuG5Ov0Nk/hbY0WpCax9H9JpEY1RgGvbqSJjZXtHZX2tIIhsvIVMga
S/TN4pl5WP7wzh7MXOuSgzhGWjAvR9xdc0hV5AfLocTKxW7I94IY060MA/hr
kgqFdsx2TnSmlAJrs7UecbqKLqpE8EqNSEgsdp4ZKlEaJW+5OcVZrtqpoT9P
8bm0M0ZghZIHyNezaQeFJ8cgoMgxG6/DGzQY2I9Il0SSvuybsiCB223806Is
ZdKBJDwdBXDh6YWQy2Yk/p3v5J478895j6JG8jVfoKBPJY/dc1uS8b4mqYV3
t8FE+9jFkepG4DRxJ8YmDGXoeWhZPS//8kCtsNuTlBBJjgE7tpWsdxi1lhUX
dTvuOvbxEo3WHXLWJRZnPMQylNfgKS4gamyk6qdioYBMJqZP6bGIbvNWmrjg
IvyAeNe0HNlVo5R81TD2HYQ4I2vSUtaJvgLI2qlo64Es5FcWmJ4X5pX9a0I5
rqJzX+kiSZv7kWOHDAuLJ1OCJqE1cuLv4lQ2IgMQGCmRXO2sPqVYA6DxooBq
PJ3yRT9/CzK1Vw2NqZYuc/4j+/qdYpd4z3yFdg06yME3pqzTLd1BDcBYBJpz
aQXcPIDUtsgqPNWf8f1pb4Pc1CpPm15z+6XMRnRSwHESVeBzEBZfK5AHDKhX
YeISmrq7J9UV4Bfg+SfowgmQ3o/9XiJbXFMvyr01iO4f/wDX1HPLp10e7WmV
Tc1kTGRBmjrXEBtUJ9NSvAG60orBdpCZ6iny3vhvvQkHJSSYM8FKNmK6GUqb
VZZ7EXu+HDJg/BRlXHhPQ4xYVsYMvpGLPYv8DeLdOW/wLrnHxnp1RazjPoUs
iQDip/TtVn5wqSPG1wQ3uTDPHgc3BLXmvp/VR+C7z0/4cCaYtYHZy8bCGB82
lrFzQSQS7VpHYheuTxEpc5ICHNEOHo/e9UD/1kKszmEWL+DGEXG2sxIx7uRH
6uTBPNvJWOJN7SecHnnxk1goYHfcH0Ygu5XCT8Ad6C99zJR3XTPZs5ESF3Eb
fV+UBEOrnUhR0+0VHAyx1Vo5ljghL1H6HtKQjNZHQ79y8Nr8Pd6cHTHZ2SXh
Xnr30i3KrHw0/lYzTbfLOvUzt8xEDwWpNNcgZiiAWkRz+EjhQn/dcaFhUSpA
BiQZy7yJkGXvuf7NcijreFSMCA3/U2QF3RdgXBe1aCsaLjL+VUOyLi0GFDu1
93d8b9Vhj81OAjABMthnFxhy7y0aAlKTy4Zn4GdvzYHyL0FbFBHANXUxmro8
330hQ0vphnIK9apbis/yvF+XJZwD01UlxhI/N+t8sVmyG3o3kPV5gezOi22c
2ELhCAtzrx7Uqp9Uo71X9sUlFlcgz2V+oe0pIuCQS9WdBEUFLhm3wjXOqeot
uKzxaTh/AusxnIURC8+ZTqx+lDFw0v+2GNg0WcwWGg2Wu/lDW19rlyWvxVCX
rkM0gKAfq+56rMGUON6JZGuyF6dnroZHiJvdbcgHYldHSRxpBpdA0gbwCxKg
M3Idycd9upp3ExBO9UhIwlO4DnHL8o0TLuCvIE6whA5lp3wUdZjIpo2kdJfN
Pm92RSgD1ghvrnmOD06y/yQOydZ4VExYf+u66livaqbq7pX6qKp0AL9hipT3
G40jO7JvofJ/NNMnvDKJBK+P6tyfQ+3sLDkHoot77ZkfshS0i23uzOBIEAZe
4VvHtqXIGcGucWAlFsFXT+h7jnuFCSBzPQWO8pvOXtcTtWvnRT+1/AlJnsmp
FuHzqZiU+/Ka918avP8SNz0l07UpkmofsYcPT2LXhMFoJ8vlO1vlbjHiJylJ
9gGwz5Wsa4d1tSGs7R0ehkbGMivyvV+dHEn+px3ZrE2InnHO0SuuM5YXkj4I
/pWbnM/0OgqEIXn9pixVZX8KJCIJokuO+8/our1ofVDOVJpVwqTkYyjt5tH8
ax80pvtc6J/MFcem4ykTrHwSmjx9eptwjdDTBpYKh17BC/Dmfx87VyzhJLa/
EUQTCRNd/SMYEihFb/butQIKikqAkDGZd2Tv4qpj5VYG/8ICFG4DR28Yatd9
W5Rw1uDvuXFtdCFNt/Z7gEQEUEKWY4Qt9/5bB1UDE41hYzTPPPohmzOa1yVS
wA2LcMNMbwOollEg/EqcsMKF+emvbfruN97Uf5iOn5sop24F4tSdhwjge8Gv
MU8YkacmRrxvjLc402kAQireeL8qqf2YhPj5V5C6eeMPZ75l09VP+r/c+M/S
FlGt3xlYHet18Euv+NLghyWnD99DRc7zUcJje7lLOdlVj9FBP1Vwy59Za4z8
G3LGzUNlLonOfVcr5YWBuXMwA9whHmqKZriyx7Rd1bE9JECk89muV1HDyZFc
1BBiWfo/Qtonu9wiFRap6mzjN2WuwRamzSZO9plaDAykv+HGvpw7PavVJLwo
Riyjkj5zgN5NSzqMz/SFz8saiJ5QAAPB6Xjl2h1KrVdCbIjyFFH+8e8BW6xg
Omn2odk7tGPJoQsO+sd7wqV9F90RHF/nrmKu6By072mTDXwmjHeFG69TGqKj
x4mGPZ//xWozpLxqD+H92IvFUBl7hyf5H+1AlYUFGnPvw/q0ESN4YiXliX2l
gSrQ7esy2uYpy1ey+jo3EBKkN8MtC7/sdpKIJg7XaPkdoBTYIFzVAjqiFK/t
aVdTMei42mnBmXB7YEmjYYqJWdTYLJis5dszTe1Hp1K+4XDHqHO6iqZZqG95
z8LUZTkNUckmRbXwpF0za2BtKTSqUZJ952TjAw5xw/aRzBTZAw3CBFZ7Foyx
z+DvXN+mbXL/P6+oBowobTu3vBxinmJ/vJxs5lFNtrMzumpq4xajlIiGCY/l
YHxRoWf+uYV4AVdjs3oblvHX3ybExZbFvAuJyTxfo2+fu+f6I5OZ6GV32hi9
tg5MVKCUS8LVoBEOscHa/t+adYZ6tJjVAs1xbjmuwcuHBzFE9D8joh0y5+34
G2KfolTzxMnE3tqUjXrO1LXnwlqB3hB1N3B94bj2ONKZYSQiHWW31xmwDCkS
ygakitS/sC7GwGbfRP/itcI5d91eX9u2j1pYz+BZP0fMyARO9Yv6L/0GITxY
kHPZqHmiTMfx+YTf0Zaz2d3l1Ug4cmWIHUA=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyKBU1CjsoZsgIFpiSYTsq7ICHt/ZgXQm+7S96Hv3977JrmWWbKEipt+5neleH0b27oLSrn5HFMD0oqoeK5LJxOpkj5Y4jW6WURvj0rfnlVQWvvMaJFjoVT4yr9W7kFwC7LU8aFekYHf54/RNFuSOyDNHvpEjsegywYoOjxChY5hZ4GdA7zqI/OiNBGteoRCD0SO1NQZ69bUPW+sUbl+Rzyf6xCF7mVZoy9mt7neHF5Aw+vgcTL7W7jwWYSaBtT5dGfgdLl+qzhRR1MY6ufSjQs6pyWh5A++x1sUtdk/89PO9o4WRoqfMAbPuTq9ofaonsTd0dJfdf7SkAgAkQgStKPuIfbdtnROZUNn1pyxQj4NQm/fppoa2crcSEsbDDwaGB1FMTYR5nuwjC1RZzLTfaFB0h5OXIMQh+/LsibkH9wnbKJvveQwp9ztU05QmTzv5JXgQIVYHpyZg7qls1sqLJzhvMv4b1aY1fhG9A2VPlcsRFSOxL1YQMGXtAAR3zyEVENFbn4OO70Sf2xzubGeKt0y6fnJ5wv13kuabtEWY7iQTxLZqPHMBJzz4P9/TS7MI3QICKb+LlWk3nNBjwU7WIHrRx6W6wygvGYfabjNVcLT1R79fwaZvTPZubqUDF6TT+75kq/HK7Paqu4YUU8REAs0Bg/TtzyK1eMox42/uFN0x8Q0shbRTptHRwv0CF63vyrSWzU0aHtqkRk+KuQ/LmoZFeTNw+yi7Vuf5rBko0HewKX3BVWP+sxgt2E2r/OwR0BLzJ1fGXbQBYii2Q3R4mfF"
`endif