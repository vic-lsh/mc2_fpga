// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mCUjjBu6dBZDhoI+P3sw2PA54qqGoYjfJCjk4an4NXBbEaEfClBOcllYEc04
0JrPI/t6mlmUSXfdHv1K7QW6v73E/o3jWtNLn4sPpVTGdlo0eFVSMC/1rpp3
UmYIAq7N7l6kGgyZGOBo4s9/PnaW31gOjgP5kfUUH5I6ZPGzdnRxZNkNeiri
MMl5tILMBQ4BxtCC8rPhJZg2d5P+KBk38ULFhE28tAqUvhOT1aOkoP33hTkU
BGt7Y8qiv0tLywB0vr1EFKc1/QlNd2fij9E91YAh/MJMrg7GykyO+csLu45l
NhSWaTuFvhvg6U20Olj3CzMLg4wrtlvOOAg2SRf6eg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TnhKzkRVFAzv7Tv+qXicRwWA8NZr/lDwE+K3689XDe1SvCsNsJxXY225EVzr
QdJoXu1u5DrkmOcksMaXw42ri2hY3UA0R2PdlS+LQAkuq4C0UZkniLGCAnkK
nhMA0K66C5BabmUz0fjjfziC6+ioNgE8syxL9/H+o8e5016+MY1npxU+asyC
XXQD/EPV8qacEYck1bB/6UtDzfwUuoDoxgjdF40rPoSzojkIq27il6JaIq2m
BG/jNft4h69aJO331Fybj3tRDbFPbqi2MhogGMTiEDljXt7cemq69H8RD7x6
HIdQ9mF43akmWQ5dbY/j3m60/eCyRrCxU/ivpUnRXg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fAZEuZoe/4EURyO3BUc98xSFyA5gxadZ3zMWjVb6+tBlmnEiHj11szsqiG/u
gtj2jqqX6c5JHokIah1JXGj/Od2aCF9dOfTYkcBAYMFzR23VDUzDjDDmpONs
ZA4nWgczhiDfvTOZ4zyi8WJsWO8DuADl4+6VeZlJr+KSKORbqddoSJQwffYZ
Pe+v5Tl1OWiAvWSal22JssNk4MmPY2I8OT+iy+Ad5I3eHheLSla3NmsENg8L
ijqnYx3KyRjUfxkrRJbzHAFAVX6iiO+R/UYoK0GHA9bqff7bqSbSIWthfBMK
YhfKFts9sCXSg/E56xsOBbbwzcooo0KBq0F4IXMdkA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
loB5n3erErILGLz1Wc0VlvrJCLXfuek3AMrsll1/1a/2f/LqfLHwK/RiVUhn
8JwxGMqX4b/pulXRozPekASXhREfosIutWKJ/6ZCjS6xwGyne2e4HsGr3uMo
hkdq+S6x5fNd6PtfA0YBXJIJHFNGfBwGpx8Mutc2IcDEICpHAibbmqmE96y9
GB2tguNuv0fgKDGnD+WINSMbbLaNR7dRUU4J613f0PKnew1MJ+WOcZ8tcmNR
jQpARVtY6iosV6rsPlAzmoTSIHP71xvdpMaiplSx4LcxC2VBqOnANw+5KloQ
k3x4HT03P6joXxxKs95fHQbzU6XZ0Hn7TWXvlc2WrA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
q4ndJBfZzhwrSbL35KOHGlPgS1c0RY/kjR2nEre8K9KSrm5W6/mD+4Qt8Muv
YXUVycjyKhv6UmrrVoXynq6PsT3BXqyQ/cU9DcG1fQRVcXnPdp8SM5ub+EPg
ZvMo5hI9jmfItNtkwQwglPQ5l05gV6q1JQTdis3ucgAJalb+RrU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
v9Q5+3kKABOM2a7mXKwgihUbn6VRpEXuhRSwL2MuS8dzqqUyJANDrXoSAB1L
enNKG02tP57hSGulzDvPh4U1vvq6cDY9m8AwCvGChqKW2RKZYXv2xzUlk1IJ
EjTPOauAwFVDeWpeFn6we7quTGPL5XkIttHEYlyYcAl/CzihdcQ3DcUMGGAX
brIZLEeWP7psdc5qLTxsE86v6L0NeKrmREYrY7GJzDLAx5gnhHdYdlx13h4z
9KeRRtxika09GurvIWULonQJ0qquwICm/cvd/t56DzRsjg81DGFKj/0I/E0Z
HVFl0/QtLeaLgPFvOSf/YxJU5bjnbnqf3qRndtEoVzlyZxpGeVtDQiGqEQEb
ZWcYtKtSczyv5kklL/Ry0Q7TkGG3nJ2pOIf7cw8pOVI+Hc0RgVBSbh0XKaGl
rp01Nvm4TQXpfFEg0b9AMuqMaIesXeaXIUme4sR9FI7c8Th8DGX70hUTfiHW
GBFwi97hTiU4eG49T6zKnANVgX5V7FgK


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qhIfHhuBNYy1MO+6OSsHs51yvwba0shFE7elaCjUoRY+0Uc7brv0KpUv9ZWv
4qLlhNLMCyQLGUDEtIsi6mg9Yq03kw0Kyfz9yLyu9rmD+Q1V9DZMcuO4uI7X
7WlLS2l3nLt/2BEH7ubT3l3G1gss8FhmepNmJ0hzAp1aFgBtqS4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sx+gZuHsJpv2+8+801MIJo6Pm1Wfw8+bPohTqsGNwNvIub2sDyapm+mAzhVn
3L9aiaVwBC3U4amTXA2+5ZRSgR3t5kA3e+0/r2S3XpITw5i4Fd62x8nW3Ub3
HcipZ303AIcUwflSmnCYzWTIr5DRYEDfrPmG6PZhFz007K5FSVg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4288)
`pragma protect data_block
LmYcAgxOhUsYuRxQPuD8rXZHR54xlGs/IArNS3WoxR8CxGgUIpLTwmbgQWgq
5qyrBvaZBopMkrlKVeAl3TnlmZmTqgNbcJAriiypL5w5gz1hefqJk1s/9wqB
RBDluzBW6kiugtwrGd82yDq+ZXOrjF2CxEzmViQKNF92hqaSRnADsX0JeOVL
C4igt4V4YHHqs8GVfS9FplchiQFsRIsuQOyLFuZV74DfE3AvGnvDMkCrfIOY
TkPaQVByz1y4YtsOKRG6EXNcXvOgPN4SsLenU+PcQZdZstcbu2WRPlwl+kGP
n3sRBzdE0bvMnZcYvy5Q8YrRV1twtKNx4+5QS2fbkefFsyUBmNCSID7P5OOR
YpOiNBJQgQwKcHy2asRuMrJBIXgh6Z2rfHxJE6xJyzNTDytBlMWme5avm6JA
C0JWjH97P8S1fvZ+yYSIjl+PotMBUaE3qMUNvhH7Gh9nXNe9hWTCviLsbOcn
3WGl8VqjVspZ4pbsfA5CrmzHuj3PHTaTRJ0F57WC64zu3pwknhor5je11GP8
QCmk2eDTcafDCN0sxZUW/h17JZjZkzfwOazhWL4h1ndfKqsHlbeAHtzISCMP
Y3YvdRxWMQaF7R0PAfqFFvYYfDoVPh72UV48JSwXw5ftd4lICN2uFxhLsF01
OkuM7uLkBRqIsqQ8d4+YCDt+pChpOhlyQNF5fbONTaBbGGPOlANo73pgzjfq
NqEZNQzlMW/PiS+g/DkeyDroNyytJar+7xVG/TSmXFpJPmffv/b26yjtjrpl
ms6pM5lCgwEREaHOjmetcZ4VZM5rcTRa3Tm3qaipLo06kn2oQozR3i+NRk2f
ZR90+DEN3MIibBnw9O3uE6QiQan+/1C4KiS1VhXaL01l6JFL9ZiJBPkOFaUg
mxWJXvrU7T38ZEHzeNOnTGFRzJGf7WhY3+WYxI6UhzBD2uk27xlQYNPKEZ8z
sgb5IKJq/gGcq73aNZi4zRdpEubTwUkhMu5nRMwwnQ/AhiOrBJUO+6yKqool
Uj9Okub9qyqCuLhDt48WWXZwR2x3Eb/5OKRzL/ckh5YxMZhcGdk+TC2Xlcvi
Pwnj4cz7F0CX5ndVO3dzMd7AO2B5Ws43YeY++opuIBPNaKqvDlPnZnLuDLvs
gOWEOCMd0y+42G1LyV+mEPqgDfqApuZ1Qd2P/9P0UZlokWiF/BgnO1HaG7ID
eIzTXt08ybHTiMBQLwhagaSIYvJ6PiGCNx//M2t/49qnGjFcdd/w82mgCjAi
pxlOTPtWVcIKrhWeXQhOS8Y9tWUcFXm6MgkNj/v+wrHborbMmFWDkVPU6ctc
xMVMMwrAHkhIvSzr6ruAJGiXshPWZ35eUnD3/NJ1r8ETgnV9P8fE5woNNQ5H
GxO1ihYVscxcGRR73jmwzAGE9cO40n87+Utxp250fX180npTiD3XO6NMmTFT
CWBZqamiq7Ucv+CH2/8JzjGLWihKAIM73Iqf7FvNL4REJ7pA/I5quY/fSTVL
WhEWG9JHDgxg/sH/nTB1qaGwfGzG5tmOBmAoSNhNzFQ9bSEvUvJA9WsQ6pM+
yjX5NyZgsV+d+w3BUKsIm7eqpYQa0i5GeOiHS7bz2zJWC3kKdUX9KGKR9yyp
nYJ+PtDCEBzj2nLWbE6ZRZIAfdNOsuB5/9Rx2IGrrQO+KO4ED9rWxdIyiKDs
++mJ2hmPwZBFhrO0xn+QW1OJFkE2NJN1O4rlFc7w2YEjRe0YnkaRFiL7k5ja
5Cglg6TofCsf5i+KLAkre68lIk13uaR012tr4N1u3CUTIdJHFZeah7xUWLFk
XHC2HV8+w1RVrRFFvfMlKmu1YZ9v46MQKZgfjUlEmksQl33crmFFQK929C8c
b1X8cvZOwRL1BRgu8X0Kx9fEmrDYWa+IA7MktiUFCP38a59cdfZeXMP/44CM
FU4numZw1MQSj3ZKmcrVai5zq8dZL9jMYTbu9K35oDrDwySV7I0penXyJ+3l
APr466NQi/XDIw3NY4uG2CTNulPgnuNs4U/RlPadsX81ufaR0982v9hcvDTD
m+m4AFt+sUBL6TBu3GfEaEpxtPhN7pyq0ddG+k68SCY9YzERhNJFwK3dmjci
u/J7PQiOIyXUZRgrN8oyJLXTmoEUmyFTvENPpThD7kwtpc2mkOS+sr27PSb4
aIcWLQGYbOm4n//IDKpZ8ikiNio+ElnhhiIZuonpWYuGdjGAujdkK1KvqiZ5
Dk4RDfWtVByixGMnKE/BSbRmnkvGYdSvm4UpeT4hb3MqCEF61HSEn6MB4y+y
mK34uK6Hz2KdHK3b0nHIX2mzpOgXuvvP8Ro/dtcnX79JX7sdwV3Ra6IJLptc
3inCQ6j08IY1/SXj8nHeHLuA29TlY/2yGC2cb0o5t4tpam8LCvYDLQDKff9C
kIsCV3LGGjX3h+XazyLTQrHdIxCJSYFerEvS5G5cgnUlTvEHOjst/i87FjeS
6TZbDhrtsY1De7x6TMGs7IcPXHWhazVn14ZNGCCvbpwUv3VdaIFSN4YlXe80
Zx9+dBpjvN4g65LqGsVvnQfeamf41EvvdMeuLhlKOLugRbykRutw/OWfRc26
Yf6AeZouKELrNU+ZK83/gTo0XeH+78wyGpaRJo3Guy3mvpBaMKlFmAKBAhF9
R0cH3M9K5qX++dn4NPOdExQrUT1WTgoLXh5G8gm0mJCI06mAgfHhrAV3DjBb
ZFJUImUNjqPbedeCyPT1mAdN8rpXaes4BcTJfccytQAbC2C8sDH/b/bVNovS
3Ehg4SrO/+i9PqSX5OuyvNpTpRE/+y2BFw6cz+633KZTTBIquhSPwGzeeF/a
2JzIg/ZSaCjTFZGZddAZxs0bMyJAl1WwayO8KhWQEyTd5plEmCFsKhCubZFV
akHMS8eSvR1ZlFjI7FKz7OGnxWOW+Eptp1z+YIEeP0w9kne4i49EIERU7y66
hljYhFDVplyOOeUwe286I2LS8o7/Ei5Hfryv6u1Hp9nXLu0hkbm3H9HJFw6K
HYrA+IIUVYdYE2J9+J4a84a8qmPesvQwkqi2DjjQemigDsoavSQ3D9ZHEzMo
HMOgPWIzSRkRx7A3yaJTLTM2iEpqfELN6tY5OcO6I0VcI6SOT7ciRA9ESLQu
JMiAviikc7EF8xBMjA0oeJbDjfqr7HlT6Tm2UnRZP/wNshX5RyeBDYUC4oJG
dQa+ZE2ae9h++Am22VGbXrEtswVUvkwdcErSVjs1RngLVj9CjO1IsJ8l32Mn
gIXQ8Kma6S5VHQkn64JD3t9qKwtlNhpFxfuB51+ktJqbwQwtroqx0rwVVKn8
w3Z/vN40FD5a1DNp2w03wFrnzJG4bNWl0UBYqeDRz5veEkPxg3HQjbTenRpf
CjorqofXfPZhSwerMpJmKJWIL1E07fK45P7hkQZkNCz0tYT9gcEsJP8j5Q7/
FclKhWdp8Ezi9caDJlHqxMRr8ugjoX+rivGhque7/jVIAxkXQ79hjFG/2l9S
G3GQB/f1FzBMw4ftEzf0kaviD0WW+u5h981VLLn//cN3Vwf5f84yNzw0jf/f
Pg2RnN6w273qirVcGhQTe2bkdUkjcLslm3RBppIokK00ECs6fPay9ZbKMcfs
DAZw6Vo8mssqQbRWevNR6gcA8aumGLCiblAi+1Z5bHVDQNx/QzZu1pTmlyNW
MbSYSNQ8meDHdgYmj0qfcp+LHALzoNasDmUVpm08rjmL21ebqhnj2OOt2RFl
cV9zfWGKi2WPt8+ZbfGriUXJ5bVQSVmT9tdjfU/FKFPZ3zkBYyHiE2LZuRDI
lvAdSoXtL9y7ZddtenilSRN8IBvoDdYZ0WSX/f/vWwFGBPMgW9mfVQjhaGDe
zTflRxhBSChzKcz4OfXy7vVI/VYVOMbi92yDRM4fuR+12jQJccO18LqWF8G6
1EAvF3b3d8wBXCXbA6IwWBUH1b6kMGnu6zejsCXnFj80VG3ITOiXSOsEAe3q
zAqs777c8jD1MpsRE9in8kiww3pVImauZ7TGYDE8DObOdyhAz7kmVIQcgMAu
U1Xs2WMBNGxTynXaAWi0o08gtI5CXJiSePH+c2BThVBQDqWazLIEXVwssxgX
9iJMPomKwQJJC3ha5qdk2tDHDo0MosJE6vIy10xlRsHoH6DvBCunXYQQAG22
GdCI6t5smx5OxneKVHHWT/hBzI4WGfSLsZnjSBAv70/2zG8BvT1JNL6cXVLJ
WQxRlt8NYZwAl/EHcNC/IAQZvSk2dh0yx1ivfhNU6sIqrS0dE0wQQc7++kUh
z/4benvA+feHfy3O6j88VmC7bEMLBAgwSym5SYTmH99X6o2xuwLo1fnsRrhJ
sdovDNSMARvH24hXVPAVOMf/YdVSoHgvrkbSz9dIWpaC3u1K/zxCGOkVqs+t
vwQlYO/PZGsbW6ndNw10715FW18RaEUhkmV0PXVzANzX8Ub937e5v6h4l6zf
xetX72nzZsWAe5zSQXBo5tQ8c61ceD7Ejl0J/kmDACpUFqktnZXRGx7sels4
AOtD9LLWuY0+jWFUCNQ/iYrljXPXjoN+VHUAaziS6ZOpGu3qkY27ofrFnp+h
nh9XfZNi/+SRLJjkD1ChMIHbWEqg/CYaAemXuEuD99MXUcO5ZEyWJxA++4MF
1z2GDu751llBe3G8U8BwNfLxJB7ZOeHon2xfm5v9HHJUJY5aSpXKErWjwscp
D4xF2waABzcTiK4GxAIsw8bVnB+HEsh9L6qF0htYM9rAubzfPCzs8++RRkw6
pNBj3czrkP+zYg+2+tpJJjxWeD0f0KzhVz4HXFx/smazCEQIa3yDb4VAm1qL
tDpJ88C9qSxfzCdc1DDqE/yZywpziwmysPIRpo0qvcGWm/Oc43QdOg8pVVyG
awSmxqA0JM7IMgtL6UZiAQh1/u2at2Io6deK/+84iHYeTgQwhv5JTlDVtmGj
WD2G5MpIjrt3v9NErI2VOj3F8YeZrZVmqMIa+1Nxv2I7D5um5tgBc69/QrDF
jS0bpfyQLD5HPONaeyNAmkkon5bz8oYp+DOJgrqMp5yIj9Lc2OVsBtVEnrBG
CvXQTQu1nX44/d5XWFFhoNVHCMull3FGd4gzkx46swkFiOGYwYa+jdVoRAHm
IePetuNQgAw1D1AuQSKhouFuFB5Zdoq5Lj9A2QfS/6noyDlU1KrbZWuJBJH8
sT+UzNuZ+el+elVeh4lxjd4Kpz6aykX2Eb7Haiua7k16mc5UcikZqsc7nch3
VXTsp0SMRRilC0RoM/0+LOTdkECH3qYwVM93pwHqpzi7cXAGVnwdLkgOv37v
h5o4Ceg3D0cvQE/sze6tH8OiEzF3nE2eXUjQak/TG8pXtGdX+uLO1n2pmi8o
Z/9YsLE4nXVR5E8NUmgWAEakun8/EpCkkOPluVyGsBmdQ1/d3OUmbVGdok2B
MaA1beWjM2yEpaHt2dOmsWtABQExtwVO430jmDVhRMjlTt+6O1nY+8YwhKkz
18ZUeBI1wiSf4ccfiy8RCkB4p2Qry1MjDlqqffdx2XnWM52KnHbTY5mw84Ph
eo6LDF767Nn47rPbtV8xmvGjqtRX+22iRSv7ZsiEC9r1Rc1LCwWifwf13qCj
c88OIo2eKucMqUJ1iA8zP7oO/AE4A5Iwvn+2q2tICvMIUknedhULPZ4zn6Ev
l9G7idVf7j5+QV9WqKsCPEDKDkYbOg1Wle/jesPFHM1OaAUHMWB00OZKU4lV
ktgREUxRV9e8jjg1LA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "lK4MM9NDeLrdcSiRM+VIuNgpOLUAzWAt6nzBJ3Vw5tvBogzjtStM5gMJjD6PMmMyupOFzYouKIpJuOZh/11WnQBMmqEc6gvbtnHqfGmxFaxYyOv1rddc1B279ac1WEgUgi2BHG6DRj+tHk4+Vv2VvppW/Z9gUZ9e40aCxOYZZHwEVb/SJ8ximgD4Fihl81LOgt6U1JRoR0S/yAHMZXIkaoJ6FVEBkPAD3J3ew7MX9EzJcfgHsyessQd5Idvv87A8Pfki64qHlo7nR0YcnvYtwC7//1Xm20EfXZlKQFFrKGp5YG7/jrcY0gult/ltjEHkmyUAjbAEFRUtu5l8omwGBz7ZlXmUJBW3BacBlgzbhJh55oE2a8sJZPiJPig6QAa6SYztQwlYjB+xMKCoZWTpKfvKVtWW/PRH3oLUH4w/HxTzoje3fqlc5FcOSTJ6iTkMdUK9Jk6+LL1EMhS1ZHfUD8SdE0vA9I7gwmA0l5NMs+IPVZCMm3iRX8kXsSjxzv/YhMCbkaB+uTlqezRrj8lFq+ilD0exwsIq2NBEi+hm5KnemNuAJQxNv9JQaliqCvhWNqJrlNXZg/npf3tabP466JoWgc1iJl9F7xRr2cZAHM8av3lrB69Opjd+DCSrmwJ4ySYOjic3QWjnGpRSOTYOEBMWWAHdYxNTxO8FPbjgsulLJy2W0TtVx/YXlqMOt5mUUpxG5ozCFU3dWUuE5Gh+JrTgpVBM2vY6efGj2tviGQjLXuo5iBSK6eWgA0LR31WxlPWz3DbeVMOC1jRUnWX62TH7U0T200yXTC+Gk8Kpdb4TrQsAEDW8M8emNbKNrEJzA5/tULDPC8ZiGWlolaI5fJp0TvDhHmNT3IPY8zPK6U6W6sT78VcgVkpLpzOzPTBu6AxSafMUf9hchvkBHze6+XUPIBIC0FyabQ7qH3M/gw0dedA/tq3yJd18TDI5tZy7xDGujQnYY87mWnJjfuMDoFZepkNrXKVgF9gD8qqNGHkgUANAOYzbIktWtnhDCl84"
`endif