// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pMaTwjDiO3Tmy4TRtNh5mB05kI5pzBGmvWEkRU7PsMyIEW+aBELZPjUHbH9V
DxpFI5yCyoak4ld+1BGtVujplVDd10Vgciagou/2zDeyAJ1kokTD4Bojsq0p
kaVXj0KGnVgLLiuGQmuJQnDc9xH9IWxQvbWVh/A3IHEMJbTiVzuFylK3uXxZ
DfMmuV9uzq/Kivwj5wpwJ9MUEbOprkGLgqEUdyfugspZ08Pd8gfYe7BtYsKd
el1ZETT/SeRpbOpBwu+NfeurlQ4jO3vFA/Zb/IZJSrirvIumw+Le+qkCyoEP
OFYlcePPrQGrR0TTuq3PyYWVa1C92neVV9sLqHOZtg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dEEQbfqc+4PtKb4z1v92bkB1Ph/gzdb9UMILMLRCdl6ksBARkzk+fEc7tX8y
kqUioyris9Lf9F90kL8/0fHjOWO2liOQAsUFynItIWqHo6vEPBScmHVuZh/i
D/o5yxj3vTFd+uDDV31u4VIMpAWR/aDor3pttRTxQ0XaoqLi6w0gpd2mCsfo
oNEPpelnMXfi1Uj1VDnqRfgpq4gAmDodHTCUb0EwKx5dq5vIYuClDDIuv78R
/j2XsLqt0dF9AvGgI5Wo1qrr2Lnx2X94T+7s5dLR9SWpBfeCqKXmwvv3QFDG
EZh3Z8tp0sG+mGOnxYw6G1Efq3E1K7bW0xnd7bLwjg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
o9w+cR0X7OvzuvdAcMQgauccUf39lzzRIr033/yA4AGcaRyV3n4QGpT2mgVZ
Wc79MY3aLTsYyNDvswE4V4S77v/zeEh3e4/uo5S/wNInRyifLhjqEMwh1HYj
QyYq5Ftyci9brIo8mqmYS6w+WhBy8tOokUP1fpEcJyqbNeMTmnhKAg2KA85f
o6PRUW1+6AG2B+MqYimnm0mtdp3pc/HmPKYkK83hz0BfjxuhwvuQu6r1If7L
T4QZ2C3EMBNCCmwBW/pOlEZsl4wbIvxlyesjNmnI6czcxiSOtLkHCLwyWhyK
FnpJmkSRZqrrOwELagnQou17YWxA759yk0SLCy2bLQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bONUFveOA9DV7N9jiOQWeEYyJRiVqGMQk+nEaCsZBLVdhXdXxpKEjVMenwKh
PwOWezlXlP1UrhF0+dY3DpSEy3j95kxQC5euYicjwOi0hW+kdTZHedqe039V
/CFQOHPfu9xh7r/hTjZiXN3HSsvkM7JqONwoW+NXfcXbod3K2n6qjOFinno0
Gfmg/rHvmyze86Ow2FYJqQfJUuoFFqWjCXI1m6T2BacNu/WpBx9STM8xV7ry
RVO1PPef0kyHovdZqK2pNpNeGvn8YpOAMHEk3g0HFeB9+KNA52/1GCPmU69B
YJi0dsV51ad/hvPuQLjoejhp4+S2/CY29F6eMWHaHA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
djSItN4JGTimB212g16yXsvzH0Ucfv8yurLd/bkC0QH4RSfQg4fwdF6VmGcT
D7piLG+oDwDHBCOi+rXAB3RSCdZjIn7fffdq5XCpp+SIqNjltbwOscUwznaM
x/xun4KToG/HYBd5m1sPqRbqoizxGGQ7h9O6nF20qIi1AZvKNF4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
vSBicH0e75i1fC9k+gxngr92OGDCobjSHB/a21XjovC/B+TYQ+CNc9ic0fD1
c/L7N7p5THWaEZG8mPoBPyHGl2PxZNHWPsGsrCHcrm09ojEklnZD4riVldpe
rNOCK4GKBV5PzGFyY0xTs4Ib4SfOYdU82J7XK2bOdi1+FRsM/f7UkYUzLfKy
wdpT1mfN8Nv0eF5KAirsG+8p+jcGeUiDBCSUDnxWhi8QBhvAzWN6NuebVMfM
5YBq5JtoIPVCVLhEIS/54En3yoTOZHEUAJuxdOSb0gpbLcNC3o7rZ9Hg9y7C
QwWusV9kc3d/13n7f2Db4HBDQWD/diCuM53NfykgZA+y9Vm4JROH5Il7TZCS
0UcomoUZEF/s6fzqnVhg4mft2QdtGv5Gl3qkcGI6+QCorUOCJTjlE9Zfu7WC
ZPiajbXbTphIU3lxjFs5yam0ua3eL7AoMePhm3CJFeYey1cZo28VGAvnwxZR
SAbLGILGbRZh2aDOIiY+25aM1vB4PcdV


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dd8z4d7Su+0FybqMT9rX2AImecN/tFjQlpiU52mKiVOhzxYG4RIj6NWktrzH
CUPlb0cODDeL7IhegDvXl0AJYjNqDfQrtt6D5o3/V7CWCRF/2VnL6pdmtodL
1hhJy/vq0B5OTT8YVnGUnC+A1VUKTNXr4JfFh8pOzbWaAh1hD9Q=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZLRSz4+o9XZjXXi6USM/tWWNhZJ0FWH9zhM6g5fRiRA8EvCf3cZzCKrsqhIs
JizqQ2BsdBaXd2RLqY/Ogvm7iX/cGxdUAaqwM33miV7QTxBftZieD54OIE93
5TkQOtY17FCurME7BbcAWjTnryciQNKNbEBj38EP1Jeir3TkZ58=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 27680)
`pragma protect data_block
vVS6KdPHkuThhk0Oj3uyonpmwovP8/yp6EM6rpnLIlWgCnOr2B9xNjovp2N9
jmwHL48/vix6hLfhEJRX1Jb4I5lafOnujVCGC+oazJLfWOZD6A43w02QlxJK
BKSKWaQwQrm0cudEfBDYDpZQgJEeEgxA3yxiRAyjcHcyg4gEcLGvzTjVurCn
5WEgXDHLhfs53hrzoqVBR2BN4/GeWR8lGCDUNw98cpH4p2lC7K2nHENfrGA2
Pno/nXEPpUrgjmkyK5YJS0jZZRvJ410fj9e+a23Sd+iXaJED+R6jwijAeZRK
KojzYWFUBMHDKJAlgWKM+nzEcJ6VVJ8iAmbs6spiCS5wQAzE2kYlYi820oJx
thIaDQmRRZCvGZUs+GRAKvVAPDWpqJTi90NEv+czfBax2q+wjmHXEVrzZBVc
kwPmoxCwdWvozO674MIx35ZI/kMFfRSLxmAQ3NgXPbBIkwY2/HU08y5GW+Xo
w4ZxL1JdDrsK1VJYz14N4k3/2qyCJ4V5w4bmJ2rR2RNCCQX24//mglSM59Yc
QQ8CUAf8zY7Y+7auMhFGtAfIu4BtkEEwQ7itn0WWU4N5GPFUH60mvheYy0ka
I4sqz3UhVh4C80pcQpyaOruT7/g1OE7Y6teshHNlzKVX6lc6UUEd1YMmeNFb
+k1LAnCMobkQKqDYU9gNCE+5IEuhEuhU/ybSPwrknVufvp1Og3TeoYu/Rt+l
yi8pRMn/FX4Xof915wBiZc6xM5BMy1DiIeU49pTce7lT5tPJ3TrDDr2HvUag
L2EtGgVk80HddRAfQa7PhJGR0LmPwcpP5J0c6YjCQ30hUPjqnPnRselgjixz
YIiawyuUT+tovgHrjLPa2DqK7owoK9lwopySGmPH84+Kb8zPVW9fUOdQ/ZJ7
JCgSe2w1I6TE4wsUKNNqoXmZEiSAPDE34uDZrvTD07zT8C2twDQhWf09Inof
iuzNGvFwy/gaqNAK2NwnuLrJU6QzggUoS3CM3B8YLS2PgvDSi6elMrsedCfK
mIm+9Sf7LnQ4PkvOH3tnK35Hs5ALufrtQBH5H9kN/TXoETKNZlNGSuFYv+QY
PTlB4spoOpl6iFgYIZpsQbAWs5gniLqQH35UCRCPzWUGP8MimSkFgv5w/OZ3
Y1Ht9Jw7Kyf8Bjgggr+pXe428ixAHyiUE3PlftUEZvUVH4iQs3RRpwn3cR8R
+zv1467L6TBCh3hTkzi7o6EeHrHkT7k29mwDfRkebQJoFaGcl3ddGwCg4Ki9
4pkgiQt6iBtCmiCJ6LmHObHTZ6+2N0PauB+Ju++KJ3Zw90UI0TfqRX4LK/qk
XBNFsJYzK8BTdGF/3wiLq6a5N+IMsVi4v5uUHupwkyEwxzcfsAU0MeHeRTbE
MTYavKstMwJeQD8i2BNZnzfKarCHCIPbGKIWDLqPfdA0EshFubhHhRztNVSE
nPvBN8izoG1sOOZ8GiQ3VB+PWV33HKBEl5Uy1QG45IEENfs4d7b/f2BtOy35
BHnJuhlR0i4oe5SYlrfxsNpOnhgOhaWpyc2a9kbwcsvxg1oTgEvRbgrZeMZ+
cohJbpNzCT3Nac+ckRoo8hQBfB9Er+UpLiaV2hJx7bJKhsiGvrUyrw28T7Fv
jKpZBlzaWxSb9gugVcK5xXSHM8PutOxq/VUjk6EgvOuYgl2SGEZS7EvmI1Qw
9acasaukz6mQTSTLzo8o2mX+7XjHyFHZ2DtQnuWIh6jLZXbr7bGJ8XDFI4Jo
K4PJ7D8pJwcQ9AcwvtsjraqvaGKdNTdWh9fmqWBZBIIcP8T0Kyn9QIpboKhp
4JL8Od+/OQOwFcmD5l4MDnpImEw6dZZBQ2l89Knoyij3mRJsU/lRLRd/fHLh
JobXdwk0pWjR/pbXIpCTSRMJR2t2grQ2IQ/MhJr8J3pJAycF5B0fojOBgjio
uIepKMkciyhVwybtZygRTjHeKKi1YvRv5Yb8i7qf0AbrPzNr7pl/fp37lvuZ
FPU+sFR/btPgMEmkbfRAH0LYE+w6r/lm8hl/nPMw6S4xwRsSGikuDBLXI629
CNTkj8OaVfDMUT+36sHVzsniiQWvtiD0nBH0/V98YtMBHh5A5c7V5Dhe0ib/
8xaSbefT2EMn7SDUlLJA4/Ph5mHrcUJlng9wzIbwTGAhgfMR1+foU5ff0Q3c
r9WSJRqQrGSaQI0Z31llciSdfmx72hFtXCdRGEOgAs3MaFBjDJnrSXXjqvuX
gBAyFMrFtFlTFCWUrVwkc76xp5o1cFa4GVnVvdF3LEZ9WhQRVsZ4EBnGZ4Tr
7vRzvNXAWh8OgmkuCgnwT2KdIPL5pCNosc6GY4v8ILtuCnJIWh0YgAXsKzM9
bhyZW/9TGu3c7cATKUqYk06xOTzc0XHvHk2qiJ9ejyf1P8aXXzNtxN5vsYQw
jqb0G0l3Kn1QTh1dYpqVSCFGdYWwJ2FGBlGOGNSr1pm74XRGJK5KH1dLQURA
1y6GFVDn8AM7FjpOxwqsrP1bWyU3hDQ0djOdpY93betL+h/5hjT2t4qna+nn
COO4gXlgGmcF9xKTPwBc/5nU/bIqDtazTcLBcXHWoFFmd/Krw+llU7o+1S21
pd+Ab71ARYbDxYEw+uyQJU8TmPG9un+Hop4sS2e39jjMCVB6xHajAsSPO0jl
pZ11JQDd7SmpVN7C7PoPlKiS+BxT2P/LYlKevcR9IMiO4aumMrARA9Iyd1GN
tdQTvTSSRQ7Qkh7HvpyqCvF0mVCoBZ/XORD1Fe1DsGs3FQw3lQjT2FqXKPZa
CnoYkV1ZEZ/cxgjxscCxK5h+LdVqFmLevFAziJvmufiIfu0zINgWQ3sOvLVG
PYMbkci81fqzsALSscKtj/AKcsfBzDo3N4CDsgXf/dYxcevPtDz9O5EvAdch
N2qEfJlDAjQa+z8eGZM2ckqw7pQS5orm4bOWojFNAFzIyQLg89aINUV4XXNu
85c+0bSqDz1BxWdCjzm8fQTvmqnD1Ww8hsazQdTHhhiypigrN8YGvNmAUGEj
F9+MBL1y+WkLqGwQQfdlQWqhJu7kTjZIup7v/NXHKqsWJ/DUDv6DKECXY5Lh
VVkRMSCC6hoTI8J+AgCRkkChFN0pi4A8DOGnopJ0XPE40pW9y6Ll0iZBFPZG
WAZ2Pr5+sxVCp03f6frIaKdBsp+I4BqakFdz3abQL16d/3SXSup09AgsGHKY
0EdxkCF/P8Nup6/qZJxpd44yppiD+3nJtX2u8nvfs4bzAoYJb32Zlf8e+JzE
4KNQWtOV8yyBH/qjSMn2+uFQf3yKUNnfY5cRDGVI+vonX+Z/wLRjkavRMCBd
W15+q22UzXcE6Fj+z7GZ1/+0c1UxWEE2ZLiVHncG2oGtsnpMPCCQEgw8/Q2M
N+C0bmFA5kO4VG/HUEiSg91q0l76R6MRt274jZEs3PnVI0TSiAraJbaXz+WD
OWJfBG7CvBhBGuxMNZ4Fh1L+FpGKadi2wxtdL+3SQ/sbx6ZHQPpTb+p9oldO
bkkQMc5Mu0+Vuvh6MqW0UOhga64t1oOQenKZVpLPavGAPnsmLPTqQzlqr5Qz
MrgTRdnA9ZQdhjAGwk5YdBpwdcGrMm6m759QPO23fLUk+mdY4L8GSM7c/ozI
nexBsLpcNGIfSkjMy0C9C2dtVL653b3ifjqOAN3pZtmlnvgl7vknwjeYefn+
Wsxu7f1Shekty5Y7WAv5v0SEPCpczo8uWtlXUraGvZJm5a5hjb/MXLEhkwOi
tVVy0LiEauC8FZNnVImKvzdoqFzawpIbM1h2lSQyxO8hLi0lO1rEjbwQmL9Z
hkqZcfebpr+HdaCRAbS4H838SVyrMuhGuCN9EqBOnK6to/KaU75bpUE0KiAZ
1t32miZCDeoa/Yf1ixBr5/WxqQ33OPHJHYokYMqcoXvEARSnZ8CTQwPcYT/e
kKL/mtFDTepks/HmNPrYqEfpvh0DKdd5a38yff61u8F7Lp2wfTwGfMJLMK5Y
xqCVzlBFCAwe+JoxNzBnDSO2kUzIRx34NV2f60VVzBYqc454+6TB8sumVRKy
DDmwBWtxgwt2fiDzUTUD3h0OZOTSzP1c2JXd9D0mUzz0RQXdFbfNtDSiYSsa
KpjhUgcBCWQExNNcik/LAElGXiozO978L18+jlZ1lquwbnO60OupoFFf+2pP
CZAyEblmyD/GTnTjS6IHHa5MUWtvIBZVw1Gioc1ZEgaZH+sO1edgKQeF3Mnl
tHjn78GGHmFg7x8XqN2jMB4qGFX44mCORDjwCgfwts3UdDdsgQSWVO4Y/bzG
s0WeySe9coBpdLN6sRosW96VpRzNepB7kcJ3xBhmsUhcbPBt0igQvGrtqM7v
SBxa56WCyGoZftBcm7okJTRb14VoPlVoFkBb9D1wUFoaVjO5tp2EmlAjqjuf
Yxd3JANKy40NKylUOdykie9kgl7vNrxdaJg1rn55k6jlWdPuxN3y8+fyIx00
b4feL9DPPVnM/K1Z77RC8nN4PrYQHsKf+GUftIURYVDcPVx/gNqBDdDZ1yuo
5fJQ6NLbKojOqpmkNfI6b9ty51QYqbKClQt/ZASJSmPGcyyJ0gMPJUrjbFlf
+/pnFO9t/k4hO1242DxwZEOfY7MVKXUv8xDSzsM5aFlT7AaRdgexMm/6jc0g
EL70Z64Wyht+xPrjEEfiASCI+t4FaQGeOE8qTZKaDsIyAn+SMqn0KuXi7e85
zNkS/+0TzkXlZffD5dAOYuDFGEdZUGYIqqz+BoV4CzTS4GcXpejtFbtwNwIM
fIUFbRo22y0tvuCPZh1u/PB2dWsoZ1dVoMI6TvgdQUMtsuEZj6hxFO+wnACb
F1uQhqZ3HEXlnAOM1VgeZNsdwTj0idulSajfqNo3Y6PZcfAvYYInOFMoDeh2
zRg9YJwxmkVw45DxJwXHNrpNHI+b3QmlfxGCkmdGIC+Nx/iEsR7Oq1sCNyed
bK4+UhTJUkHHGfjs2ZaHE47ghR43WTO0DghSUNrHHSrMDq3gQvxjHbZ8TPpz
OR19usIvbPR2dIz1fH0UJyTsFPzQSB8omIgwQutglJ1hGMUmd77xVqLwgCC8
joQO+XExuos2lepXg6gni4P0ThI+Ekd4BvjUgiqKXo85P6MqE7C+WVc//DSA
QZsBOulXEbBbTu3ar6V3hNjKaKUZvn08yw5akzhgaegkSkqGxjfjTTGn973B
AmDvu/9HpEcp/bY5xQT+IvVw9fnzvWyFtNodxc6+/55nhgj2B7K4t4D1QFR+
q0mtu5+qUDlKDWo0lGgB2mW/39rPEYI6Nw4pexQDv50EOLY5HDaqMsiBnYSB
BiJv896tO2GQL+3kGdHBALTu5Yd/la0R7yPDb6YbBzLTHXoaVGOo8cL5iN9r
OahNSEgYombhsKj5haI/1c/xI8jhi+Sh8dTW966WxvLpSpAHJ6Clg108mT5Q
FihBWbDnpPdeTrfoZDEdNVVLvgk6ejAGqMBizAgr7H+aGWCn2kNC09InHr3H
W6dggcpd4iHXK21StvQPU5YM9VEAVf70BCCOMp5aCXD8mdP6BTV0vRC6yEzt
yYudRlcn+pczk7DBA0fBLkSeeb0/B2UZf9GqTsQ2K6ykfl7WjwmQ9q7hx+v9
sy7Sy18vAIs1gwa7F20G0ypwsAZOW552NOgWOHUNcIPO+g7NPCXgUgllj85m
5AdWXrBms64E7eIjgeNvGnMp9u5IqWGOv25RwTjUaR49N595qbPzgG0LMSRp
E0cUzMV2zQ2rmdP0hv+A6K2RRP+m5hdTqZOXGel12oM53EsQA6MPuLEhtHib
Ue1jSvwSOVjGy/6nCqlwzJkrFVRmO3PEFmKX/iCvy5lsHyFSuN8hBgWNbODw
09WRz8yK9Jm1VmSScrCdNfrC0WCBFHaXTpywZj35mtU2LN9p4b4DkPrPeEAH
ZKKBnyLl2WcgS+xS9S020x93oQmS8fJk2avArQtLimZXbLswkca6vf2IzC88
YAO73vWfQ3lJCJ4JDMzGQ7AJcCf1KFnAlyq6A/pnlc+GUSt5t/eQpAUIVnXn
DeZiXyutO/4p0FgrL18o1Sc+tIZ52GurajfXSpKyx0BPsgxLz9BtaAK4aMyk
es5NrT5psUo2V3PfY1vnxYbtXhfCreBBGPKhluCpXe5uZ8T/4iCI+OVk/VNM
3rK9VJIBbqDAUmgg3YqgasgVu9sOl8b+WPlcdFm30bbJGUVujdmmf0+79od8
MMMv/B8xcuwyFfpWRVnhkKOf5RWYpMz/ODw35/0qV2pMZS9bcOVrgbNwCYOj
xM/JW/62ikW2V/opuBYL6LZEsqmnD5fWkJyQd1r2q/D2lBBdDfjz4GIrZAXP
d3K/MVus5WLr4IBu/9qZYlxig9cePCBsjXP2m/omtqouqZxnBsfzkyAXA47n
snqlGUgIP5XpvNISDFAGg6G3aRH0TtgZ0UYy0vRZnT7/j18Ra7BlvIHmem9A
dNezzAEX6snki9lXbflfwIX+vejjagZVVUobNAgTWf8Yp0msm+0tpeKWsRzc
tynm+5jhYqj/xmlzqyAm0PCrLJnsbVJ7kccu9yDLE0a++UqcQcNTxZJY6Ym0
ijgyyTsEvhowNZVbG9L9fvM0bZ/durrJ7cCikdjcx7O4pfYt0Cxn8T8lY7FO
hta86sZas5YRdGj8k74MHQ7SpaawNoamqwAGu/5fqW5MWLX1jie6vwau8imh
ZuzKlEKYLMY0GjyCKJtGbKCeOk59+9I7aaDLsSJiMOGb2HKeyperEYLSsH8B
V4Oe3HD2nninfraRcNOyIxQU4TPZiMMOEkH6/rWnnlbot1GggiH8E8MuBJq+
/UuOOOvfLLFPsjc26/00EpDMPfjb6fQ1eEgjfwOSbPpgF1PwnapbfYhlW7Az
do7TCofxO60BRaq/xcUld9gAVYNrh8HcrPP7tcZk0DtOv1PPc33VXvQ1QDEA
2QT7hC+QGM6n51g3hGyZTwJmo6z/0HQ3UM4IKkCobjF51pYXHzOyTdWDBZBK
aa1g40jr4RpD35cpKriLiJ2xa2NkCz8+fp9yeTDeLgPgQ0VX7W2bbQS/Ste/
KNcU2AjHfahgBvBc2OROc6TArDweSD5CQF5dL9Zle6DRhQf6yKMP+/hlX19f
0BgixBF2TbHe94GQ2xyAAq2xXWwLZOvjmDnFo0+MImmTsyPaUseFIaZtBT87
gfgtq1I0hhJv1IJHE4f6yLyed1DpAsvMdJnb3zjWsjmBqorZK6LR+vvYXWfl
3PBnG3e68CFCIhKpIxqVe8ll7+r1oNpmVPO62W9L5sGxwGl0JICfwCABi6CA
ByHGt1xZ5f19RVMnGmwl8gqW9qFMf0by+0yk0h/eqHVn5QYaURmm84aW94AP
w+u7uBZIbXyDE6Magztt41Vv2lHdVQu5N93bR12kgJ05LGVyH/c9zuHDu1w1
ohVpme16dSx4Zh/4TyZUN3J3+zKNg+dlOcZ7vT6o7TbAFnnh39r2byzcf4lx
NzmCd7L0nDfybNqpkr5PBHCXaYdcpS3YNi11V5pB7yQRIes1utJymmjPyygJ
aVigTbYj0yiw4f5P4C5mXEYuIcypGmTpJyU9GXGhDXpmREjk/tRKOBXds4Tk
MNJQvxicqYJ3MHb452DFn2cILdYmz0JUU2bxPaE73v067QJgfvlDypq76950
68DISqDxzPqC8+imYa1qHqPPjs/0/5YExGECqt0bHV/eVtibmTlc7R/noQOX
j5g2ByrYyVgJpQvRFir8FOqV9SYTErzDAQwel9VrLFDfRlp5CTg8UwRHIS/I
3nnzCgxksbhYkwZOhQIEvo7urCvdxn4J2I1tlL2Z1hDZkj8S3uGzyD2hebcQ
HGhA6nxb1jPicnipLusRZcmQOXqQvGFOKg7dAIPRPnapU6orhPZjk4tgLrVb
BKvx/nSd9UPagJ4z8fjarj4wZIkCt9AcGbUiQj9T5xAxdvSZHDyrzfnoOm9a
ZL1M5O4BluDDcXamostlWl22xoU03m6xNws1UqEGZTMz0VgKLNHsfXS6zovy
RGSF4Byag/KjkOEDzVnNvQkkCBM+/dsCdxal1ZtzsTGMqIzKAi8HOes/fth3
vRVLpBZ2J2xYutvGInPHFJurlvvPRi60XCQyLaEDAsYpIAj/aUqxblXaaXso
tnFqyKnvGhh4ElQmdtQmk3CcPiN9WJoZOAJQOvHCyZTQJYQU28mxvGqZCUDv
jR86380EpaQwTTlCn+EVDs1hgvDdm8tpFOIba0nSqLaojImXvLWYG7DcshDg
o2p7HSSYxvG0XMihbubcjhXIOoSCrWZWqpIJMUFe771ou7Fe1gdvpyWtTfkL
EaD4tBT3LREafi61pLqRPtZEF1f7IVxEbcFVDgdX+RhHHk8NjH2YCB4CXB8I
uTPp3avutCfsxnFPkqogp+28rMRslM2szZBE9aFJXXPDVRLNGQE6tJK+J0P9
Jx8mkj5YuG6QeQLBWU2fkCrOrjiswKQPlYtlS4+DaOpsfALwFkpPhKh7ysML
qa3OmWxT/eJWxxrKcfdd4TfHUo+nURhfSGPKMFSlPIIRL+/QGqZGO1Iwttvw
AjX3gYS85eAKd0hgSeGjrzNqg8Dxn7zmSq4B6VX445dt8xSIoCejcFFiC5Fm
GWeIwiUdLv7yn4FsPj/LdzzuodM4E9ZLVeSZZyC8loLEbYoqXLop+nAdZSX1
OkyxClnYYugrDTlHrO8NZ1YJbAvrVWmEYv8i7pw9jG6LL7rbgWNMMUCZdKOK
RP9U+vV0S6tbXp6BvRvZOtcsiOHifV9KTPVKVSYYD3igc8WvLyMiSO2QkycI
OFyNdz+PXlPK4a/yEguYnGbFm6IUtZjXh/1WoNNfhn0IDiChhMQ9Lupw/qC0
DJwrGrAC3HZDuTcuLKjHULeU8wlwdY66Rfl6Wy6sDHqWbxy18aQYIb+8J5wI
GYFgxk6PkD370UIDv//uN451Rvv83Be02S+qKMA7Ckhyu/mWiAT7xDfiUU+i
/zZZV08ATDpmxXOCRyGNuId1lxG0FVeUzf46ty6KI70zUwbuEerFsQ7X2FRL
8MoW/mYnl0o6PDbx6JNk0R1RpUR251lnllR+xzm+ByhZHlPtCIQGOtEmhMcl
4q7q1bhDRnjNjZS0NNsT/nD4tRIJZc8JvmfT8XYXJHmWqgSu/IrOWCNbNbvw
3AS3oQe57UjKoP8VEcPWlGQAzRRAbrX9dxtwHfIhidDOufk3TwslLg2jygQL
R+LaPSw3ZrqWc3D7nlxoKbsDFyXRNhQCj5Z5UdHDT6oxBr28BpZ7OKoASTil
V1n/VpRRdQZjqGO2atGxKIvh+GxlpEPpII/5jz+gbfDOK2SJHLFPNOtnXlw8
cLW+sWfV/F6MrdUv//yxCQMDV/V0UFqf2+8TlOZ91/R2bEDN5SyCAc3b25m0
AkaxW18D7zF+5uNt4+mUM8VTZkDH/90xfc8dHtJaVnvj+4SzTcTYevjHvL3Y
g+o8UCqSFkU53sRJKX+9VL8LPAEaiGdqcosEjKERROocYycmNJnj3crn892k
px+/OYE+4O9LqjP9mXG2vfR9bP6iEpGSTCN2AItbjz6ZmBEp7SaIfzSH0zEL
DIVwY9GztzU5yngPCEglORuPypQia3XA1bFjsXvBHgsW6ZAnf8XK2Ble5qOf
JJFY3SyVEGvD63/doGosvhSqOR0nFtv1r9ydG90DmUhQdpB3JmGgQE1wZzli
+Zakyqq/IKb/D0aewkeFowDPTL/7CPb7RZ9PxnPWrLOThHNt1Y+fWh5SEPyP
RHvBRtfJXDdRsytskcx+DuF/O/9z7N93sULhVGeoBvGNHNTqdB4DLo6/qvjv
v4fwnBVB5dz1sEbdcd/K/CfDOpFEvUyDmp4rq7gtrjY+GQxKxBHbh+xni0Li
4hr9rzQKKH9aWYep9RKKhZwC4Afo/C8Qjx2atOhszLb7Yl3nySlT75W8ijB+
j5sXbZqJnKbIPM+dfe/imuSJCWzhi+/IOYAaFCxoIlbGVuD7miEwO6121XMU
ocWN7PHhMBLenAiom2/bDMRUzgVthVqhLj5jlXX3eidoV7o7NW8CqA6jUTII
16zNsMv+v7nRFhQnEiWDVuDE94xWofgFWKTQMTF4GnqaMi/iKQ78wco05Gfx
zxc2I4UxJbphwnc+y5Qa1AWUHuCWA4UULfaeVUaTBwIuLcjTw9TphALOQ9gp
mTvy8fPVdzpJxOAGPUlgr4x+ILvqSG2p5jgwYouZ/8leubOgERaLuhlsD3z1
ZlRskMWoL/Ho4zGWd64Dda0qcrYGfAiQyN401gU7vtzTxLYVOK57JL3d6BGd
thBRV4drMmEanj0bMemn7Yu0ld+Q/ovS6Gd5D98I0u/nJXVq5hNZadTHgIHb
yn1pbDxtaq6A7PNyomVp3BXbjTJ2fmqSNShaSPleY24fixIRSZ0DhIIGqPWb
Kp3AwqNcJHFjG/K5kgn5IOVG5hTrLMmnyNO7Dj9RLGLiQQYXYMi+d1y1jFB9
nijLMm0R1HdPDVB5C7ZJIZyHDNs+/MwARjvzuzvweWqO8+Apq2og2lgQKEJE
PY3NYjFvDJYZksz0BaG8riSTXRAS98/QE2yhE3HDYzhSfJC3aJz5rpUv9JcQ
ZwT4/rU/R4jcle8S4laFKXpzJkblPYGN/wVtNS8BO9BgWrmbaK2+RzhaP2m5
m3lJzc08F/yb6aX4YCzQh/Cj62VCNqF0S+BkpziJssN5WyJl9strZiklltam
APSGN64wbNVatcv/19vky5Jk9tr/baXyh0EmMmS9dQRCDlRBByB468CAdXAo
zDRbTGN1yMI51QIV3T3WSKayXqo4jdzasvyRmwuKaT76TXMicnGeVFInHvmL
r50OsHTSmpVLe04snVsrQ6stLlRLrczVXmA2y0rQpiHtUsXtKQuSdBfh9g2w
cTT+lA6vJGsx1QgUgLVvuqcRr46Jp8APnQRl/NQcV34eNAxLcE8yFZbnJARb
szIfyoJIyjYQX3Ok4CEqzQzVJxO/Qes8aE1I3YXDZ/1bZdy6fdU388uoqvJj
RuttiAY8GGNYl0oHk8CpO7fHoxjJWQbKdVz0TKSJb1VcsozvBG8XIXNUQBG6
a3Dw+rryWmU0xYoSFWG3zMgFOzt6VAoKI7IgsDu2RpjQDvZQM5jR/84zapKL
Dfy3nAHC1aS450Vii3HrcT4PwwRxHc4fDSbE4o/sSgzZ90m9qp12Igcs0ln5
S8XcgB0E9e1PbTCZpxZ0xV0g5GEzUJA+eTWVvbpR6CmR3PwyJV+qEMqNuFZo
7t/B+hkBrGmXg/qv2Ti9qxjCyRMrTmOZLJzfnxGQmufDPpg8bnBeLiqwyJry
daIhCuqeebNJA1V20joZOMxTlOpDR9blefk0cX2DPlnnvJLYLzXXD60NfpHg
fORGaSA39HwgYNtl3jvCXQilac4W1oQto9MWOfyOw5e0TPKqCevMLIl4gm86
VhIfztWp3KDvEnFq1B3sfdIWrxCIPijkx8TnMQqnKEFGmV3CiUXVkXAnI87m
mikB8of4KspEiySELjMB/kEdhkm5tPaonEzgSwRwxTuRsowXITEiqHKCaKry
BkyBtROiJOOu7qsb57Tr2TtI26VmM9vQMhnYRU9DrpG9XfAAwSlhpwMK5/5z
yaswo8rLb/Xz6+nj9BeWv8oDnuqCR98Rj/lqWu9ubLIC9w2JwAYjdUGP7vXZ
0dYUq1UV88AMfFRouH+wTIVN6q7IKiRQrOmZvKzHpHCvB4NJEraZtruFlaS7
yWt9HkqzKaatIrnj9FjrPsKirLSstPJsNZb4WRDUrnKm1BbZG01PYvFC/RyA
r0Y4zfczkiuIgeTjc+HA5lVCjlzcXmeDR7eZYxYj5KQuw/tgcVa+4fZiWHxk
UssttSC2c2XMXGqbGi8z5nKtZtBdyuWleK3i8c0Vy8XvfTarGbloO2fx9Qr/
QKzzCKs+G+TOWHrvOAJJr/c+6uibCUXOh9sotq/+fl1vRzBQWBkDC/ZZvMZK
EG7Ah142nyOjlEYTo0K9JcPYHw8PvA7QfvqmYGQKB3OTXbu1OSo0ViMo+a7D
mERrDtmPHDt9NYgqk/NbMeZtceV79LF5jHoYxsrzNAYddt5bvmcpximSN8Mp
KUIYdkor+eF29zKRoMftat+EW2FBI0LFescJvXPZTh3cR/iPlKyneGzKENA6
1t82i0o4nK9yoP9HOygJqfZ2Pvf+LTmz+Hhs4U3W+g3kVuZZA6hg1/SzN+JZ
MKRrpnuMiCnbBT2UpjpPif8mYqGiK70p60D5ae7/UoZib/X5AXjfpbqe9Rxa
peiByCIIoTVxKMUUD/3F5pWXKqlGPf6+y+RqlHivkBpWvxIensX6FY9AXTiZ
N6n5QadM3N2e+U0CqmXV2AaoI5mYv+vRQH9celZqZpvEmsSsbpKt5i7f+4tE
ffH0fY2i8jRaXJ7G107wEiMuRQMCv81FPxnNmqHzvvgcY+zbjrFCSCt1TdJA
5BNjUdYkHvmgbyEfSsBHz9danR2oKJcjVTZ79McOlBdx9iLFOCOC3V2wiLYO
pp6DZKFjn7I7VVt/sBbXVmj2zXdTshI+Nmnf6QxAPA2FYSXygdD2pWha9QUr
NP5FmpToCUAT+u3ifRh/t89GYnGYb3XiW+0L3bQ+l6VBLb9SeK6KYGQGas27
7iKQDtMqEm9xzbwRNS/0pU5Ezg+pcTc4A1vsZlHiVvLT9e04lDkvLS/RnRLF
3OE5P36Q4QjtX0bY4bY57xFaOtk6YiIye0TsH1BDOsDzal1b4x5kgH8CMMol
knSU77Px7djuEdGGWjw+dGCM/Vj5DK6GKqJZ83lepBQxKG9mGWeGZp4DDrgS
oC1gCpUXY89Zx/ieKNF5sgIWyYCvF3ZWkrVi1pkGqCnMm5iR5gsMihLs3MDd
FRwmWnyYrsfbcsSqsoXQKeYDgDoglZvuDM7AZmy5qjn2AWDbIPDwz/CDUnOy
38oL/O/kpnGTgavMnZqUvUTH6309E38qkXJMVGTanMuwVQ+iwQMnYgmmq3+0
I0J89m5pZKioe7esRmV0MP6Fsstq505SYivsrF8VKRUORmW7JV9W58LgSc8i
gKa8dLn7iwKy5kmgiTuWJFqlcTVOkr5dMlcbS0DBkLU/Yf6F4ONY2c5zYtVc
wSWRsTrg4kQG4IqJUjTBRxqU82JTUVfUdJrh23oqZSolsoVsm3ObX52Q0ZFt
ai0TKKe7UTFd9omiu8frl+4rYsi2JPDc+lbWB4aax6WYmoRH8+I0n2+Ie8/5
qNKJhgbjrWUQ5+chKAq/u8w8Xg+QpvCy4FLwjTtWrCznm5GZsS3CjLlvfUT/
pknzzlBhHI9UqW11zrFMn+8E2PkNIZfZmDzPrWF32+WqgRa0KxSaKkURPCLv
jpMIg7mh/fMFUzTlwNtOZTwO0RaVGyQNViwx8m5GdLpl+VPvKjZsP+8qUHOo
GdZX9lesuRvsjPMRTMc+ri0WRp60nSGT4xyftTafZCd4iIGaqVc4ijyfu/RY
thyrOG2U53SzBXpQIV3Aukgi5Hm83wFoVbInpnM0T/pXJaSjbglk59HXK44x
ioU/9Fhw/JUrPwJR0zmVW4Z34XCGhNb6Cnv2HQoZjH2XvOQE1u78Bm88drwO
KEesflRrvLmtgVcJYqLvv+Po4o+QyMJHxOcC0nff6XxT2rc6CX5vizn/7HVI
oi7yz/GlAAqsDsE0jHfUaQpdrMM2ofqFbe6GNEQ43zKuiQooSzoTknhXfWzs
EBzPhcw3mccFoi4ajmH0gRCNsfdzBo2kW0+ZK9A1DMBsKY3osH4f183uYwgN
tBuXKfLW+iYZTkAqcX/pp7CSWAkP5N/o8PRQzJvEW7SiHmR95EJP2ahzE5ZV
ZK4ziwBly3byT2cG2Mvo5y6jIAnZSogDxJ4K3AQl42Cw2sJGOiHVcSjg9uRR
0iaNlHPOHUyYEV+np5a5PG0r2TNcEYdd2nTw4GOw5fDKMVly80KDJZ2wVeg1
3jOsYsW0cagq7t0kgHFurklNaegDohRhFDar/3ObtbEChKOPXApqKEBvMKO2
tEM3pq+cYi32Ett2PwaWU1P7W6Chsa6umvy0M5ANfI+xKwgLkkBYffVGq2VZ
nCiQTpmyxnGhLhITKvqDpI1bn2byIOnic38/OS/DXwuj+xzXO5OhI92ItL8S
5Ah0UqWUmHKqlKlHlzkFbvtPvZFnbQKJZNjp2KjoBg3mXp4DozH4cPIN0Wnl
mZN1w5hzYL0K7sohxmFG53oP9cF30GgihEXmD/Axee5rKc38i2FpSaImBE1Z
gGC50VFo4iolC2rBe+wWaQoEzsUkqQ/RMqnAki0YxYHGrgWlKo0AeYt/vcFD
J4iuEoVrQeR2uQuuOaifWiACQJ4XmGvltRnn6djaQgGuSVag+aDV442wmPTx
u0ViluoBRWOkI4RI1LM0O1YYlvb9ohvWeZF5jZ4SUD7tOAMANSqae7zL1G0q
eeYemwtZmUWlTeXpgR59fiwLLtkX88HFrSf9v78l85JPksF6CmewQG/q70Bx
pyspqreATMZCxYB5+dVFCIYTFBDlHRasK7fL3uX0gDa8zqt2CTbmd0+149+l
zrWYWN2WBq505x4yoXQGWWFyqiLZ1GF9ZLND8HeQCH+wuexvFfEliWF/LrSM
HHeGIXx3SgG/n1FoN6++hGH8uTx9ZWS51tN23QPXJhWFLF2vW8xy5YMT/wT3
zy/6gVHLdEuNavY7u+5lM9WVkgzxsdZWkIONZEypaJ39+0XmMOMDshOk98SG
VYmpjFj0K0mKUP8xmqnhWTrMKqOVakFs7mF0U8aPUThDr4Bsxa9t0TpaUf3B
77euPqaTjymnIgcLzN6FGBHg7bkqrCnj1C8/kobDz2hFHcTJ9FdScg/JzqOS
8RyhJNQtae4u2aDoT0lgftQD0X20Q6p4osSPiDj1UDL0+0VuCrQ+NIkv6hur
9YhqKprFu0yTk6d+h/fMbcjjuLCYSxV2YRhVo5XgTUnKXgqDks69TpwXo7D2
NtmOt0c2k+cd+vfAYT2Kp3JJ7OZzYVN+pyvUhFxucs/S/pqVeZwq/NU9AaqM
wubQb17wtoW4qPXKR+YFWjl0cmjD27rSCsL1sx5DwU//rI56iq3/t9UD/OTy
zTe7DaqRb3gSBUQH2R8VmPTJjeTBjsbtZ17VnhP5wKcjTb72gW+ajd2NoA/W
M2CWYVqaO5dhWguf8bp0NCU2/DehZvYG9pdGJoXx42TotHzIKGSWJgbPzBzI
cVtEwkBqIjVjPXs+iBYpVu68RE+oe2LObctTEQgOYcgkyn489VDvqxABlPEH
32YknhdelYQw6xYFlc3EWeS5rhTiQbjfjkzcdpQQRRlQOLppCKRnyDDuJr/9
pqMzxRFaJFXvV8RqvW740iihWJncjZnyayLCVugqzqU7aoDodQKxc/r5AM6x
DhJqj3HKm/wtEKvfUN7AsEOL4XdQq3pJpYcp0jw3BLRVQf7S3gBp5g9Bfvxz
cFKYDZkNXK8Hd7UFs01X5pjUUvRsIpuRJ/br2EQ8xXPbs/hTYc7wqK73NBOo
v4wBTwyrhkO5hQ8VblkyPDJ1x83El8KgLOyK47qv32MAOsRuvjKJDYgHZ70D
+SAVF2qxpsOmEFe8ZdBfA5fHjBf6TZPiPGHtyRbdnLMGgVK4w8eCrSiTBbYY
hR0Hu6pNCSx4arF6AcKmrMJ5rp9mLDkk8vp8sjrVqNfwyJAxg0hdTa8U97YB
mUCgQZRCPubEZKNs9hTM4cm64WS65/vF3CL6djhP1QRJR1DuYebWo9o/cYnN
0fqsBqXZozlsyb35TMHhbgkB96arlB//Ez5npoGFuG9fhoaWv8VMcItLWTiv
JNRrjy8xx9/ynFm4eQaq1YeqdRy17F+S+bxQWtwBPqeS6BUbFJzZv08HJpkM
P/edLCrmbSawOKVykL/M2xEt6Uc5kHNg6xCGZ3dooCZf9FMhiTCAdb/57FRY
Y5W4Bwu63wlnxNR1ZiRBeYrIAey31Gw++ZoxCFeJ7AEtEJospZGZ5kD5BaKx
t3rnO55wrZzo49HMZrhy1GOhgpHID/7zwaftT8MA3w10xjfzfvkDeg91mDZP
Arfu010hvv73VY67AUH6tsEzmK+zDYyBhNFelWG9uJ/X2BINX3eDh7sIPIa/
DYrpUdLaYpV2XuLJNAjkMy+LZNRkPxMpYEXo0Tt+60ueHOPQGkF9MDaDY5ga
8MYCDdvE1gqSjCOwIykwz7eucxKUuV6BZYfidtZkgcmQCc9SDt42jRU+kfUq
9KBWec1rNh/urue7g0XzTHk0qiece2nxsWKxqlM2l5NssKnu94WoIvii/DfL
YW0IhXkNbkROH+NZxuVZw8+lbSW0q+Zk6hF99xzeT8isbkKehBhDKMKI6Ch4
ezF884TFPiX6v7bv1hXGI4NX9+lZz2PXUOBxWdzvmOGQFx0XqLwFR10q/oGY
AKSbirwMe6AVpkkma92qJr/t2CHuA68nxiIE1XUHebrcIIo0yUYD3wzI5DBp
WcCuzMByC90wwt3RzGg7kPo45ArOupmahXIuNLwQ2aMFkOgaxr5azxHvyN6L
f6KiXcrJruYTCjjL/3eyCr8j8xPQV5QUOWCKIVEKEo9DL6H5cKzb+Sl8jJ0N
KrDocTSfZ4iWM/WYFhXqMZu1hslBW6bB+6cVB5wHjYizNaaOUjCsiJZKI6to
E+ZIN0t4qupD4Mg7yHfvXZj90XtIGoKt+0+WMtjuKlCkr81var3YM0dBpgG4
zFjozBPLBtSKj2FWvCOsT43LmO0T5ntMbXZiw8ZNBoCGYSDn2fcF01f/bdC/
Lq5PIsBon+RmIHhBIKSb6f1GkIqMtSh4xgk9Q6lTWJZdA0XsOYdR6noxXVVR
/AaM78GDyy8G/rMnncgOxXev02+lCKX4sEej8kmaK+OIRKBSZe3fv5kDyuex
YZfEhZoJb3gQL6vp9P/0VDG5VDk4WZfFehQ0NQ5tUBTLL0BmKLg4ZZXAxCC+
8+uU6TQaoyAYhiB6KW/eWdS88RGQKuiwhtWWJmLOin2Cd8jjeVS44GdSxGPP
jOvysa8CNViyud6t01cCuzuwnJ8aEqKFbauZPGoQvuYKB9LI8lNpDqSAP7FR
kHSTo6QvKFsXfVKe6AmR5yXKYq0HWDvXveeLYVrHbH2Sdis61HSyNgXFQZ4Y
nNgr9Nw+PKpR7hccslqXxAZ6ZY7tICErnFyMkZdwj+p3vLPqTHoVtTO+Pgde
GQ0qxIFx2d8mTzPWyyS2caE+Vz9Nx956cphHgSPnv512ST+ofn4q3jJ7kIqs
zzD3hSMJYs57Y9g4unOU3CLyq+VmbPZx+vyK08RWtSs+AskTdX1ne7+TADro
39RtCia0wFZWU8O335Kxyt3j1wQBfP1aj7Oa1gKdp04sPMXDISSMtDnrqtHT
1QRsvZqKppxGW+itMHMkTS3kFMJhBIm5JXEN4qwz9lPeJgEzhMKc2qBE+p8p
LEsbTCVihxcE/KbrDK5RtBtJcXmhpuEV2TOelmNc52cgL7ZAYC0md4P0HrU4
sycVtw3L0ggyhM/hemp9yEnbMqJeXiwezvWEfYLOeYxNJmT30Z1YBIB1+WEj
PROcTZVuTV2Ssx0SW/Bb9i6aiMl1XE2FKleEN8mNlhfZgnDWlHgyMKD7rQ2Y
DUR7bdD2SiHL/JsDFYkJs+EK1g7F0IwC9UxwjuHFZ0aZEHivVlrwpVQiQX4z
utBTr6a3CoHtGsaOI/YvwalEHupLRX/CMfXZ4/wR6wMnmnmQEsly83HTxVAm
mH7q1ndt10hU8hN68b7chUFoPRSWuEJ+kYZgqAO1NATf24IpOwtHhMS32MOQ
UeKRVA0dRWw10AluLq/nEcnsAeOv9E07dsYvq8rkqV8vazSHsX21ANXv6THL
Lr2UeCFiVIiPmVvBTETK1fyqXhsYaIzzpNpOUqwpxkqCU58jAae4oSkFs9Rp
HVVz1H1EhoE7irLq4x7Yb+YdgCsGz1asfLcSeb9pPEjoxYShY4cnBIoi7pa4
5k9akZLRoJE4JCj8IxwMugn+yKFvRNZtp/PNkqlAJlX13PNL3R1JZ5UL+Q3Z
0BK/DDPi3iE8mD1sNTWKsgNvoieYhBWiVV+7EAM7Z3liL1peJQcPxN3lyO8W
EQMztYVGvfVArTf0rrXOdJMxsgSYioDZyCiwumAc1atbldBW3ty93GbyRq9k
hhYPwThbBFzJWfiMiYoTBwWb1+1oB59UuCmaZhSXLfWM4Tw4zeCwSPWildDn
5LcUD1HyZm5foSB+DxEJOjqBOvI27XQa/PYTR/6VN791ognKa9A9gTA6LO2G
PEqTzfwdL9iC29+DLNm8mKhitMJj+eEjdMC7/eogVSQ33uVxrHpbUz1W2BZ6
5SUv1ULm5rhdYoCZ4rIn6BdXKkCoBctWSZ7vEU2EAwYeJaz532tkUzW+MuXm
KosnbKXwPOG+4ThRovZnVsAA0YRr03OxuEydvlgSmqQl/8r80znSSWBqCzEe
xrAbBfiLlL1Mybd+wGCXeVXRSvIbK/g7hXu166K1mX6M9Qv8RmVEqlidiLdi
jpGudpEvC05LfyJg/FIaLsoKGyPY7gW1Q5PyUGQtrgRYgGzoCSCaYfn7n21a
sIB1IxYUXUasiB+aOfaDKSPNW706/bgvTR0KqPcqLCwO7R8Soi2+jsGMneGZ
ZEO4Xn2GN+uLPjFZs/0DUzVEqlpl+0iEAZR7HU5+GH+jL/LJXwN2QcJ0VQ1N
D6q0G/qN0sZG3i8RFb+vad/8u+inWkGaU6zxdGDZvZcthKxq7yBpf4E3Getf
o9R2ftgHKlIabPB9F8TntRUnbkaBp+paYRWEXoOj1FYNqegj4Ilced147W9D
vlLb9t6OJ8D2U4eUjMxxcJxQRfiVFDJ8sbZMW7u37MxzAhfFnI9afy3FJa7j
1MNOLPEgo89zm76UIAP+Al8xOp46Jn0mIMK0vH0DGsTWQEIPm1YgEg7F4iov
1iUHY+ceYwyoK0w4JxwULfi7Hojl/d9eam4Z21yhmUEm3oISVzBi/nm7cJiK
V1Rz+2uRy1VeZZFCDz75MibwCe8Kp7ZIdj0GHXbwMPZtGyQZTqVDuwQaCVRk
6ij/HPokE/nPuDg3yOtXGcegDxllbiipYscmBXN2/z+ht/mgBtiX/oGkihOI
6DGhbPTRTpLmdwAPwsau7Cmu3wg9MWdSeZmt1pvWCmfb0w2LU7e3P3wvOaqS
5Inhl/g3jjpkGQNBbX0XYBmSRuYMeaWMboZMJHbwAhNEhizzAGfuHqsowq0f
NOyaQrdtSwjKfp0Y1GiPSZ96hEV8+0W3EFROJJo6KDsgzOwTJGI89YfJql/E
HjMVBrhsKhOJsJdTfpIUREZv9TUSGS8ZDvbYbCjs45lcUpEJZlEsZk3tUKrn
eTMvs22+HhU/F/98ElDGwb3IRr3gTwfj4UPy+daXsFxIO8oe4+qEHs41gAPZ
8v2JBh5y3TzhYaeKs1jgashXMirkm3rXorC/W0WwR6648fIFqjogWxjMn+oQ
+QuYFe585+F7hCw690niM/wgFZ7a00Y0yKIkdMr94XhSvnWihkR1gg5P6QN3
pE1y2ZBkIPMc2u2mS/Lf+mQU+2D3bHnuiGoVLGADoiBckifk/LLx2WTovAA8
cX4gARKLUbF412oFUNNY2sQUoeXHmDP3pwbZKhSZN9IkVBf8icavfwNgtZzf
KfO+elxo58NtIvE3EDlNZ4EQsGyA9UMIiWDTWX4DHZAXlmdd+t+BXJzeeCBR
wIUfoq8fF0PLbb3/yRxGb8jVKMs05Hna+Ptd2MBoQKVx/o5Usag/hfUFIz3d
G6Ymucz4EddUsc14PDz7Vlh8W50CTL1MK1Td8iiFt+h98zI8g28JO4jdpv5H
4C6oQLZTXott1zR1QhUTVEXUugTevdbIczgc9PlO4ygST79/bno7JvTWTYei
29VW/6EwOfwnRWWyvgGWkFCxdQGRNrTi/4bsSfsKT+mg/pYLl2TJ5zCwVKn2
a4RMYFsyizVPZtCpfOooFmRzQVRz2IjvteLIjz623XzMV62iY74yRLg14sVo
JReWdSp8eqplHLDyHOfG7oH2fOoSxeDFDzo1V1NU9q5RgEqOloRc9ChBczJa
BJ1OfEar/Z1c7yO8ZaxeYlUPZo7GHZNdCz4jn0X52SnqfqEl1/s8OzW7CAmg
EqxECS6WOuC6w3Q6zpipihmssWUsqGxt6WeOAZ8CtgR70A3N5Ga6pywlOO0V
epzLYNuNMpsf0YmgMvbVskOgMnPO70vQRbtLYE8+a7OevTci7pg/ZZBnphAw
Z5xJrAW1tuzJ8rKmPA2lGuqPeQ1+F8/WMEMD8yNtJHmS7GMqyXwiCSPHpuwt
/I+5j9ftOVQObxZq0LqzPp18bJcEH7iAIzm3wk3WR2oqsbmfPzJAjNLfiDz2
YabKEzkxZQKntVjx4YAAvU08VOdbfajXpnXtO+UTJqa+5tBv7WDiArsE+ZsS
Wpd2VmgbWIYRke/OgK7dtIBtl5nhrc+0xF4Is2QO7GXQsk30hQ+F6EDx5aJs
fD8auRpCRm36ZLz6NrkI4314D0hr1cD/lMXbLkF7CAc8BnWBmTxix/KUt5Ey
PBkl52yTQ0S9fTqF5o2b7u5NmXvIqy6I41rT9hEByg4cacuVvFOzapkfbZR5
Ou5LFFsh0CvwjTTlksVEnZ2VntEGwZ5c17NbvpxflazlVNn7etKO0jP5aa3b
w71sV7cllvYWpuW4jP4gJHiZaP1Hq9FDO1UKzvudCH5hjNFYkKYnk4pr/kdE
JGOwx5RgXiwQ1A79hjJ3LFpjeZukAxqfEPFFMHXQMcujZ3Fj7GTRG5fUKvBO
5NeaqQHcJk7wGjd3RHjOa6STDvQldQQvCnZomDbkGn/SBkFGQaKxwBWr17wt
QkFL8NxUNRLUF6JoW3VV0bpugV0jAtaaUybL65X9djSE0S2cNNTTOgBjtudm
ApLDmCc6qVVTavAVVZj7DOK5T4USZDjxThsDC2CEyhW50wkJIZ8y3ZkxYGKM
UQqfHsUFF9zF8e4ot3K72p0DQUkGFZgkbQfMEZfH1Dag0WJc7HryCf0QY6vk
5TyO/QJSTQ9QyylaatpvROM3uXBpYgAI97kSQHyBM4ihMC/6CAanjO1LdV8M
UvpNt050fpyKNYEex/PwuS++8ZyzoqaLCpzOWk1S+H6wwlrqQ3ktz8zCPWKU
MLyudMEqK1FQINisOlk+t9Y9vxxlo+0fnPjyA0YSGebWo3sBB7ScfT7vXZgm
1b+niwSqRuJKa7fCBxtwhJPd1o1JPLEcYiCN3s4vu5xg3tuUxPwK4VR55XHj
et8p8DHxxnafBfBBYMgZqC9sz56cDXTfyc2KuZ72v3QuqUtYpEZjYyDy/BVP
gPP6gn+qhuoadyzUu32ilKpXFdhxzmYqCyd7tkN5p/LZSRSosKZR4sAEf7d1
f6MMd7g1L3ooeLGMwCew0jRIxfqlerUsyhidUUuxenH7DVLpllt/IoVIBSQR
GA8fCqSKUDxoFTq3XCCv4UFx+tSJDWYdSR1Xf6I5vx9tuYUcvzahJO11AckE
6n5OG2qh/VdqunhDubEdRVxpvwqgYzpQmWqIAS83kQn0rWSQc94HJQCB3jd1
fF55qRhMRMpVYkKYyn9UNi2s/yE3nWOUh/0i3KIwR5wyGqyDx4UqIFq+dv2M
mnYmYDG6LkM1lv54Q+zKoHzmNcLV95XPtI42tvL+FKpZKwPh8BE6OB/TX6Xi
NOjbAUgNVZ1wtRL+3jUaaOPGkHFuocHw00tGNCF8124JMjYCKdbetdYcSPll
c0ru4olupw5AerlkxAKt3gKUqsqTwGcs7eFdCIvDEh7sZiSCoP3zPcXhbvkF
ID8wV8mgU3nUySsQ/AUedTtxdz0rYdwJt1r98Eyy/ou5ZOZyctT3fmylJGDd
eUHuYrlq7rqHx942fGSt69r6Cd30s6EQfbLCh7MNBpXBJtXqV3w36fEVxVr1
gU3TO0zN/73LYFY86o3klfq23857fY1Oq6a+EipfVlEmhVNuhteCaVnPZylN
OuWEAm/HtklKijD+ydNbgtVW/h5OHVDaJvBk2MX74S9EQAXe+cR7AtqSUY3d
Y0I22hT2Y75we4DNzZAMsWi5G7xlFsRITp6zV0bA3EkhARMVLUKMBD2sIxfB
WxD7YGbMPEmNetFmL+MhJ9ejCcX6MNbroYCRO5zEA+IOtPbwcDf1hYTaUjgM
rrZhunvzgq5uAdlRTddijPSO96WIOOuypZ3K4aMtD7uFx0xCn/HYy3FxwV4L
jtomMAuhrWsZ51DV2e0vIhBPRIZkKG6hRZi9f7zRDqwimJIPivkR4HeZyJOC
GchjOwe4GmC2TUbg0VcHVqt06VPan/fYzKai1kDeQ78N8BZkZ1ruPBc3WHIQ
IQSHc9nm0dqLFKmQYOl+tqmqoyp86jWTBeQcc36F4BKFo/MabidGx9MfkFnK
ErMnT3VeQc3zfh2N7cLLBcEe5ui4akYzsU4biXFGgqyrV4HfF49sTKqIP8qT
7iP1pbjxpHJ999ApXJingt0MJ/YFO9SOPHf4sA4Q/OfUNzuIw7GxFCx1fHHK
35Akjo4omj/7r1PWHB8DIUNUWA7njfxdEkk+K/sEXcjSuPWqQjInjxPjAG5B
m1TwJ9pknfWLlM9d0hq8odA2Y2DdWXYxuLV9RTcnyEDRUzMKAqFYjQJjjNMW
pgR2a2JvqJqssVOAAbbkrNEYFvyOsvGNs3VbhkwBBS7rYIAEE+6N+UTN/scn
+GrxZJ/HZZyHfc8sFWou+aXrJwERpZ5Lh1OVkN5DqhT8COo1qVMHpBeODYzd
oigwX+aa9DgzYt0u8+0GU5zcfNS5onOoH1uv6kzYXlfZu2I9OkXCdyWAEzlx
uESbNcwGyaf1l/nE0fddehrvvz9R8NO2pSj8inQElNAPyjUr6E3B5YOc5Lhf
bUJINQ2D6IijaSiFEgrHtjqw7owrs+S/5aoVlwSSfGZn1gYYXN4yvfUpCUyZ
0Ofcb7mDFF81Igs32hOBuF+KfZz+YZVt7K7Xq6qt3jG3/MvKTrp3RYxK3EC/
LdL3hgAsOPmQrQEh/ijTiNse9SnjaGP2We91OxCHgKFLj+b1DTduYyiclwiS
Nmm1Pgu7Ea42fBa7Q+xB5ksy3b0EtQQFsLAjwVzC1XowEmxOawnjAQNFulMP
c0pPtrETL53FEXXIrMdmcffUc7w2GZTnpSPR+9S6yBasCkaYqJki6LnFIP7g
rJCh1W9+7e+Tt+KpKSadffVLhRWi97izUesI+u0xsMo8abCXmxne+qA0sMiA
ElT5Hl90iFDRZpjwCAtZh0PAg00Rg8DsDChp91EiAIqtkWX2zCHetqH4Jy6K
VW2Ea/LqnWIue7FISl4PpEqAEx6CVLSFozxqWnlmuK7CcAPu+a15kCwcey+t
Nwfr+r6y5i6sbDy5AwFMZwad8MWLhZv+dQgPEUGwf1PIUSKaUA/+hU3rXVXw
FLcUyZjr2tJl63hneFV+vJ5nohURIKWhRxe+lRX6q5Sc+sTYgM6DiyMx2FC/
QaP9axxsbCqbOoFnin9/B8q5vCv5khpFR1HzBo2ViTGGt3gc+BAQ2kwPzc5W
/aVtrJs2j3Ukbhm3sMdPy6VsnRHAsZ0cvMStxMEcrw9n+6tnMrZeuafXI7jQ
WNcIQfBAgTYfsSgWS4JJFHKVPVKCh78f3bAL4J/DmC9+uqOJu48cor5pXzUw
Q1DuBK1K7lbLa/QHMC/FFaITl6sUGLMU2q6qgiMqqlw+9NnSew2XcvnyWKB8
jD6eS07ifzLM+hPVSh7YtHlUFX3G8xNuYDuBgol2lUlUSWpPFPb0VoZeJchW
EXx7HgROSarKGs/xck2P+Cvqhb/Hamzg8IQT7zxSTbOZfIyx7dtMH6Ybuvgh
sSVnLEVIn/xzhGPTFSKaL+KTZQvfVjzzTqvommFdaz/GCxN3m1U9M0sA2bWm
SzFiJOolVbmSxO5gu6T56Jz7IbW4XZqkb0gR40i4qhbgY0dmAspuekieH9jR
NbRw7TjbZvW2uZhUjjhDiisyLzW5mW0WnEdgSpsdGNAcALoZj8Fys8xm20t5
HbZL4U35LNzxjk7OhSAMgxTDyRf86ErY/yL+K2i9WyfGBbhMEke3UwHFDr1L
I0FiYKCU5LHAaW28xsfFdyTPGweTkPSQ21LBEm+mcH8FyNUNDqzBtKvYmMIN
OyjggqiPcwAxHh1axFIuiyxAzEwx207Tk7Uvv77ENuEBxH/2vczZMsHhnYa/
R2++D1Zc3SmR8z5lEHqReJDuBZnrqhkgmTUWO92vmiBwjE0iosBdHKeKdNkt
tu+ZO1uPajZ73oCPChLXMfx5SNK2/o4AZazXc5bPr7oHekRB2CNnMLIB3F1r
+kahBKGYhaX6mUEiGEAzxPVHFvR+4wLei/Rk6Kzlz8GkJAX+BNXiQ+anVOR6
TzHUyF+7htl/ekFXr7zC7ocsLGIwgVr1ZwABxfY7JyEB7HmFbkk7XQSbV+3O
2bUk9aZOCquj5dMIfY9NRNIH0FAkhO8PmAnvaKf5KqKxugiTaHJp0gtEEQY0
jGzyBEQwe5Q9b3t2ObkSLkOCKhLhzggmmvS4z2OH/Uwk0Vhp7o61KTHLzaVj
RBXGSKk0czFWaecijG7VeDMQCJgY4PofdxvZwftm3eECLfAfdoHrEXSZfsTZ
nWdwWCk1i6HukMXUd80rrnfc6aWvg2VdTD2Tz4MvsW0R1blaA/cqrTnKjv4x
tHkGYxZrTUgf5u37DiXMctj4xL8lnNQHzm4BOjFZt39j1/hVwG033aFTjwxV
KezON8KJ1XXBMZxkULnMsVskj3/VB4slAsxY1D+ZqAvFrjsFKjfrDKeuSQUl
5Q6mdd5W3eB8SQ98r9IIGXWYKspNgDQ7TVGz5otMPjxFEYX/i6F0JOwtVpbw
gOaz9YWuTJBV247ALtmfV5+VBe7tHYY6/GdjYYYB289m1FLLvGd+DDETeXT6
DLOlneIKm6SodauDjhvVS1I/tNxxgWv3lDInIgKf37Jbu9OBE6wv86GaIdkR
/n9FGveCC+XRatjqzOi/bmi6aMntPX6+lvnRMr2hMnndMQBaUGvsTar6A74/
t6N/wYQKpUU7vn2sIITDCU3O+3B62fUrFydTI9gXK4rS15uPNG+f6W+D1eBF
sNQUHT4TrBvzo9bqpsWh+DIjKMqzBZ7Wtp7hfoQuInZafqi7btRUq+3S8Llq
tVFwyw6QV73jRWoJxNM6XW8ztS3hPMZgrEFP4aLK682CE+TKU/XuR2dYsUOd
mvjf1ySnJxg++elRuMETjxevSFtYvGkifzVC20WUNz/GuLKbaX55sUPx0jWl
qXr+o0lA9JTMMydI0DXn7MQi6Nrnfikj+KcxKJCDK4Im2uMVN3Tj4584gJ+U
qyzcO9jivFLrVhHclBY1rNf6Yr3fwdOfd3Qo0BqzdidOqD/xMy0p1Oty/oJG
FgsQgku+tQHfqMFuPqjMO78PZwF3rhPxtnl5WtR5ujLsjXqLsJm7awCWIdPy
G/O1d8iXX6aOIPXa/U+T4JYD0+P9TulcAR+sqakIMo3xpjNcnkxt5o8HBDNl
/gON4QIPN+PytZrIfqgbc1A+pbboiZgtgsLldRPXo21ZI4s4Ud10HDf43GWh
bukB/vhzwMPypb1di0WL0LNXN3Rgg1LL7BfGPJCm5wU1BLXb4Y0v18dLrvWT
doQ17XKkjIAUVhkHxB4isFonxcMl/U9f4gW0HVTWLkHvLQFQ8fqusmY5hKir
1Z9RRq2Wj1B8J78rvpVfbezaD3nbt2fjNiT1PjS8qleM3RGTX8RYICaWWS8L
k8NkL3pG2lG78+bfa9nHbRoM85srQ6lnB8yOow2VA+BpRQ8hVWmNihbWaBR8
nQTUIoN6yoFbB/kfrWc86f0Ws8QFIqgCKbBuNb+4QlsXV3aOdF3NxdjvOYwu
bwO38E1h3rk/giq55RvdrvrwfkeWliVRXilNoXkibDHoeQz5s7dFfu+jOLg7
CI/XpoFCeoESZK7GnSYoCebBJ6e41qEtPxILdB0s3srSMiha68MtYgvzBt/i
fKXmRD/SGfXCzm6PAgtTYN5naOzbBYKcAIZMvNGaQCofXagEnzhZPQhL2Y40
efyW0R9JzL46ZpmClQVV3s7S7lAZ9nytFHkhN8dNlH+8QvU2n8jxPDdrjLLG
zstOCjchhMoZXXuyVz3cwAS2lR1ucMaLfu9+Azb5Kl69HuLgmifh4i5iq87P
00UERvZR6Q1dvqkf2RpuQlRs8fZpHeC+kxML0FRQeYy0k6qpSLU/oOkcJta5
O7CmFy/U+xevcVH6g5igRIN+4U07QidlB/2AqOpxUDJBLCpOgZcbBZCA8zMU
4A+GBhyZGDcBzBa+NvHLRYs0BlImPt4svlgWazVusiz6oFAvkhqQ4FCsvgyh
ZHbYwJvSc32LsHgcO7TJ/pjHMYdHa9AMeHAInbCqowFddy0UZh/sDqT1gtht
SQhPd50dFOPIDzk34GF2ladP5tBR/TWmpKEp1sgOBrN8xA0Xy0+Hr/DHb1aA
R2PZCmv8UYZrel7uYjqEdN24dVMSVDioHKZ2VkApAr1KM2CNxqe+LU0Exw72
xuq6AguaEPO2XkRqJTNQG/jgQOfzNC5jfc4VhKyJFItokDMYKl4JwPKtCvyE
cUFRlNppl6fnQBTcAQB7txyCZYZ4dfYbcGmZvVj2VCheOLM2Mb7HWrKveaZk
rEpnN2EFoBlNwtI+hh5TQZGyTy7VPOdB12X5qQzWeRxKyuFVkSg3uzMdSQvi
NL0VLiulUG9W0mf5sjOdJNYHAp6oLrg4ciidemVLrvqg2p9+AfFnEjHXI99b
gSWQ4SiQ4TjVC3sQh3OwrrcjbLvVvsktVm8G6v2qCRDw8FozPaMh75wUTPL5
uC7Xt6bBah4hgVqtc5Oin4X1j3R9ROaZ53vws+hN5q49zsvvFY6NyXmDc14R
+aHHK67qaojVem40g3JsLVo9TCCs2exksSKl3tyGv4YkMWVh8zDPcWilEZrQ
LaVXvNtHRUfw7/2jlAF+3a7dXGTtYYNbpgVLt0ll6tMvFwQbX84e32WxJrr5
T57YxDtAAuMtJDAjP7s767sMoUqk3SJtxAFOPDVgrqpXrRjjXMm6CVzHohh1
JmGhzggc35VHGu9sOgp/ITUFHbDiPyu2aBJdOQm4CTULSPZ7tU/PBdz0ifrz
aymF9/RjfDSrHr3HXzWvNSl8VP970HkrjcwbWXqSLqFHDUylS1Vhfvj8hvls
2TnNKrVgDrvfLiauxJ7AEXrHywxuDCCaChED+mpNFTtYPXcEPkBVs8fRYtcy
nL6bMotV9wunV1ORNrbug2iq1cgS1wULgbQvxUUfC468GnQsaqQ2yZYwjPFg
xBU3qyhrC44/LMcuIa+ZanNAPk50jJ2Lgc+sTgB3MI+Lw+3ZUywZxsBFW/RX
vdG6jYdUei9TIEceltOLX3khh9OfDPy7jLdq1tTgmfst9IXHJUOoXA7fbePp
6kww0g0L+aztQ0MydonaaxLvhWotNDOP/lsXgv43+dnMZTtRX1ELMiXoss1g
XhOS9wPooPVTK4XE0CsXGQX+H90t6Psu+FubI+ObeMeoPAHGeGme4m80YJBH
7Bo5VSysFFRlS327k3UM/hnt5jaoeqQ5MJxX8olIEjX6hs8cDMxFiFGFadxH
ga3ACEN5sSx2lf3bEjvDie8sKI/CegLSMp0/KZYjEaR8hUCpqQ3GR+MfaPi/
uLLmY+HUG7qbJV9MFXbvYcEmexHCDQt/av6LNvhrfLwyoxETtjqWVpYJqF05
NywiBzz6ESMuviswf+wDGnEXWBU65ZNU1/jfJSsmRCwlqKbymL1RyQqfEeaK
+MMzbdGFVJ9GXn1w4IwBDvwQ5gU2Z73dJyeXT7Av/sVrHIzsjV/g6ryKdK5v
v5/SNtIgRCdVnjx37GmBOFz0GvOSXEwrz1KeGL9tmPmNkDFxObvM405twaQh
BbMmLTABLE5GVY0NufwI2F+5IZc8Jfcq7Uu8zkhUh0QNmj0KRapIbd3C1Y+X
K8YTtdzb/HDCHmZaVb/BAvHrCIh8xgtddbfSNQ7KJyJv08qbWkT3TeIP9r4c
7Q/6euSRl9/NePUepyemnHbClSnoJ4S2tdQkLkbuQtkBYrxJOCNQM/PZhiPr
uwF6rRKuNFcGH7tP4jyK5AU4ZlsQe1omovQoXTucTjqLKMosgHNVOMGz0jnB
OoY1UALdMZ0hIAF7MCUujuBRUMCwPUnED7kEaI0RU3MgZtTXaqOHAgd4xKKT
fSO23tCqmRlXIqieuYfL3DlZh5JG+flOz+f4eWP+eESCzQb5m4cKsEdCCCL3
ZEGqfnFtTB7Tn/8fUu8ZLzCXmzLnW1550j37SV9opqLivCZ3Oyq9eoCSZ+ly
UfIZbt87HsWSCrLcTBWVT2A70M5r22epfPHOTwBmh9hw4HjB0GeVz8A1JqK/
jS3A1+BE0T6m6OdTJnaA85FFZCGK939Er86ZQt4KKten2cLaxlISpM4zCzb0
VuAmnw115ui/4ADIyTGEXx+s9egH6URWdB0oCFOLNTt7wSVrLFQKfxGf8I0K
WbvX//vb6APyAVaUr+x5eIA20CdDMBLr40KxtPGF4c9pAx+FtR/9s96HYPmg
AstyQjyHCO88RIetAxN5VeDh7Byo0/XkyKY9XdXTs+uJndkRQ0zt9nVs6gWO
KJSL34OW6GpifvpTN8fA++rNjAAaLWzAkJ969qKWxkeARMU6D9BDniyGGl0F
3b491gezhePEklnC9tP9w/SpVhYaVz0qEA2PZ/sYyCZ58GGlDpMYOXern2Yq
U0MxMttvLhHdexbr6uP2uxFQ2aqwoM99xnRFwgEr0e+my80YCrQoKIEDjnWf
JLcSZ4eA6TVmkP4o3elnD9YMPW2MssQJ24N5IsVMs9z+xu4WpiiuwIVoaGIP
Nste2aqZmsMSsGZhtqOMg6BZuslbFxf2oU4GpiOkBV44YvXmzh3GZ+h8YxFK
hBqGvnNcKmCguGeM3HHfEosxjQ/FRvg2NL4wLnecPHCJN3N+B25oEwBb5d/2
TezT9jGoV9hoZQ/fy8QMkeVsY9cvxMvI7ORjCbpE8j9Bx/kUz7EY+vEMSygx
UqIz51VmI5cXlKyoPcogYBu+bSbPGTTZN1bi3HTndj6KBPoYQICbUWplyKKZ
13D1+61UrnFK7h+uqO5HQJ9619ebArn3ATj4f+2iNak7XJZa/udlth4UakHi
XGIO1XnSleZUAP1ZNH2a+v/KIXJHplbz8NmCB1zbHyWSxPBmHyYos5o02f9F
WDGeJ7KOrGKyjSdgovvjUNGkL30WDUf1p1nlxwqRIN2mdGR4f5GmEvSyciL4
njO2+/+Ta4/w5scufD7qXRO+JmMJUwOy1k5Pw5tiJ7GapjVlbHjEgVQHd0ZL
I2Tcc/1xq1aT+Yvo64MIbCmUYUDUutKMg0V1werGgiXkjLqQicD7bwwcukbT
Q6+YKzepNPRV6RUDX5M/RSYmPxhuBhj7t3WSKvqXqLg8DYIzxB6Nx+W89CVv
I30a3giJl1oiqyKj9/RJlQ6UWxqEdQxpFAD1z0aU2/OQ8kuAZhjFxig29ZQ2
ri1TdaO+pzWEMbm6OunuaXaR+0ccZtzCwxAPsr7YibdRilzBc8NyqBnYmks9
4j3DytxwT2QTXqv9OO2cujRa+YK+mYSOcLYjwgMNlCy+jNpCrmMxZzmG2N1p
fUF6hyKXeMhy760sJPC0YRoPKknxPzobzUoEGvc7iCAWMVsVQe4oS6gU8bcG
14xXAZs82zEjat13JYi2413ZX9mrC9dtN+rxEKzQKYnxoDiATxUVpyIkpGYh
x5yL0a3Kpqj4sTDw26PczIJp2WPFnJvSaJj3nnEFMbWmgS0+zd4saphCDy5Q
lvK1RDEwwhIifEjolmzrvijjRuhYTh5UFOUoREXqHndeV26I7/68XBAzSl/b
+NK3C1ZpCgALKK+mvmMMAISqb3VpVX0zArM6QjRpxOG/rF13608N2g1sv+r+
g91csEdhwTZqSOSMDXW/jO6yil/xX2XZlLAKrLNVuitYJtbGkKZXjHm6iisZ
oglJOXrre0tC7iDwlQGEYmxL01GxNGHLpBwlmmGQ62NzLwuRq87Q+qc2PYsN
hT201swyQxRP5uvDIlKLH4Z6rqckrl0Kd3YUBa6WYhFXbbDqagppL+0r8Ne6
h68RIpc6n+KU7Z3k4uaNCizou2gjw5+Z76jL18OwWSqFZ2V+U+ydVUS/jDZ1
SIZxrbue3IduB6WiqqJukvggVGDgYfQEg1HviyhjdfcBPDPvb/m/slSUFxWr
Tkm9hCsOeb1qJKWZIinuVVZYCRX+g2krwEH3MYbRUahOJZ68OmeEp8OYHgbU
+4r4DcsoCqPs+Z2+qao4hU+LYkxmMg+B5sbRycGcpozFheYyj0n4CWvkpgq5
MdByLwhR4J3Fuc1EP6KKfyQeEYihPTS7qyd9a7bna8VEIQaNIxAj037Y4lCd
LXLDQRPp5C9GB+V4ptyRRoVmG1gkTr7BhB7khooGsW1LVpg77uk3t0ftdW6N
GXYGEXWSIH75gs7gsDbcve+NbkGllnnYDk3nrWQr245KMsUkTTeyvoWDdyDO
2W0TqCJcaeQE+2RPsW+Dn11PEIvoDS/uaIqku6EgDhNI43TzRVTpiUhsO0Cp
ELjvYu9FkuQl8avuKPdTqvrsS9MNKeU30ZYfbym/P9bSKLne/prhSffS6HPo
s15nEsxBUdJQkDacbOr55WSqIl3g4DBUZJ5v7cCtR5IerEAX1DK8NX3qljqM
ediIrjT0WN4yvSOKpzmE59kuYkBh6vOwQ/nDHAQ27jSFN8LLPgGZ9Etj9Lfm
BtgEdn7tiYbWKAOFHwKXc7CJ6e6cy6QszmIpVx6cvBfASpXmNhtTelPxpeNX
LMIKI35zZoNNXtme1hNUPVXeOuN1h9/lrLUL9KUNCs4sQr0cZjslRPtMYsFG
eMoqbte/NMcJ18vzpro86pLluFu2iSm+/I7dw3h1tmS8PNi8IHJqfZ+jVZdV
xo4wMLyqNJQWvKgRdCIpMykcoI1lbAP1RZzNI/R+YpISfqqHyD/tSPrOCKLZ
kzMr8VXPSEeuHWZwSuFxOfreP7TSG9aveUZ4fTMgIA1noyLWwhQIfNOl5Rvi
r6BR7rGAEaYVgQHPtISj5/4CEZd93pT88+Po7N4N8K9B7222lfwn0hPHn5LI
FokiGh6uCNflUtD2Ej8D1xDQynyaFeJRhW76ztXyO5SsP/ZsUqMzL0bFv118
sTWUYIknOEBKlAA3fMMrX+w8Wi0aDFw2uUg4Exvmw6vTNQ50UhVnzJKqpRLi
RJFF8kLExTJ87jGY5bphgcmMpM+Vv9Dx8ZmF0ksBc7CeGhkDLq9Uw7uQijfJ
nKjvGuJZZg4nmkTuI9/kW7qvjGqDZ4Bb0p14RnHRmrb3j8K5IbvSkjU7ffWW
aCl1gh89XhsmMAoLqXC/6xDW4SlOrDYK8rnZnF74GlWX6htLqT2KW+r/Hp4w
G8vGCFeaNxSZu570DkuFqMIXhqFLMtex5qkhua7N6CTgekxYION8QoUyJArC
0qrZ3l/3AT7hCPu2OYW+K2+jlN5q8yLRciedwhtrAdKcD2wBHMp9z8pnMhR1
b2zmOwx8DOiE7mVlmcaQYzRNnZHyV0NECo6Czl5DFhu+DMOYWL0lVS98NRC2
bmi52ETUUpte0zzhYjNR+CQX8bZ+2DvoVd+17F7k3VD3pc3QiU9TzXYxbm7Q
SGf5wCrBk0mQ0J/t7P0RVMO0wZtCJovrJYnOyNakZtMFmCSaKerSkx+LzM2i
79w4Uovjz55DqW8FcQ9303eP2rCoG8PI6vEJOySa9uiszWXQo5XF5spIOiUo
gEpHwQKMVOZDmI+MIFvQeFZQFe3wf5PGGnh+G2xDuVfF9k8mSVts46GpRNZZ
4EeJMxnhRFLy9So+1sT8L+RenuDarvzV0+Y7OXim7FB1UWDMi2STXjnQ3zxW
oXuJP/vun9T1/KEXiEsNkJMafz7QezZBEfnu3xBteV1CdHoT9AdvI65+l2Iz
YnO+RAv6OjMObj7XHT+q7bT7BdMIf4rmyoNyymz4EeVEUYh2gpwmEllIUf4J
KQg2gOMSLppmuDcnQHHYCzTVgzA28tx8L97LqunVCPpLeMLNOggRV7vKF5UP
2YvS08Y8mSwTSjvVyushE4cG7Un8UC+skAPwrK49cdB+Yh/m76BdoN9DCdHn
b4wUqeRnKquNFYwbXCLbFzm3hGHjscUHmahLQ6jIY8i32s6ytYvEoqmC+3th
Wbd5+wx3xAdVHP1r86k7CmwapJPDC8h9VHBONsMjFhJTPuIh6q68N3hErw4/
Seuu/cP4rb/0K9Ja0XYrIuFV6EE7xJ208ez5uwbHo/JXkwJuQt9H7Cx6L0KP
4FCClGrb2ygYP2FUOEyMq0aB/q955PBDGbqn5wkuTn6K0u5ZZUo+u2O07x7y
sZeNXmlv+QCBQjM/kKzlvveC3r6KkuEX5hw0SWTse7AQggrarmLvLy4dSh5m
6c1ybp+4wbzTJQrMVwhPAIQ0Z0If7MbYPxvOUzyiTyBkKxrgcbar1BZNzXfg
87mgBvDxs4bKMxRLJsV2xaCRiOeOWMT3dXP2FtGTAVu1v7DuUXkMPpMiErUu
vEfMElw/pxZwXdeCA/gy1d/WmjxSjEva8kNlWwfA8bxNCgH2/8ajvruA6I5R
mwOQZlYCaQXyk/O62lee3+txkggD/+Zoha7kf/OHnO91bGrD0UoHUXRFWuIx
MQ7eXlgnX2lNR2cWsvZ85hj0OKJ6+iuRKg2HUPWa/9EZ7x0mqhuYbQ9xEemA
IYX95o//wl4YsqtY2sgJyLLu7S16clfeMgPnOIU32V2AMiZz0hVDdoa6OFRW
14V9VdSnA45MflMmYycVuVQJB578BYStM1VyrG8M4/qGgdO/lnKyxPkYWdpq
3+AfmqVKvIa9RVWSNa2FAZLppRbLfBjrJT0/oyuEgPU8rXscrDirDp07lSLz
XxvDtesKIXsqoeJ+EB/K5klRizlD6KuRTKeYIIAzBy3T98WGuGUhm5TOKJ9I
dVE8F3bXDYqChg+QJj4kRDp51ElTKJWbuCGiVRPQvfdPJXvsU1ELjs3B8mus
kC7gfSzGDbXGAhbi6Q2gl/qYFtAUj/0eNgsoZruae0Y9IMsxOc76cau5XpqJ
yfXh9jMLPiKwjWGmbCOPA1mx/u8Ejl10SKjHv85mwlWrH71uEKOsYk0o18YA
hyieflg86hplnm9ZHkSSoVsJSvZ4z3jrxAyRyNy9hKPOyFW7EjK4RtqkvXow
jFp40KBIrOm4AkIEW2foY+bK2/1y9kZbVsSLKxa6roQJxp5yIUmpReKfcKpR
zfgltCd3bLnR+XKoQmF3IrEkDN7nI+8xqSDLtkte2I+6YbnETd90ojVdbHnq
cqQnTonFaN2t2U9afyr9aPvVGNY2cn6HKH4b+gJtvSU0jXmlXiELUavT2m23
fd1qhSanzpQnfmVwceQ5d5yudQDenQaFXYcMvb++/IZY/a7Ya+HXTd/Mzegn
1bk5iNdq6tjw/D4qYMlUwoMNvvGc+V8GHFeewiLgs3OCxGx11mVLJg7LvQWC
vu+2m5k3zlB0QnVBVHfru4Vea/YKEyigDzn3yHXBaN3DYV8NdFetJJ8UsU6R
jKw65I7zr3JUD6s/H4AvTzECuVXrZY2cRuPxggsm46089sGGvGl8SCiSvT7s
DR4ew//BbVyypdDe1JfsrrTLckr7sbhfDa1IMGBhHaEVMBxhHa/6+UxkhmRS
XAXFxxe+e3YdQeInIuIgIkOmkcpl0En5BwPiwQoloTuB1+BVKrhRYCPj1UWv
FT+xBYb4DAS0we7O/fbQhjT1pWIip6Q72TXUd5DV4BNSgCet0VGVtoM1J6Mn
npsC0o6yH1Cojtyll8gIlJ+wW8QQXLj5Vbx8+Wu0QwsBXo2v5wGxq+fPljge
2W6ROWiQ0IUQmCNJ2ckF1twlw7YNBxqRb/vQwovTamtqsBJ86iCs6ucukU11
yl3sYUQdbU/F+IG4BBH+Plw0pEi5v1jmqSUXHwDbhn9a+cWVEaV+lLHdphtO
EQ2k92buf9zyXoJax/9jmRfQwSbiHqR9ANhUsJxkaAZyBkqrY39NahIVPTMa
E+RyLZtaoBRp4B4kiLlJch+d2z3zySprqJleYG4+DpVGHNSrSV7K8xVUpFBa
EuHePnnDL+uFxeooGMhEw7VD9SUK6d3CCE0szxn2R2XqAG9AXqcjpf49h0g8
wvgvKqwH0AN3mNaWCAIklwJeK0fvwABSzaDOdXM4nsivf7HFAXKqnsdmeGns
HgfZpC77t1DORiXKhalR5lwLLiGG7n0qFWx6KAx31Y85GnYidcT3fHVUqYKl
fKc/gllY+1OF4fjwiajj6Px5ZppF6Ef9iZvr1JwVp8yx49uuYdH98EpVdmB6
yZll6rgu9uSVI3Mo9/iGtaiNOVjM+0BXyASjtk/9ZZTpV/sL4kNEwTOCYo9X
YPjtjb6jroYpB7Q+eLAB7yiZdE29Jf8lSaXD7b1+5o5DD0YxoHd+MqejFvBj
tNdHXsyYWBkSB6A5Pu5wRjUwlQKDpIeHdANHdb9PFkLZeCz7xxme3f0zWP0G
812iPruJpx561+lFE4G4bBPnBjS06m0/XVgFhURizpsml3R4Z8/gW2epAJWJ
inMUGPP1qipNH8EorfHVe3t1eUJsBy40DJg98kmOVkXcH119TvsuMxAMa0eT
cEWgyTX6vGaIrewXd9CysOUQXjQx6cz23mVCO9Jo0GZ7mXW/4yASAsyOX6e2
BmivFpPwo6TEVsVdVrkv3ZXOIWMOBfOlN2KdHCWafmn9GD9MbwoRuPcaH2E8
sehyB0rOWUUWIg/yx0i4WsNxk6np018Ugspzv0WCDkNtOItn1yJiW+bfS6qm
0jPE3kVeG1Nbm7mLJxtr5qGqDa99SdvOZSIEZ8e+D+4h3GnA0rflkYGgFNXN
Fl42zWimxnDOjaiSDqwGPRUOnJ9luoX8i06Ay7OJySvt7LaBp08qFRf4SVtD
9fjt5CRWv5bIcIPcWT+8B4UfbmUKAWeSPUbgyOoDBqikmxtQOb5Q23flzObh
0QBylIGCQ9hubmFLc8MtbSRlBn/yYaRJlyxRyo3k4bXKRNLjsnu+brKEDghY
6KDWQLat57BeaMKRyzK+YYbya2XxUc+Oo9rSHsiWPnb6IwKeOqStAAtIemrl
CVeqDq9Fqhf52or4m4yXf8pWFSvd4+xKQIxk6uffdj7ijnyxXzI4vVE0kyep
UwOyiuGMDBbukrDqptCgCRdeI4t/SVjUv3qhqaSLyawWYMfrF81fz63A8lze
qxVqmasLGY2ulAcGBlO6gENNF5fiXowHkpsEJVKEa41ILX1x/6vS/SgMGaqP
QifQ1DenAEx5ydJUoM1SD3Rye0o54uShcCjrB8ODhVyN/bDspVrkaaY/LBWQ
/WQl7GcRKFfcOzI8M6ACe9HkuXsDI9fAv0k7FcVoDuCWrXHQfKydQ3arulXV
gJJZ9tV4/sl6Z6Gjv3pN7zwJ8Z22EywxMc3u5FquGsRQJUc7u8DLOMywiTT0
APs7nEZZvEd7ybpcU9Fk4ROXjuX4YaKxKMVuWc9gkqsCPRoMPqItXDJt5Jsk
voBruvytiDt8gREwRUNOIwHqJT8Ilr0hzEiwWJ4FJgsp/Bj1NM1BBcXMgA9F
8IJ6bQaH+isBJykqg8ahmDXz5ofbKBJPeDP5jNIT6sPCWl/OUW7dHbh67eCQ
Ussew0no+QtFR0fIWACHaESikNgABRWYOkIYDMMNjOjSOBn9Gz678P0tToIq
gI+F6TNmXNOkYpn6SKwUpf3t/f80Mssnxm3tyorQWEmBsWZ21MDGvLn126mt
/IMcJlQTsJWvH9FI6wITiydxJ10xwSouHxRMAPf2p/656KspfZ8YZ08mKPWI
uFUKrH7wYyzouMrnYJby/T2DDDNMAzYyIaVswMvHO48YHhiSSdAoJEW+4nqk
VmHEgGH25fCc9xL/6FFgmosqXLSWNOixfhUbyy557X1QkFY1ckOynCgcxBAt
BV+f7RtkJwzlPFtEaqDH/9kef3yKxWeIMesJHwre1G4N8hOqdzg4A3XbgFIL
9kq3x8syMHGgM1zYpJZqp0wsPoEYngitR/4OymhaDW7SWr4mp7s9sVFwvgr/
UlGL9edowzMVfDE5b/Ut+T5mf0QBF0QkJsTenW0epAyL9rntNI37znfAN4l+
OyZKWse2fNVUKPgddS6Xcuee1MoeUIBGJEb1xjBVNEgFR40PSjFP6Gha6VIe
YcjSVE9FcnvbatEy2vYRxYm6vtrfl8zgjgIk8XElRS6dRhbooch3D44BD4It
yNf8ewRsIXfApHxhf8uRxkyJ9yO9DNyd7tXkif3IGbliyKdQxK4J5d9QzdDV
cWocVeMo2hAAmNsPsmmpTw++7ZOknZhr66jqOubwnH6rQ7vBKAJy/YsIOUVi
VuhyF3AsEV5gg9n3N7r8oZAC89qjZgGkNdhOQXmyHGo0gg2XOw39kTUQ9PzE
xDyXLxaiJUvblCwdRmBFIc9NiIOt4C6xP9A6EsXCjBF2PG3bUzBCYnIM73Qb
LOOY5gvttUO2Z//KAN5IsKlU1W/gTqSt/jhD10aUWUp8bX66ZUll9j5yQ4aa
je8tT4QNUOEsFIoVPIHvTaqJeRVeEGNL26dZZQUeUC9ETSEgkz9xakyr2o4w
MI9m/FVMnSnVL1s+oTl+R6EAPk/JZVPefnptLbtI+nyHDRP/n0D5mT46wVGV
m1VJkuT4/6CN+oQoUnUFcbt4NXL1LzWge9NSollX6e3VaN8ZBf2xpt6DQpaM
mFUIP+67dVwp/Nz/xiTgrqxGOlLv4SI6x+JzCYCkvAkvQmILeuXNkNTCt9v9
et1XqChKiahSi8eOZ4XhkJjno3i85Kt0/CJsqQDtrEK3IhMM8jf7SZci/jJX
C9F7FvI=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+Eqc2kVBHE3sAx04bULChhL4TSFw37vw3SrmV12HeGjYg0vMYPLjF8kojZCn9D2VEKeIPALOzNWKrxcBLlA0u2ZyB6XRvE3Nu9c1IDjDplQYOKkt7uDdFfk98dZXlHVgblUUazTgRHQ2azf1xL6sNd1GnMijzWhE/bjEBZO74Te1cGDNHDv1RiRZfxGmmuobxpngsLWhMLfM3CofzSSmyjqC42sHVi040Ufnza81bnGl6QfFoHHxq+S/3NpRkaZBMCrPAiYHQcjMbyFK3TEzQgutk+azSz8woyiRrLFyBvzP9YcmGcVmCm3VZ64QDk/1+phaYH083sRM7vQmfUJWSEgGi5kwbi1X0Oj7+kmN9aKW8OzyRrurNkg48BxXPJ/TNjcbTvK6KTrsNgI7+505WD731LbWMBBu75tBs5niQ6Fr35xSGn0QaSfxKoUauLqUSHzbwWsnF4D4i9zkIT7ejyBiwRgcUVxLZuZJv3s41wx7fKqqkMECtb2PhxZbfSW+2deSvOWOC6ZQerLFNtHoOE2eEcxq6tq+BU8q7M7QVOlfu7vqhkXnYpbuYq1KG1yeNJl8FXhbePBIo4vuumtmPbj6BQseCY0DaB844AUMYoB9Wcv8HHVZIfpilhodJ/0SUefJ/NnJegIZGS2bdxxd3pf1qKvCx8FW5mMOOHXHGZw1Hf0UBx1UJ1twbJXE6uc8WDyDrXqx/0nRbZci08RX2uhYRH1F8V85BLj7v5fa834kv/VN6RBJlxPSELK2EXxmBYxffTnN76ipuIfr1eQzefud"
`endif