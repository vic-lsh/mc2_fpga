// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OXawStC15DCACj73CA1DO5AT4jrJ4CyRlBWnU3IspgobAka/8AGZWVEHUlHB
AWkpSbjPeJ+uPqTWj9Yizz0rSX/x3R/vQFkiNIHavT/7cV8LPVA0TXAekeUl
swXrh+wHs8YiggeOVMl3Kxy19gEkKR0eWKUwPu4Y5ZdfYH9giR7W2c2Q0org
T3urT1S00jB3bguFdrWBaOEhZkFFGT2Xy6pJL+zqBzfj3a/kGCNty2yvGjQC
w0J+W8VIlIlVOMJwb+tlHkeSP4Dt/qRCN6C5kmixUQvMKetRjaw5qVh3ppPh
RwDXH+mjjEHk4fe6kjgky5U5gjWa4mIAduifjvyGyA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UTYaTIR45z5xaZp8009epZSaOqJHyK2s1HD10McrE3ixa12gqIDHBPYehGNW
PZDM+B0KzJDaeQUN1tyqzdH+VDs7HuGAsor2SHDu5m1X5lwHmMKzfv49vuvh
6uCRdHBKaFwmhvVyi315dIG8gJUd0fWisF6s1VkQNblMXes4WYdounyRjJPZ
HchYO08E7EbJAvyo1qsi6BrfRx5aGOOXLgdjMa5sOayjpk5KZbBe79R/cIdb
zbal42iF7jQSkTPHbaTcN9dmhUg5V74ZtyHeplrEwkuQT+EkdgxwLjFvXkZd
RYBvi6F6sG1YgV3noAqpKn8d1sxJq2L4mjqeDmZxDQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
utbRU/p01xN7NN0n4yr0jgs6H1rBbLHi4I9WUGMfvBUf7Y00/XYEmQvzYdPx
BM66xQVit/koni8TsJafcKE9UBRV4GvkuzSem7HlyYgdbwnqZV5gecmrmmav
W1PCR8IY6Eh6F9jYt86xJhT2UC13rH8CV55LfGXSxPO8OUAIPyoIi3eF0cjl
VPxArxVU4IwJJ/Z+KG0iZrmhleD52hB5YNTRNDo+5AVY6MF5eVhw4gg4dKVu
MHsyzw8po3NIknJsaw+PkD65/hqSAV/tiHO8TF/7P+ifBSXtpuCQ6Cwa5CO8
lz6sXdRtjJUxZPC4/LTC2gLVXMXqUp/O7vRrPqBMeQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
F9bEPobyPHDt5xfb3gUyveNJdcliXJI4+aJMa1i9VgTr7xs71ALedXvbguBT
abi+aTUxy/GwHRKVnTvgVjj3XZZvJEgOZ9q7o7MmtbiTJaipNYyFu265zt6O
Aim0eNsppZebE4TmXuDvYtDh8RyqhpEqQ1EFcTDhcQVcAfPBMGQQo6uXOVzu
/e889XJqKMOP8f+f/GTCyW669Wo7bna2GWXAwJgl2KqJGkOccbTZTid00ffm
6ryIWLKlmgh67HR6UXjYn6994/nzxJPhRPOrwevn+YS47rXUIVSdK73C7SDk
IXtTfv/q0uSMGWYocKf6SJnq6dVUF7xNyopbSaRgvA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MVPaOGV4eLiAZppqpN/9kQIfbn0oqh3QI6yus8YAMQ9218MOIpOBXC68H24h
sFtyPXJipnnGw5bOYRRAi9SMDV4SgG1Dneu67gNu4mloebGU/gySfrM7ubdP
cJ+GyAO6pbU/yp6dKTOT6ukDW672kh5ccg/u5nt9mIPdmE7QC8w=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
b3bF1js+bDfMWWDmWhw3ltM91ufsccXkTguSCw+BOP8pEni04aseZd5SIjwn
oYF6PvF/BwL9IUtRZxZ50D5xfkXMo/nvYTG69K8ZHBUouTqTfepj9zu1Ir6O
9NEc8SBAVfnrwYEQ201XdEuwvVmlwgjsnIzmxXA6WWJnTNZ2/eDR7N6sCdST
ofIPHubGY3dxkStum78ImErluG++eiEEsV/Tg+zOz84GQooKCW/DE+Isqu5+
Cn9SKPuuLScNW2PgDaULjHa6SPAriIRqPzdmxISWyeY0nsNEdtP7HmGpmFuh
9HR51kUyKzkjkH8TB84s7WLPLMzfK6E82E9ObV6chkjczTYxVsw86QF1unB8
SXndq6X1LXf2c87aXS2kdbbkXLcqC32l7nnbNNjiGfyJSSVmTaMLPUZu6yMz
w/+h+lH/+3gT0Hre7ogIrAj9e/T+jTr1VMqSlzlw/2UZQBUgyXCfl441Z447
ab9rWkxHK7VjDP/gsVSJMVwJHNQHOJHV


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
a5zkqS8jMaRdmtewSnk1APGmsqjjGa2ehnASVAsVddgs+B1fMEstGAKI2xyk
LRgZf7lAJn5I6ejnamocS/d8CxVFZNM4MAvLHB2C7cJjd9Jm8oIaaAHiPvLH
FROS//HcgCwnFjIYUuxp0BkfB+N1xCTae1Qe3GuQQwxHQz+gTc0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hZfqFNUhqMIMR4rGMDUEbJ4DOHu1NzAFua3WMu2q29tK01B3LT6a/8o+GWFy
J/bCRdnUfjQ/EgkYXnem0akbzl9v7KAtbIxWyO1WEC/ms8kaKS8aHgpWUo66
G2iHrx+70m4XaBRRvPLVKlx4R6sZQWKwV6OYyJdpl6p1Qu5R6vo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 93024)
`pragma protect data_block
WkvA2u0nzc6LS4JIFfD6p2mm3ljZzAgkdXommh7jbM99KoLJbsLCnmVDTixq
hsRc2sA73nsOKtvkID8R2x4p/00My3q3nHw4o2Zb85JnH6YCUIurLsMOaoNv
vVlvTtPJ/KumRZZBDJMzdjGyKEVL6gF3vQu+QaHfSLWdHSdJH3pkHWo3GtIb
sCV2ZqjODMV89BXGRBLLIEAojHr8WrEjynerh722Bpg38CdwdHnEGQM4xIzu
Yw9InnEUfH6ojhkG/bAkw2X+N6H7lBxMKCDeATFsk7D7/GsKsJcxqBCqGeQQ
yhkB2IzKysaqhYDl3tZMxRcZkFa1c+xUDaEJs9j3k202P12cMLSeASoJ0rad
aAlJq/w9wTizCcAH0wWuOMb1o+f91Z4qNfljlBi07YO7RJ4g/tPFxcvDGA6K
1IQrdoq7oQJufc4ZTiz022bswN9Rd4ybB4r/SvTJl4vNxoLQ1GSN+h/7QXvB
z438VRZxiPs9Fr7ensZ//yPRBso9zxyxSTyEacXSz528MtR4dbLEHXM501bm
PlckIsfxORwdKSl6T4oBJyPL0RgmPsiWh/Pso+B+hn0iuoInfkIWmk1QxSfe
QEPX/ENO9Uzx8zlwmDk6gfardwL3eHuC6mEW19eo8vOEUNdAVCc3HN3WLLCf
V581UM+t1VJt6fxrhYlFX+oor5iRVGLAbtaOpDGIomrmVymqDttDg3ythw+N
dgX91fIKbLGtvM67SLcGLmnhh78WBO2yDToKdCMPq8c5dXBNM3nqaKccyO8I
/eJX7Gk2V7vvv/q8jBCgR7CzKaLv89X/giE0B2Rwt5HblFAbQVPokszW4eEv
l5+KT9mXHb4Km7bITDdDyy7c9AUkoJaNLWLAldKJ7XjaM4YAFBNCXNPW4LDq
xbzWQUmBdNC1xhxmeVXlcEPrpMCoMDUsVKlny6JKrgfITYokssl3gz9ahHFb
bwNcuVJaFKP6WMJe0f0FKMFniU+hhIUiBlJxnpZ2DtuDCdjxc0phZ+venHdL
LWyILZtzMl78HIthHxs1uwIx9ZBgsY/L9c/FaCIJxxTSdon8tdXVZEcRgB6v
9zGOD7mdgDTr394hE56Qsc/864STtsa+iupBCwm8CHtWMrVbcST2DCE0d0kZ
AAT+TAPaJhiUptSwAjtKDklvFCaRHU65XM3ZQn7h7AFXJHA1neCCrNlQ35HJ
y7bVptL3KUk03WC0iVj92BJmg6WrODGITAlQI2h+3bveSZifm5E8Svrih4kN
UKw5Ygmxv4yXe+gfOQyCqntUGi581MxhQSJIL6UpnqtweBhEH64vyw/TTZ/k
uVvkrV9QP8mvB1MTHeqdH+HJOPJ+6EN4drVE+Ni+OA8UZb1zQ5wp9he/sN2j
n53W7ZPr8+VNM4DicB98EY9hUVM+Njekdvjnt2lKKWq/FgsN/dVTPhK6+9pS
UpJmU1ezjCsCUTUAeLHgmxI0DmbMYgaWaWefajzCHGflYu0AUkzg39DU/nQE
rBhhzmNvqrWaWzkhie3QOeXRskKLGWV7DUtHljLxWZKihPUPOg6oBFqe6VhE
ugA+kJ7SPqdOAWW4ZYyxAwoG5Blcpctl1U8EaK53BSqe1WT8e8/VyToG3iib
5IC5qrh8vzigYv1SN+mrrTLm1ln3wzlneEPb2cHvz3gS+yQo4sg83/t90ayy
xACCMTtu15eoNMiuR8kPifmvIa6HTKvB8THRtp7I1oFPUi2qQye5Buz/pbHr
WaSHMSdahq+CRAi46V7uwid8VAkQ3xIBt2t9kM+hiWkabTSQZKNyeMKv/kOu
YsQFkJO4bEnvS2jW/JLQ4UDfW4YpLUouIOCMHSWIHcUhfNkibVFAnPsTh0gL
RwprFokbDhRA43BWoC2yCnMRLsMnKl1/74usc/YuaDccJN0hDOZBv/JzFltL
Z7kjQJnfMo6Wa7i24VWgpF5LC5i8AR/ie5VnaLrztX0f3t/WPPCFj2LxDzUm
U7DBbxddzkfBtqh/6tTtEKEQo2MozHFWnFaWPo3uMwvbgsEadPdGSUC9vC64
g5KpGXmnEYiFTxQVgIxQw3dRfIWLGv0AEva9sAWY1/Ml1GsMZhodI3gxeknK
Bl8vt5f9867Zi4WkgGF1rsJRsdqGatl5dmuAMV78oxP7MvV8tWi+HHei+UaZ
HI8CsyjJdRil3tZ/G9HMhybwAkDbnObrSetNgILDv9lR8xXsNn+kWNegH3G8
0QrlE3RaoSwQ7cmVsmOnkb1vlwTrWrQ9aRW4uLpg3ulBJWa5wuD2Xksf3882
3FKB8QMsXuz9GO1WycXoOBXps13NG2dcEQCJVYWRN4v48eXI6sP93ZJ6L/3G
K/wpC+YpFTZGd0PmQWJ0oEr2GRntk8aqmRbnuHw8vhKY3B7ArJF1VKhVEPRl
Ln9xeysCu5qx7HWHStqwys56uvLcDldJe1Bsu526uQ8yBLMDqgBwPAQLu0VG
LtwUs6AXKnzS713xHqH4XXyBnjU+TZ+D7XfJSUcXORvVfbfivKma+VTLdmur
6hBSbPNF2y3bjFXaRfSo75Pj5As6Eih/llQLordHmA5gNoLv7uI8roycC0P1
Cg62TzbwEE3m/rVnc+snYheBRV0X1PyYzshtWBlqxwsF6VGErmeA1OobxdCL
Ndmk8pKDcz35nD7xoAb4oaYKRTkKZArHFWB8s9pVKoVoB2R1DdoYo9Ajsauq
VmJJvI7pv9vBTW6gg7PP2mMjXyFRrtcvuARobl5XFcQSnNsJVCMs9fZQ2doh
gb5bx6jWmHsfg765XqtaG/GH3+rvXs2XPBwULddnFKORral9V3KiOSutQci4
E1cumgmo0M9Awj7ZcvY9wgPTCvYI14NS0ONke6JYzEei/iUN2t0Gn75gTUCj
ElUt5x+fR4WIsS+zr1rz1OKhFNn5gAAwEGN2m8DTdvXaAEbFc87RLU5T5iUP
7pE91e0/PMkf+Tq2D15PnVccl6/wu5cuNDj9OxDyqjWv2rKSloF+n28B/qY7
yb1N+fViZmV+EbsqdoExb6yX8giD05rk2Mj/RPRxTocu8RBpZyU47NcnQNJM
NL1g4//V/nnFxrWkudmO+FDKJxCkvdlxmUpNrVHP76WkGl6JzuWvm//iD5XD
1iTwxNPg6eqYhQRWXyk2Ybj9g9E9DJsYVuy8+61RXdWuZR+JdyCb9I0arF7f
qd4upm8UClrLw3Rz1HGt+UZffi/dGCy4nt7VF5zEVngRzam8SLCwhk20fKDa
hAI1EKv9Xk2gVhv9KatAv+0rAhNX3YCAdG6pA6q9CYNw8HEKpR1EHs74bBDj
rarGwHhxZUZ6ZM2daGW3eTTWaVyMEaN7062ld7aboOjv/BS37Aot74MDT1m/
PUNJ/7czl9aBKX1kxN3gEyu6W89EOUlWRSUey0P+V94GUQVyagvuTWyauAjp
XMSc7dxaho51kVTLKVwaN72ZGhL4/TwwR3EpmKksBUajhF+mJ5tV8VPUiOGs
fLiEMV3Wo4aYk9XaMvyJUM357/Kbj4FAXJ7EUY1Yfsy3AZyyLNJp1mTTARP7
IeqNuyJub6l/2iRSrD5FbLqAaRsZcr66HLBVmy3zzouSd0N+VTx2TWhqv6OY
swJsBEjiaYNo0kykOFYXLHr474LdENpVK++s05o2aoC8OgMUZwtShOk05uP1
0MGC0/XclbdLlBNsYvDJrMqiOlcCCrX48gUcspbz4Zi2Gl6jLIK2fLZuhtEh
4P/6TkNvIe7LXzkDT2kqz6UT1Q+MaUafTCXHstukI16y0G1dYFyXUoN4yPnp
+rKfTTlN/ixCsQ1lVurKAYw4yx1GibQAreRUe6yI+q9l6He2xh/TVgimkei7
0kVsI5R6g4bnDme8xQOYnitYEQ7k7Xnc5l6rfrAaaelEaP0BRVDYd4lW2Caf
SowvMvkqyrRzfvT6i2+kHcASlzXpRispEkWREgbqwndLyWvZxCOyXLd7mhT4
5MFbQMa5Z5+cdzGYQxVqtgbOkUfV0SVrXBbYO627tBkOA8AEg1ktx2II1Gvu
yBp1APlRe0OCbcwXb6thHUp+vAMgwF2ibvF0H6iDKMc1CXt7QGAYqqu87NMx
oxRjQ+pzwr0n5holXUBEVApOzR9H81veqJIOZGrpO4gV/RcQQOtYZW1iK9Vy
HvEm4mfO0r1M+TSPP3+ubgmq1pmWfCUIY0HOhpoT13MdsojusJwyK7m1jcFh
M9pN/t6lAEjG+hLENKK1irwBiZyWK0lq+L1Cv+MalvvFS6cufwUuk/ok/Er9
eEubUoPX7X/lEbnFwSW+eZkIaxc61I8EPRn5E/XoWKiydcy5kwJ0wcy4fe5+
WvQT4vcnPdVNC39sZVYu09ROSYJMbBs6qGrqS2Dcwk7lNvuxyTUuSa56mkYV
C+T82iKwg0NdYl7jr8uYj8slyoC64w7dqz3cMVUGT9ZwGeNnNup6fh2bp7Sa
gHkTa0MPUk+wPstNFuo1EhvLZdbBf/S6t+cA/ICrK5QB0yu8t+clx+bH1iEO
2L/kup2RWjp4JFPa8RLpmPuQD374PPEWAz1SYs890BB8CCEyQyj8SK9acXSn
x7gddC0l4+4AwQYuHiEDgkuw6RoHWPnBDf4jJRHk9g/MOy0x63gRMx/79PmL
fWIpsNQoWrJ4UkKbHpKlBuEWnJ6j4pK8AsFdIOnX5Q8seeGlwEEVPt9tpQzZ
O4EdoPgHe1pNiTBtzbWJp9XwPKojquxhGbj9U/aMx42wzBofgs0KXLL3Ir4q
RG/wwHiZd3d55My3op1e7rwZKTEcXXDlO5dUc0dEm+8qmI3CsQv8HVuzCdHB
0aOVcBODVYHUBoLm8fdSI3nG7hNtzk+Ww4xay3IbtWUjuAPC3j04Zfo7NM2L
BKS8vZZZ9MEtMU6KeE5igNRzNeesL1nhoDiwM5pFuU1X3oNPdFuBllBNdpAw
hEP5Sb7SrCZ1AkdH74JhEXjWx1gYhSBKG0OweQcVPAcufzQdhtnWZhI1j/qg
Cr0ZLIxDJpLCU7+B/+P6r9oGcwbm/lWaP/GxHCpzhPrX6BZl+pGaQ1a7z+fe
9miqvF5HREGlvHSa8IHskVNR9xEnBGTMqbxmy8KMKFLPr3sKeMNtFU27k3fg
UocNHH4a28oFXi3orRWYSfoEHhkp2/iNuHsP7Vi02S9IbpHs3CiJnwJgSVVj
eK+hgsaW+YpKMdYQlzQ4wh35nF99WLGSG4dxTCyOik7iS0OILJHXaU7vKI8J
NimO8lINJ59DPnwGk6uh1UpJzpOjRN7WmfFvQDT2Q35fo9kVYN94dl440QzV
LbDQFnKXeCJfrYT9ogf+Eg+VK2MMNcysCdN8x2sbaHKZISXbQbzm40besvYw
gEfsHHcra+xTtRHef7zOta2LcyGKktPfxi0rDhBLN7o61CHnIl0bN2d6ntVX
nVHmH6RFytG0Kcy07J09th77d56KUBWYlw7/BXzmejli86TDo1F+ktPMqFDY
qkmyH3BnIxre3CEDhk3/iG9Qx7bc3n6Mfmva+MKCeouTxymu1l+SKxWnjq+I
DSEk92J1ew/xCoQ3MdgOmBB0gbCAdakzeSOetA9wkHsE8Nm2sC2xIvJ0IMPZ
IoiJ/hiizQlm7zq1QSp/t97ugt/Y0XUEl1uJ6thAZMxX8eZRAjQ6vEUeRZFW
D85nfSniVG0OwCrKj+ptAIJWGmAGfC9VNFLCFHwrW9wTg9ox1DCpYJwT2yQN
CkKUkfCiNGhF/nhMxvWLMVuEVticzakBDjDKxH+ZVsacZN7NcEb6Ruvv9k3r
TDZiyRrmwzVBPklYMBkWrczh5pJURlzv6MtD/mQ0OdS1qW5ZCPj6HQMcMLAY
F+AsYdmE5PEr0PCl9mXA2aJJrNNSvojg7hxs7vzin0NDCEHqKntAlUUGiEaQ
7OijWoiWNJuBBArOObh8LHwbGfITDoVrAkhuo4Vmk4CCpZ8sAVbYKrTe1sun
vazgUjdRjcs60g2H0WDMiq7R0LS4Jwsv/YKZ17bgjS49VGQf3my7LzkpXgXK
ry6lX7pghduF+qBT6dC1hY34g2U1XPif66q7Z/F5LUNRp/gncrSLJrxm2nnv
ZnoN/rncTTgg25PdxJECpfSdcap6UM7RGDLLhLm5/4YYYIKp8n450RBKZCAB
u7ZQo9lpOz1newyYy17hz5UcpxV4crSMM/mTuaj1AARrLxkx6O+GLvFD5+4E
ebWcrThb51tqIw7QJnGpVW7CH0us1qzwSiR+LYwYeXkxQjLi/5SWtWonbXQP
RL0OuiMcBiVqLrGkA/aWAlJuoq7ddvCe3mrqJUGhpQLhO8tuDS8/jrKiSJyq
4Q/LI3OfqqIToo8S1uYo1Ga+lpRBwod13d5jB9oXcap9cWlZxJmPuyaiYdY+
vuOJW2N8bEokRdqscSO6CN39YdWaeSOUOsSTowbNzTlZfb+6Jb+eheLR8xSv
tkCOPGRO1fUqKnuY5LOZ+/4TMPNoPfmPlgaw3hSczyvw/OgduO6XLT244rre
j7S9aM7XTKQfZjvuDwSZDEfsnC/17otHfSgpPC2QLn3/qdhU1w0eMo2mCTfI
0r5tr7zPQVx3cyrvKo2GV6r3B+2ST0gw6IFOid6kW4mHxyvfSkpA3Ni07w58
wSAfyDWZGWWLZeqvLbeRikCjEqXE37H+wVbmtTegtmqXYsLOd87tdxPpSEPr
KSVRguGFs0kKadcNlPAqOKoNkBsEJ0ZZfWbWOnE+7POU8/8DtRISL8PjFPiy
D6p6Zmb+3STvpaqZcvthnEq+DpNiAPuzxCcPGHA7ww+d1sRqNFtZL4JWxjZZ
DkYVFVtvxXGO4CW53VGs2+5OtFgJjmVtqn4O9iDj3r+ol5i5zrKrwwbShtQC
vwSJEVq4y8/ew+tyF/BHMbuw2Zr3MSPwm0gRel5m0J7PKyPUBDwdnsMEPUCY
ZDk9CrdHHObioDOkYFS1KDSFYTweGH/LAz7rnY2AurojZMEIHBx09QzPV4Tv
IsTYIZyEX66FeQMWRbGQfO3ztmHfG4dJzHCA3aSLn8zN4INfMcRR/0NS0spu
UojULryl3fCKgh5CLNfFLzSesrdbujW7rQ8a5FECJkWGE3NxBf5090XlQ2e8
iEI43Ru8f3FbGYr0v+XeHH9os3Q9KVkXtgm0HccPm2iRMaUSgXDOfkgWfxyR
h9wFqr6Qb6UsThf4s//PoH41bOGIRHDQdxVrWQi6ppC1swr4JfVANZ1UyWn7
6YoqlNsuhk8XUnxCUaICo80wTyecpRQfJLbcQ10f1dVXtUDchZNJUUU5i1it
AzdkTrw7q7KNn3WwIbAhqyB0kUNu8wbe+hZnXVVJZi90GJNesoQvMV2f4uqK
wh4JR4TRPf4R0PHkWwGdO0Nf5kBWY/pm6EvS3k/cDLHiRovYtUqWhYwyZhVa
QURpBhUutQt0e0FC46cw2S/9P4eSUIr99gmjhem9HfikaoAFwR2ASYTbo9s8
LDvJLx37EnB/Yk7fFErA3Vs+fSKu/wflPQ5/zquwWBqrUsNCAW1buthjkEWq
pPc6eFX6Df8jUYHmE7YbfeF2htrtfUjmk/8okpA8VA+gIx86ACYBWb7DAuoT
VX9w3Nua3Z8lC/MR3c9B+l/LIJfPT0ITRxSV1JWKEJeTWoYRUeABabojDRau
/iEzvrC+5cr+fqbIHIrdXZwpCSORc7BsfdCI8a4tmRwntDBV65BaE9zThd6K
4OOfqb40HmzwFvXOnNwjsZxIk2NG8ETUyZdRowE3SOyn/7BHubyC+0CDyRah
RniZgSB+8GZgnJv+FEFYbcFxv/2K+dZ5owNg4fX8zqak+LgDfnkpTHiEZyX/
0t6ZzN97tDc/X7E/Q88I6qEyJOoxCS4iF7+SEIpoH+M7488Jvwx6H3PXdkHD
69wBG7U0x1j9II6kXgP6i0c1LTrpkxbC7yGjrpWutgb+TzypgQqWYd0umzii
qNdhY2mrNZRRWXE/EXPHaYOBWTn0x+QNtPLapaAX0IRbSugWkC4Hs7fvh7Mt
nGh8IXxXfCF0QZjh7hqhUasnPhU8gSjXIzmtxIczyonVdRdy0bsbQHkMy6BV
D77gv+r8amI0pEt2Wbv0Q3bMJ8LFQj4rhDGYl5g5NKLUb/hynyiQjMjLAjO9
66c+LhUT0PH10b7B0AKoQeUQxLz/DRxRJRe9Gvyu0MP0oP7Z+mAQrfjNu3IZ
FPvvlYrFVomUzpOCFRJpEoEnAx3kv/WhsdTBFZ0t3QFtLGOWNIro+V04fEs0
q0jk2VQl0ZsBYx5TEu8BeNUOj0drZFnwNz7X2/2Y+coAjN4Dm9keCOoIXkx2
mg1JJ+iQ5u+ZBGftzWSt8vOVZrFRY57zRPBdYLFK61b4YQox9FZexGJishI9
ljVVHsBWODWmDHq5iz76GBFvRGG2mXCJ5sA3kiOLVlzC77pSXzojDKzsMu27
StuTc+QoDZ8JT+9eWfp8ega66ryJlQuDHtlpHuIqswbfdlRXRgkv88aZAjV7
x/m+j7npazgCmoIfQAldwW4JL+FxE3LuprAkTQWlxSLC8p9YQawSUUAKhwk6
kiGuZo6Js5qQs08GDVUaBrLj8ANeMJ1z69zA3pKQkVpL4eOM7riWYCrbwqHF
/u2vXxA5no5+OrPsgxgVigyK96diVQ9fyOvS0AfN7IdpQ25fYmy/qOGEAMlJ
9lyXt/IG6+6+4nF/2Q/VWj70k6bK4fVBvsgp6ffrFOWQTphBpo4SZU6DRsJb
b7Ke3zxlWILKMC3tPhBYOnhYyDJd2xkxGybAuqUNb+zlKxrZNFImU3ZE/t85
KKjp+J+ZXJ5FJIRrl77tEVHdMq0GrPpUJxMvmBfZmwjBJByK12FbqZXdYk52
fkmU2mJ8ODW9POW9aJ0uZ+8iuSQOxuT+cGO02yFhABFEHRMG+08V1IaMbcQR
TplJH6g4UrqVWTb0c0H7LFDIFDTVCYwqRNC/P0O/bywMZHHapp3i/bJuxwkt
tWkem1wMMxtx/MgRIyc7GocNuqUb8Xm0wTn/fcR7V6gcIxM5nvBkFHXLhbul
q7aKHwdmzIRjddyUFjv5cqpgOpQYaysIvXXl1egYot6u2PY0sNrggLE9mBjf
jNB8/Bt+pbAU3m4/FGrdH0rAy/1Ogi281mxPUAozX0OiushD09JtqPFuuebS
or++Z97c7KklA7shVzQnvYTPHmfEI0XtMb2ELit4F6bFmHj4/fFwvc60gan9
wYlBFHprlo/qs05NBZGo6cRmCplm9Bq0+tjsksUmxuGUdWXuK1F7t+aMHflJ
Xo49xU+CysHO3/7I1dyaTPeTLveWu8KfKZVsceFV6zR2WN84lxPaekx+uGNd
cMSDkcRX+oq+9dMHV8uEdDYjbyI7eA84A0xMeXRFIHbWyG8TQjr/5RAy+YUw
uyQfa+RjOU4Lj/kznrrJXWzNL5GDM4nbrwFsZtrR/hoD5KK9IULCIlYbAC48
+laK1Gh8HBReS3J4TKxfM6IGsATXeWlLf3k/vWsfsGTM3156aCNYicZf1SCs
sKhh4lWTvknH15pXbZ1JQQvuCJNQSFQK9iQ1BXEAgxaEv2vgOclAWK4cjrtA
Vu9zpT4JthAvesRxNAVS2GkUcYH5LS0aqToLwLYXthaW8QA1omyvKJnhOB5c
K+ko6xjkhnVFMXv/qbOHn1m7+mYEIQ88thlJnknmpi+tlELIxbt2eEaYhhQ7
ak+pYhuGReXZemkWQ5GSAeFblofo0+OomBwAl8aqiwb80hk0f8Ep2/LVspIp
aZD4tpK8lsilpp3A4AGN1p1gSiKyTpBwoh/rm6GnQrWr17uTpDvogvffzG1j
nC7wz/6dYKLxXvlExEg8kknzl9Z5PlR+H/u3NmkCZqgE4ndOMw+WLB6TG46m
zDIV1o7tYawqsLsF6NYxqtMzZ3PARbX9uEv2loxEEEHVepfMhxZ2RfBZsfud
nua97zaknm6U2Y6EqZ3fB+PgsygoZfwSSQOkypayY2+UH5XIpxBg20/WBj8H
n4cWTxe7Z+PrX5lo6vVb/+bUrqABF7Yv8n6kNVYjFqFwU2Tzoh54363U7j8a
e4vFPKvVQeBwwtJmIl+9T+CoOhPdpw8A6LpxjlWrc608PD++0cbOSWUDPG/u
PPuKS2/3KkArauppDQONHdT4selpRfXEPi5g9SDrdSq0PG4lqr+bBAgXNAWj
P3U/iBdN5POGhGQwhveWzF4D/sQdbivKaqlTA2If06DS+p3cl4t3/BYc0v86
vArKUP9z1NRpYezmAoRHzZFLccofXvQYQH6ZPNupsBN59iC6hjepag0Bdd3A
mNIELuv0IkPhW0S7KPUgFZYq2yQ3DZ0b4HRQm3DhzDGjgz8IdIyfG4djwm9R
dAu6JGKbYNwAl4+bbhrjNNM3m5bKUD1w/LxBEStFT/Bw0NTYl8Ezd0nvTOxN
8l7S2e28W6PX2bpzDE31mPvIeEFLvhiu+xS3afcC2nON6T1kp1nHlIGgVU9a
SrHKxqXxy64HRYd0HVPjWcDrlZfe2/7MlwfY7nq4gf2V85xTZ6yPt18DoqrH
CcbfAju7XZXuZkXl+rs3+JsR8Z4pUcF2kL6NFZneRsCGiTpuEzbjobHtGe50
YtVIUt+510Jeu1brWYxWEB56gInhDwqzvQcWJ6lE5xTo+nafIg2baJKPWZ1h
W14kakk8u4AAj4Kcju1UjwASzqENrDHd2RPVXHjlHltMIRGCPbZ7zytDoS/t
lyE2mNwiSsyYgJy4xK17Qxfb/7PT044VtPY1WZuAE8aVtrP9C+Evssky2ndh
dkC1FX86/tELFZhxGM8MpjXvGB77WkdXUX1ZUcmhwcQ4LvurtqIp2wNlHlov
S1bZsQnrKVOvQfBD0uoSZfyMqXEnIge9I9fVmOMOgYiw97RLHMZ58ACUE23J
T+mVKi988X4zxI2o1zITGt1VzqOP45n24WOT/WPEJWUAl0hidj5oU4zOGTTr
emUqf2bjHQHOVHRVjTiLXttHL5UT3LaTcA78tBfu7IoiG+s+lWzIPjLjjdHl
0OjQaaBs5YGFNGIYiIgAP/0xsMHEJxtCzk5HYV+awUNLacY587/wmaoTXusD
NWLx3psxX0fcWJTkC6Y4wcmaKXrL3VOMiEzkiiCxa+plNZIWemdXdR+CEx/O
apngiT8PyEWN3Oh2C9lq/5fdT+iAE5aHEbt9soJtXvj1gdqGqNysEovJ1QsJ
1T9fwv0O0A4A3E10V3gXfN1pUweT01n6KycVuOe6FXQ0xIdKseMBsbyvSZ/g
LarshwAsvQbwMGb5nwHzizaePbKuTtfGs/1pdlMcbmnHmDYuCUOaRakS4xWQ
oFwbgjBBLkfytrha7kSCvCf9649wPT3Vilm4tFoP1gHCgXDNeYNdhylrqa+8
HPczWyqdIiDzUX0c839fZL18pjMjSu+CLwCh7EXmLdjBnwqbw/g9kZNPc6ir
V1955z2KKI8sopBW+rks+C23bhtq8/oG1gDCDVcIcV+ew4phugqdcRPjuS/I
2cxA6c/GNU0A3lFMPCdi54jTQ8uWn8iNSX9bRMxg5ouREVeXPkazqjrxAw4T
cG1SJvogkI+/viZG5zgcxk/LBVZIQaF3QVM3J15M+bAS7OI/eTcGg0GNyIO8
UkEpvXaY1yDUIT8ix4YFaNvft6p6RufTLmeCIiZourBOlS+3nEIgN4RTxsjg
m55V1J8HJNIPWw7of0xLMh1PGN4XHC29cgqC5tTDQjLOS7AF6NZFUT1W+8fy
fibeRwtJuRFMS+aeO6waGUeut94CukzjhNSXQWck4nN1Dr90RbJ3JRV1ItdJ
MtoZDJ8vP/k8ngoE6FOJBTHdrG/zDQda9bHZhv31EQsfdQHtKiQw0oqkPprb
kuS5h/wOWnqY/9TX22BRmBaQs1U8cRvRMrokgQkS7ecSfe/RFSKlpP+PKoxr
jH1Ut8Zwz1BNEvyFCLUCzDVSQfrfUdhYWwSeHRrAEwz245RRtG1qpHtLZ2jh
YX8ceHmuTDO7iShqmtL2k/2OrEUXAguLEB6351zu0w/GNvaRC0zzlU9xAypH
wypordQ92C0xhq3xs2hOcmQvTEvHesOquQju1JjIS1FJVdrTMeM+ruPwIkfO
624zGrEFG9qOoBl10B+WuuBxFIQREPjH2JfGOZBqgYVlfxTrZ3ZwCeZ9scIZ
7dGxwXypgJkTYT/SFHbMJYfqrjipm6nFM5tYqbpNYa0Bc4ekQHA7Sj9B3XGc
fU5d5xONbxdDAwwNeIzFQ1GUy7aVPGX4rUx6QKA9vI1MsvEd3z+s5S6AhDOr
jnKdtrjZEpOPw4oZrfO3wugm8bXa0sFXAuRovu0ucW7rwjoQMwWjh9edwXV6
HHy9udYO7eN0YJgrNQOnpW0a0gJ1GdnlaRnbs3QGsrG4MrUpRdRneI0h6D2o
hmz4H5FTzQY8vKk0M/9KScuYSy5eNd8MuGDD3S1mrqKx2LRaO4sNKbANXJxw
zBlPXL8Xvo8/pJ9gh1AzAa3eSGILk3d/AUh7nIJkMx4TlK8pjaEu9/jZ+h1Y
LuQdopLvOjahOdREuxsPXpZER8wgsqnG9tsZLxw100EkzXyAC3pIcm1DSDKQ
vYuAuqip/RXRBK6aV8TBjFuzw2RtJVnBZj2AffyoI+JRhdB1LNdmfLeq7pkS
l/OWhTSdkPoifdlc/tB52z+oUOSBOpdmcWBVoEoT68WVT8dXZ+pFNjFsZvBK
xU+dyqO4Qf1g/sLW8BqvttDXb+84ZMbah50sMZLTeU/AUhF97aRmho/M7dll
WxB3SpWMNRijh7OvtR3pOoOPDAFZMAew4mCOkGWyorWKGF/J8VOXZu5sOteh
+GJoTzNyTjb2eGTh0IwyAGGO2op0CNhXPwCL2s07WminW4cqxkFqaVvxXbmw
DYVAIZtWVftn8N2Z5R2UsiUe8ZHuNPsHTWsDbX+d9I0J9FJXmHgbsqsgx0nm
W4amZGbB4hLOXYs1SuJVLBuooXWsUNby/CK4Z7XZmFIySS3RVF0BFHEk4ICs
o7bKNaiywjqiaHctGMI8jNoc1MZsdRvODcL7zLs2iyeSuJjZ+7kmlfGknaS+
+Ja7jKa//Hpoo5J4zjiG6S2TLKBHIVcdlsyRSwEFYQjm1flDeO0xJSxgs+zy
Rk2+2auLz04aBlQ36crsSt5fjJgpO8z8Hp67/GrFhZP70bzzZ9gxM/QGuLq5
6OvT6qkNhalDk/REM5NrfWzjG5CiJVxWOPXMMG93DiSfalk1A0y4/yY+9w40
V3UGS/6aaiYVJtzMFG+oLBHkfCWBxlZUhzFfyRWaKhf9yw3DntL54cd2wsGA
y27oqbm84F9Ii1jgtnWtEKsFlBLHddPdO0uL5E2TS47FaMnNi2MkInVhQyB1
36ADyyCoFitnmb/3DsXLvHSiDKMGzXvGhgTSA/P+ILptcu362uONgkKhUaim
0NlUGwq7GmA/1bj2X4RVpNFYBnxYRdIry6yFLFPOn00fl/umxErKICSoOdNZ
R56TScEoDnr36bGppx8D/TrvT6wkRB0jbLUdxZhXVITjYzdCvG5GF7pXa4GD
oipijYNTy2RvWGwGOMgeWeC4wziSF5fcEmLjRT16Eq0I4MheSA4puZsnAB0M
B8uYLloKxKC1a2SPv5c5NPPWh6hqTIgmklNpLU1IZwfbdSMJ3vkVORXpctrR
Iewifn06AGZtuNce/+EqDwUJ5JEW4DcScEUoMC3Ia+jBjTb0PTosdsUkgokF
JXeiohYQpJPqziDOM9Z0p0OtMAU1QYLoeP9iRxkIxqJmr89UvaHcwNM6GZo+
bvFdqcTbZZ0jsdFkCcxUKM/kh7fMM0IYRWn0ToJrrYKg8zATOBLiWPfZ2a7P
5SnrWJuZkAERgB5CGrBDwv/F/zsscGTromPKI4EQO4B2Vr4ex/oNdGVZ1Ju2
yaiwTEBnWMjCsNkl6Um0S/N6oprNQO10cQv9ZAWTaxCk7GtPSjXZo6fiR1fa
EjiNl8P0eXN0ZUkXtSvx1yA/MxoizYUC9cI3shs+gSY02+g0oOZV0yX0IRTt
LPp8/am8XUxsZabz7Q5efnnEdN4lGERq3fZRWlsf9A+sRtJVwGl+ru/IiYQM
CHmjpu5evpCYshx7XbyROFsSzhoQkJhYWPqyzGN9g+eXgJIAkNVGnrbupsBA
p4zCvASin+IV8CX3tk6BZEvwsoWY9LBM1R11Gin4lsg86hGpTq6gAJwkN7vQ
RzVlKh1lxVz9B+BmjVPaaI6Dd8LToykQc9reBdQO2yuH9BFABCjq0TpK6TMj
WhzO/sLMPSalcxLdNHgBrx7mM5Bko6PXHQOjPSfAWuBSE8V5S8ac/QfJClN0
gRH/B+Kc9qbDmyiJNWd9aEP9mPl4orhU4elTasjEGcNUnKZOn8RGYpuewFUH
5dAtdtQC0F6S/EgpveQoJhOMhnaMeJiuo/WrnpBvljZsxwirwFIfNTIA0Sah
FmPx7uzVGTZyq+nQO/VNz4ZcQgQ3P5gjv0uu+wkJQpBNqwPyjcQiWJ6MR/OJ
B4dcH2Z51VAJiIpsJEK5o9kFsfqMHmv+N1j0rBtTPQZh45emLrStIKOSSvDI
5deghWdCiIV2TteIR/dzcDZ4lalLG7/Lp4rnSNR61Erjhnwjh8WiXNwGTJpH
2YScS9HWmIBElzjYTkVZsHMnIdEJKeMfim1Y9GOwTr058McwtrhSEH3EycVJ
KPDkTIxlcEpf+ASeOzq6iJFxNYFGP3z+1mMClm++JwRdgQOjJikfmE4kr7pc
2cgZ56IfC5VjP95qchfhaEcToxCxhnHt9e5oNH7gHEOOD6ryDZ4SScrHklgk
Af87d8d9lVI0REbJy4ixuCvVqamhQaymeV8AFTH0WI8rQguQiWd8Hyw0bEi+
1WDM3tm2XJWvXHBNFiH8TfVVsGeaz3J4YnawPOZbLAW5Q6o9nhLCkq2b48n7
3lYx4TqeiHfzTt2+uDvaBKK4rBFHblfhZDxy8iRIKiuO+AHuIuL3HXlEQidH
4sEkttOsaJ4xbj0GuJl0G8gdnxKEvEj0VExnCTTTNeM9RJQX2cSbxYnol9qd
Wu9m1WCysyz80hNyj3p5Bt2Cez4wEnl52G4pH/kdxpL8T8/fiQo0rMr8FtnM
XF2Rikp9Ow57T0opaVrZC10Kwd69Nry6vG6UqtpC9EzUVaLf30f0GBbvIHc/
Sx8MQrJGT8y30A9hz619sx2HfJ6Vd2pZeSgZvnXQY4m5q8rZsUizmByosqT1
USv4Rzag3fPwUg9YjvEhq2vC7ryyvxSx3nwm3OSdJgLOUm/qvq4xJ9p6+TTV
1B0neqIJOxe44y89QmTQtOGP5xi/23s5D/Xnu5oJHZhSynHYkFw+GTcBSiSD
kb/5muRUtqkAuILXj3wdNEbpr4ACV/dWuz6k+atyaBMXK3U9+qQvqSDIN1kZ
37MjabnbupJE4ejCeLxTgJhCq+SsZovFltmlkwxjMaaoauxF8ESPyAtsSuaK
im6Vm8Wtba7vL57vtVm53X4tJa9/cvCsA3AwbN7cNShCjuK0AVkZGsXy6KYR
XwWBm8RjxGZgpxi14c9jx5AGXyqT+AGph5MLtXbr6bEo3nLJGbXz/272Igpx
s45A+92YdT58/2WhvqwDwUfLmR5vhD6a+o2j/bPTvAuwu9pwOEynYC54i1cv
n7/8JQYce5vckDQVKrd3vZkOIspUj13ShglQnoH9B+zGMikCPwyzydV05St9
1rsXcYEH9240bALSvJflOnaBZdoVJYnjYGieKZpUTTJJk7CYQP1UdXcOPHbn
avWC4qkEjaqlIt5C+9SRBuLPQwVISbk9ee5QwQafh5ZMCv9owMHNSx2p2Ztl
HTA+wCibBquxKmT2vgBatKqqNiHCbiqXFJH2GEryvMR3nPHqWkPr76Vc/P3S
AUmZGw1+9f05JkcVcKBJCMcZeAV5E3MfmR5KMvKK6FlKGdrmzdRhUwXX0JUJ
KhmDi4L50uJR9HisKcpc9rvIgXLH2MyXm5jBxNFo0zWXLWzODnNmIR7JbsDs
Gzdg5pmG2mkRwZHoVOhFsjq2dNAN+1ohERAWB8frnYu8Qunwwrfh72TbqLcG
goAOceCGGbn30R032xYQqEOP1hY4KdsYR3bhb/a2yCMBYLhPIxx/yfpfXo5L
YC8npJHwv0DevKk0BJVyBiwPVcbi8PRZKmWrsb5qppU88qrTkQ6TqKTWqtuz
Wg5/UWOMNRrk6uFBsQnM6P1lrjJRJQhhPIqDSCZB3Ta17+JcVu2daRB4oFZJ
QYT8WcEIzL72mQInwuGLGZE1ud0pZKU8VVxZgsy6XqlrdjHZVFtDtIX97kwD
Ddm5G0b4okliNX2xAYpp+F1ryjsi3DI9FDcm3YfmYCtQVFC6pQWpaYfs7X58
pDWGrWk/DS/hybVT3mUuWOq9Axftt7M1VENo9rrVpdbqoR889ICFbAmBWNYO
egipfqQz+HfBB+I161VFvI9Hs+Du70s4rELQETYAhGkN/SQkwYqHyo/lke+k
3R+ZvMEcWAGoUE+FF6UxBry5Uv6T/3A2oqevIgXbJ1T538+3CdqRx/yPKipX
V/lQZeQvkJuqX2MdmzqeBL/kT77IFjPuV4728rpatf4VpBf7D5Kaqi5EfRRF
YyB7IEnbO4oF8qcGNmGuEokAqnPgCrGeb0l7Xk7gjI/yWw3SeLIs0U53TEd+
jDaSMRg6XbIBkCTCHpqDMB4ycfETA7W5EL2afCQhFfErMIt6ADfoRXiN+/V8
S5Qd7CmRNiutreqwN1OFdiE+hwh8act1oz1kItHrBCpsp2q9ixoGFzMwrDvs
YDMH547F5/o5fAlssHAcgUu9h1zzzyMUIGzTNHL3XnKDnll6Fz63q7ASPU3K
GLFw/UWeWkRlhWm9gnUd2EqXUY9+fBsi2TNRPiBWNQhTSFVkrLzTmD6hB4ef
o1HMg7/k8DfCVwvU/X33zxtLNVANjeBPqNbUzVR6ltUocBMmL3dpqyNnYaeH
FdZ87dUyWqlVlNeH8ePjsinGlQKnT5EUxVr1P4q7gqMnaa4W35KFxw6C5Mpe
y8eFL3NurhAVaS0fRQpyMtyHFre3xOl161yh9qLt7sTgxW5ZwezRv6MThqVI
4zb5dlAf4Pp9FfV84U0HoawuAd0+fshuCecKnB+XTYqIoJ6zSrAKHPCjFHki
Xgqw/myxDhyCtQbhb/BVe6ljeM7FrZ4z/0nrRen6L58lhiXHT80wEd7p4IVJ
U5EDVlAS7AEFH/oWgxM1MHwAecrBtubbrhGDEh5/rbDMcwXsS0UxxR12cg7x
rJxM0dEhL0PsfwM7r/Bx8fB/VpHpYOHO6GMIJfguHky7yar/wy2tDp+XnK77
fKR7HnqfK1uJf0WqODmAjmYg8ytv/alihEw2QpSwEAsDvMq5cPBZsfohmqXj
0pUOqQUXpk1aYMqJOJxeN6u52/U34ftj0CEPCaKUfkhPAOre1p9ZH+6bjJfS
CCdMuclTaHOIGdQ2piA/V+dPPj3p7DDqvzjry7eCe8i1IdZWzfFoOQt26xkF
NCfTfkUmhifklyegAQoTi3csO8VrFgvHfd/JMQ2CuJ/VJ2xxTj2zZ5VExpbR
4BNQaOTLBpw9woZcA0s1X/WGrXKIgb5crBUXCmbFvM+uevVRPMfhhk7xMT/b
i5jiPHHKrQdx68NCyzE1EzVPDT7ea1ZR38HsiiII/Dv01/yySqYUNzzCqW3A
NgnORoVdxIxbLO/mI0Fs5IzwUUQ1oLrvhOBWdGhpE3iPK8ls647yi+kG3lhL
87GxgONJFkoGatx05ntRpc0QMxJT3KAHLD8Pf4manW8/kAyZmokUY9IIjU6d
Tsr6S3lBw4hw+04RIoPDRYegjbkMuZgvkDfjK/x1IyO0Btb8wPOcLuEq5URO
sFkGCIRt50tHoHrmwMWNmbFGg5h2TNdvw+aeOcU/9MNQthFzr87QtKOi5gP4
ODWWJTAWdOpAyRr618ic8KT0ocoqfX0dytwMnPMm+kNtvT8UTRhYksdlF1AY
6x1S5I+p10q7yz/BaWBIEh9K048ej8l9IqVdfFiFd5780JekPZv5chN7dQZa
qek65rwBzzb9AG+vld2pUDE8ZRIberIx5QgsOQbSaHfsINthfpEH1Qix2GC0
Gqncx4immF0XM3UIlMKs+PRn4AW9M3FWuWk624pk4cEMA3TSzQF+jq6e7bgE
7w7JkLcg3ScAK5W/guD1QvDL1PjCy0kXBGX8vIvBfUqSyM5494PLgn4g37F8
/6KaNvV0yZrkkHKQV7eyVQ5YnDTOfVhibWB6nPW2A9NuDuF1gQjqgDSJhIhV
9BezC0Gb3XB/Z8NBSAtlLVfxN1/eCVWrOFT6keBfclLoEzn+l5lHUeRQpr/q
/zBchtCWVuUx1f5GtdPS57EuxHWmdLCUq4hVixxcrbwuBQG9ytYl+gV8zOf+
yRsw5XDguhH2gs1Zf9beoYcLkWQ0fTPQFJd5F3yNiqYlFCEY13NS9IW5VWx/
WfgF9V6+vg+oHy1A6kjKOMjmQOHoF62Pg9BKZs2KYgYukX8hLKNgOWu9bWxf
NWgSqG0BXov3FSarCynQEA17SzTJ5uQpgG8m7J0BDi7J4/GIJNx8GJqDojR3
kbSW9Ngwg4BmB3l32lLiDN1CD0KpLQs/1Coye7m1B78shwtlXHZMOoB9jG4V
ICM5iaFdYYIkaUm5SpG+WuDS0DPl25xQF6CgKd0epR1cfmNzO4nHH76Zg2j+
TJnZeo02EKQl1lfauOY8oN56nfs53mhGWG7u+eeGqSuA9Tx1fT4BsT92f16b
qPTD2aIAahpdNuXwtvquwooC3QRQdqwehhsTUWllHOvwyfTW+/9It2hEzje8
EQssd1XdwK+GJy7EV2lf7tCg9L+U7Zspo/gaQUyRnmDh6Nm/ln8qSQbwBOYG
xblMa5ND66yJnhMPE1qDrRTbT/xNDrEltfVHxsnzkTwjkExyn/xrcfmERS3d
Cr/5oxv5AvQTTYT3+EPo0TG34igFUyErjP+ll9ddqOr9AMDbEzSbu9fZ5LmB
QjsFnbnZO91dytt+zHIwqocJpu8RbQQ5AcyXT9Ich80q21DgA4K6LjzbGBs1
I7uOUO+6zLA506wfPZp1KoH9VLNpvCEfCdhEwZZZ82zftXiyVhOZevyyKH4b
UQkXYwX0NEG9gf29UkP1Zhx41PuI0BsSa8MZsqoy3umwnHJrtGtqoowCRr8W
M49Dp/bqhShvdm/s1kwWhsR5ot/gKAHKbI8QYxQNXpXkCCZm8iy2AZV26kH7
EXTorOvtDzQqxs35t7BdZf5/TxeD6P86th8yYvnjIgK+mYp5wFcGfbc1LILX
klMcZso9jkBrTmh3udHyyrqFYCaUQfD0BD2ovcX2AnCh04kCm6aaF7gYLIdC
0Nl3EMkptPH0FnDr47UyjYcXcdspY6sRwHgC9RG8m8A2CA6nTxdmFX1r7PF3
D+Evx2Hc/PlwoAufrYqfIK/WJlFM071z1jKBFNtX2r89wPjJ7L/F33Tjwi4Z
kJAAFuANOV30EbzVUridHl21Dn1dHIp5ecLnN1LGqLHJ3qgfdQajgBK8FGte
7SAyUtg9IEEHMX8evbpfhtShPBVyT+MiOXOaColZymGBNtwhQeg8pfly48y+
CkdwxofYHtScgS0nMybHJXNUeBRLrq+Wb5PMWGQ71OGKZIi4DyztL6Q21AQ+
vUMoS96/eWPsFLbOHlNmwaZmnYcKXSIeGltLtiz606sMGFLO47dXGuPQzodV
1MbBoTQQlmlYvy1jJt44pZ3QHlnjLji0yqjP4K6Xl2tAXpewjiughi+7hl6Z
0iA0TJ409UHQ/33HHMz0Dk6PAE3XNxcek4WmXakNaKknrZDwdepbDq8fG5ss
k2hn5pfuJVW63aARRJ2AkNQ+lv9Y1ilyNv2I7j3HOkD5Hrox5wyXWf8NQd1M
GnzKfW8RdE6mHdvd8S4/ghoUmbjma5kVRfGsX41TWQvjvdDaOmVFNguRdiz+
sT04yv4GvOdYMUlrVWqF1xPYSPIkFw8G7sFhJUwhf8KodcZipeI1iZzcAiqk
47vegDbCRK0l0WhaTtULzwzSIVfkWhpHyZLqXxxQQGbpQEEUiFFLSo/xCM4O
YzkuJdP3UeL9Jzi+G40DABVdPeFDwUZ4PjwkBCLYeIrrJKdEb5117pI4ZfCA
C0JrZqlCAHii0ogy64Wms/UL6UU9rliKnqJqZoAdgp+xbMtSIRQzE07Yjd9X
fkGuZmACtLxiDVK+1dkJqm+9WGLb7IaeUwRMv4ikmFGmoOZS8tXwsQXSMGZT
Rd90r0PilaVPtkvrTr4UJDMt4ssshAHxfp4VNGCu6nvGn95tBUynCKRLk3zQ
nBWL1PTSxVcpoDQeoQsIWJRnpyrqMtPyBERlVF2m2DReR0ESLxskQy09p/4o
/5++K76lQEIas46+8Cn04jrk9MYZq3U+URwu4tRkI5pRHcym6V2W563i2Flm
c4D26Tl8CBZFzpKyQC5OK9YE0a5TEG1hGL2ZvBdDTxX4RGjfWLT7lmBbrzZy
nT8AawWrMU0m50P1NHJYmVomo2Kw3mARS8gkI8j1GxXUBeorb17jkNz38FDM
JBBi36MkjrziBcxvUJZa8eK1oQO0/K7yOiR8Lfghax+N6Yob+fIMzwfTkEC5
q4jKKkoNR97hH6Z6v41Gq6k/cddhIInk7MqdDfCi92P0b142HV6QEQfrRrcU
FoGQzK4LsjQu9jM/R3YFMyJQAzjjBPxrk2G5DbycSoqfdMpIaaiRPR8O5CHv
Ahtj74j7Fw7eKHWhktGzLnPMcD5dp/ivtpAF2YrJWbRxwNjKSsUjuTRJdWw6
WZc++BPWMkILmv5gt25hKw/Aj4ldV0emkGXokLBVWXO2MWW8q7bknUiqloGl
XO7hk88bgGZy03aAbav9ew8BCrp6/kflPxhqMrLlZy4TQ0CyrXjenLsjE97K
Jp0lZCyGcXX95JK3rLNqKljRj2CQOoU9fwlfNy9psBOPR0fwsc7oHum346ez
1t5z9z7aFhtBLvGdqsPP4k1txYd16e2+6KGeEsoMi8yyCr0nMCX4QftZBBkm
6pEDsMd0pyg6Xx8XjneB6dlRq6m5O+ZNzFe+998S/YCvg1n2rB2tzBnNJxJP
LRuRft9bo4FTc4tsJe9euyxT6ZO7vTP+fMU5neTsZZyx/7hIkCnpv4ULN/4Z
ITnhmC2VFbSzAUzZC5czBH9e40/gGQu0G0KuJ5bjlHjWXVx3SIcVeD53PM9a
njkS+/sK7m1QbczvZccwKNpZwrf54V4jMzr5P8aQguDzWsdZ6yzPScjYOyXk
2aUUjFEixspsz5c6WWf+6V1IMOUMb9WTzxgN4mBWggdedQM2ExRubiNn0lbE
2BYzQFeo9Lnuzhqewzxyn2e1Fv19nngUvlCQDIedOx1Yr08CpRU5muBMvWEt
bbogaEIQqJxQXaOcxbtnpLq5OLwDFpaaaYoVpsjdPySlAwyfi4pnXtXt182M
8bg1Xuz1dldKcoFvsX7tc38dJ3qtGpM3Pd8xZJJjuyx07AgpU53EPQgT8JuH
UUCWIZZBtUJNoLWqfQP3/zCIdlHXIodcRSkWbQE7xeTVFCJlYVTzvlwFpS73
TQKYKkxcCNqqnj5kzEhsuK5rG8DeMKJ3DA+5jhYo923c3XZqHnIC62kYIjel
/2xFseMcCQaKZm8Xd8GZk4PiFtSobJqSmFVI3yxZPij5q47dMXL56qe4s13M
CA38TxKRSb8rtX+/33s248x8OWCmiXXketQ0zu90UZ2puM3MOWn+y7ND3Nq7
Y8g6zkYGMFgEN0LwwNm/csWQp18xlqhHvwstVu/4Av3AQA24M4E2tS4Ly/a7
zt77ieLVuZ310A7t84DrngtlnzJQ5B5ylmaZU8lxJAmwxZXpFsAREn6a2umN
itv+HSJC1L4P8GW/og5RNZfuuGwSPGa2vai0gdxrMuUlXEA3EXtp0PqzYi/q
dtKqNHCZSfO7D9+1dah6kz+KYZcRMGDQTLR2sW36NZKZ7+pOOtzaKIARX+60
w67tvD9d51GN3NiyHmRKFHn8+exZbxblXKQgOuut5FfrpxmDR88u6gJvhF/c
5F9wzluES8o3NS7J0Z8klH0YLnH7V3dMV3xPRGj+nQyzdQuNdZQohpyEhRG1
VtIt6svkVIo/6cT9K+3U48AWNTOHQlcQocAmsLReBIVeDLTEsg8rT2CymnCw
f7npDWu2R2oc6BfT1iRlEZzQlFplOGNcwgFs8RfaQfswGElvumVCeU5al1sy
vrLKslwZaX/FNzkHaGjMn7VBoNVwJMRkDRoa1ZbTnAs1nsuQVkHFXmGUTubV
f6d132ImLq2Mi6VgjnLVj8pg3o47BtgdMasdPh6J2fJqfiw58vl+VAgD0hCT
FbDZ96sbQQcaSUestFsmPlnplVqZ/xYQmingGEFJ1+/ICcQa8g0HjZLls9c7
Ndq3F+LPizuHeUbk5ntZ608dPiKjzQmCguRSqJhsVXDcloFWgMyykQ9TKimE
rdFDzatT1zs3hJVQGfRstVQswq3DZXtO/3ejaIJdxFC2pyDd2SG6ypMBCfZo
d2xooc4cMt5nrur5jgfjQRNVvMn0YCXGsHWPZXoS2vWuvPeL8JZuX7UlQcgJ
hCL2pCAC0QOTlkddQ8YmOQI5aF5DseWV4XnMhUPV6N4dadY+IRTsx6PdyII6
eqeJO6UhMGd9szAZQUQtYfvZ4y/vB40kfhoduQ22jQNKGSCCx4ZEWZfyBja9
Fh2VsTRUyjW2LNitSics/oMpbx70U0TPTA9qxflntZaMF9pA80i4BGajP3KO
ZQpSJOQw9T/e9oLoZCXk6KSMvxQ1I5BkJdBY2SndYNFbR2j+1Gu5jofc6aYM
oT2pA/S3dJIsoFydMgjVk6Ylveoyiq1UMyoM8mHWZCjXwp1BYAMroOLZISJk
r/OdySv85XCvomZUHAzEEUn2iPQWvpxfvt1yzcTS9k6dBbNFgzVK6Th4mzr1
Z23W+RLShLA4C32t6ZSRoOkDbjJ2I4jNrr/OWIPaXeHtwq5VQdgUnqPx0GAO
sDl/MstoPZEeuO/GCJugQHLNB9nW3EZdElLO21BxWBkmzuHDPe09tcFxxz6y
7l+7Jo5PyC8ii+XxxA2aTfWtpEeefm7tNAl9rRhjCBOvOUxjcNXyVS4Vnr9T
JgABR5/TeGJ/HCo/xyFKbCPAlBnrjUGKWCGRbbYMxt7OCjpATNgAFabnkIA/
MWLLXN8LJk8SzuJwiul6lwf20TSg1bWlIw2XMRrojiX1loA/O/KpN+1Pvia/
Up3LgtOuhMEPbi6jmwoRVyqJzseGKMpU+JzrUKdIe3dqw97ZEtMLmR8Srb2m
X5078HnTlM1BYk3qVQC9foa6DN7zEg9EBN6dg5+bSfRSKUnkQs5eR8cjHkr3
dUSaQW1EKp4VTmO9Kt1jPmi57mP0hI7fd7bUugtQFHkH3Sq5HVagCEr9vKKf
69qJFK58ahePTezYxBkBmWtHnbrfIC5qNYbfBMXHIDmgF5+UnVEzHNnCajaP
5h3UZ0IHQIazfgJl8F66jZIfnS6AKSknnV5QozcZmVTFkAOFHv0l+UoK7Lb+
7PQTIWwUefcMoVjMMwAq6+33A2ZcI9E1SWYjMW3C8eKs4z/5QAfmfd6d6D7F
IZtSQr0VUrmfBJzyMbQtPp70JWtKqs5t97m0tUuFbEvNDngl+WLVEdBnKmni
EgvhvNe2zBXkV1T9R5ZXysK3A/3JvXbp9lFNhA5en8ciUWBHvu8tChzmayVl
ApS/HiD+hs+A03JONuJD/xZbQhCvlplKLQHUPCpQ3oSCIxz+vQNM/Clnm5uo
INtD3gleP/eelmQs8d/fA8VP5vTjzmz8KC4MPgCnWkC6PQmWzqctovm8GhiY
Vu6h6OTG+CmIEPgysH/d65XnDK1mIRM7IH9QsY0dxfjr2zRdiFTCmOf7jzlf
0BZFdKaRABe8/H00LqSQX8dDGfxM/3Xhy2PbMYe1f+hcPSgqRV/8xeoh9Ruu
6HzUdwdkGzmjDCfcO0rgUnbpIzSqmTK4yIhTqNr775bI1/w9cZM4mcapMn5k
f4Thr7NHesabe2APpw8BwdoXFfPZmeX28KYqgTkvqbz92+y0m+886R2XZztU
uCSw6aZDvyGZY6ton7/WAyBfLpvhzPvooB1M5MqoL6Cwkl3hQRez4NwxXtbZ
E7iz/38tqMbLiIdAgXMbKrmdV+ujbFoyvkt3TjjOyKkKPylVpKMFKSRQ7Nej
r31zfsQJ86XvND4ZQ0St6TBjIewz2csawzHqfHDJALb/UsHtqcCBLvn3zfxl
SbR3Izau+4d7xs8JospoHqoB53I33tUBReTWDMLpubfn0OJvcsoVlblAULj3
fqOYspn9SHT3olCpM06vexxi26N+OzQfLCDYwhjDkP11+dgC3/Qx6/hW3twi
5f6IOX5D5LyN7GjubQIQxs3Fem1RbGEC40XFQ2Zdjt0Mb3aMSxWHAmY7ZT+1
KeR4gLptgRTN5mpgIBY3vCrQs2qirHoEPkJ4344RZvx+KnwndztAnALGDjKQ
Aeed8ZSEZbs0AMn0TX8Ic2BWY/7uRFc7fpklGUmoYxxQ7OOegtK/5sJcI20X
I7mR15Ij2A5ryMpkIB6SffZGP7gEp/cFWvfEkVeQrjwgKMd0Dwin6jn7ZOet
M8oOJXIgfnnEm487RcSTZarjmGSBN5oyexUn/0i2jlfaFESe0djhslww5hsF
uHIU4nQXqH58hS20z7y/SFTiwVZSIVisFRgqiCE1MjiuvQjAlTjBhQc/wPjn
LJa0QVEjTzPEQsAd6Dg2Zt783VZYXJ1VLkW+Licm0DjUqr7zSW/AE0sLhaiP
2Pf4jP2QDE7RTPhQCPBQYouIl/LgXTg+w1Y/IwdGZ4IThHzh3A4+p/mCW8kV
R3cAxKpX28pC9T219XkBnMt15RivCO2r2grMjabVVhp5HAtOZI3YCAPqG01z
ih1kCBAE8XXm5+FkvE0Ijha1PkWChF9Qv0xByeTa6tAk4ov4Dp2oidOkT6tQ
rznxoI4qoXKyGVQJmCEV2EMAwH6ETkguVlWwJa7L0P6IfsmokiFmh2tyv4Zf
YNg/jnU4U9QjY8ZgEav4EmU4IYP8M2iepZiJGpOqgz4nDhq1wVRwU9hNFWje
2ioQkncnxf7Mu5q9Yzom/90XGZKI8AcsAnrh44U96N5UHXzDTgEKwadIaIie
uydHG0lZgin2JSsBwmNEc8RmyDYqtEtC1ygvY6fSIp1KRzsxrpsUE9LUa6JO
MuP2AnpUOIf08Uu5S7h8Cts6WXDSo10wC5IE2Vlq+FRC3j4KyMXXMeFRwtCb
OKm9abcXS9AERiFPH8x+fo8wOmCKrrffL3C2LdGeDCXo7rkXct0xPFAsUHOx
0OEBFWDQ3OGyR/6x03dA+DoJLEGw2qqPkz39+HSWDBWrM5sLRZJueMzA335R
oYKHesF58PCDYai7vGNKvsScZxpA/fmmkDxPX0eixD10jvwpAhbjxVhaGwFf
xosemz+SIamU2rgFbiWmTfoCdv7iHi9TWT0J3HjIM8bmNrMSQOoBREZxZJj3
s81SLt6nt64y3FMre6aDsGbnHPPh4tCV1BHNPjwrtzQlpnbX3lpqDTJtklri
qBNrTcTMlE7HhdwiV4l/sWfItIVxkt+p97KrrVkgXmBSfT5zyhGXG/0WpPT7
3PhA3sdaZjxkV3VGA7yI18LUDUQnqUepvQGiyIewuHg0Mq28UtXSFGLyho6I
ChcQj84fa2IWq3YjwYLl7wknR+UlDf439no7gIzBp1NyyspTO66A9zRreVW1
0MYWXCXck+hApwmMqVXMh/adImQJZlWr5ds18jyS6M9Gho1L1m2M9UYSpFFh
5ZUr71ZuIyRAr91OD/CKbJCtCHtjPhpkiZbZLR39IwmS0M7ePr38MgcNa64s
YAqar9yQSUg2+IWMu2jXd4TQEmeWs0JW6yfa0jPecuY5KmXNqfsIrSm2p2G8
N11goy33Lu04bW66N4EEdK430hHGpjmtR4C2nxfuI1Tj/oTQCRfuTy77BcQh
kSxq9CJfzRtvtCZwumB+RCP/+i308T9T3X+9uVZkt/wdAcfrEzfE6dPjUtMj
Lf+84W9vUSCq99OSioyOKCjJcWZ8ovWMuwfes22lx5Y/vktkZlQxHcdQco+j
6y+ymqzcVT2WfISHJ2z3Z2NRfIrrT0hnv9tdfwBo54irRKWLiq9ktKapUECR
KxkxtYYPPD0B1u3bCkKdP2N3w1vMXwG5OmPQubWDN/aLpmo+nXJv+4iqa6cn
nyl3B928b+SrDg3fAFGuZZcAIOSnBvM0ZmFMbkBUaIUenwe2bI3JHwn0krHT
7A/rRlB1cRHbMKVAciJGt5PjZG4wjWzh/zUuGyEa+83TlPKaH+OI/ecI3Q1T
6DZyuZtVBHE6A5Ld1pVLGNKE+bqOjx4TQnYAweRbHNLSWf4CoIpocAVwFwu9
QSWXEVSWcenlUNnr6VlLLIwFDMpxDd7sy1cGCrwInrnvk928P2RI3O8sJ2ez
iuXj9CXJy1fAqY/R7XxYKTW0IwkG9dKsc3VCBAXHc1mltwwsghPZVWOkss1M
J1/VsJkj28ivGBm/6PYhu0r8XgZo4ru6RGdbaoGyeiWg3slkuHDVBJvWiEYc
W2ArdY9Zj3ETzHDhAxS4CAWxP6fol6OaN4xnzfgpDqolAgGmbeMzYsowYJQ+
QvtkVGmAaDtCI+BNeKFTuKF75i61gAVTrhugIjeuUBXE1eg7sJsSbQA6um+R
d9Cbfh38QRmsk+tULDOeCL5OawdVXaYCWuGZxrIJ899SxWC6BdrMDDp4XJRh
DF31B6jjjlZxw6GGPOF3TWPDeP1P0Ye0JM00xQoEE9Mh13lX57RkMsz7nyMN
+sb/GSJTH5tXYwo/3VJ49odJvQZd35BQv0Ru3wEqOrtsUdp22zEII1TQ7ldX
KRhqjVhliBNdR+Z7muvKrve0fhQ62anvIAjqcX34d//Q6j2dgzmXtmFY8sgR
Jqcn60AqOtqKiUlWv2b61/hvdE7WLwvmOqVuSsSio9rAB0Tg1ktO4Jc3m8H/
BQ6lPMYMtwex3Rfw+cYRAiKLhUT8BwKyUjMybP918w7ikJTYL5jZAaPhuqjw
FX9zWbYTEJg7LyyxaLfw75zRFJAfqCrf+8x5TGy0lojROwrdgk+pAoNW92Th
4D2JaeqNCXgvpKTW5oC09CeZ+owIV0m2OsOuJnK+kRFmpuQmlt72X1XuWuyA
DxPb+RK1fytzJC75ZSNUEwpLfyk+0EiI2Vp1wtzO/yhEf1saphgu+AM9/UAe
7em4RFoEcteXkX7NuLtk0bZCUuogQW3k6WQ6nVC4MnF0ShkEFOuYzjQxGaS/
eB1gcer7EjobqYHF8+UVLX1e4rVUE/0kxPrUusCa1oDGzoAov8lV8IALhINK
RrS4nTygp2vqmg7XzMCvWPQVgLenVUIPmsF/MKdgaPzdzU27q3W1L/hlypVZ
2N83N4Om/7mUPJe5p4i3A70ZrHjUS0VNBQRoXIJExphL6opbWzAZGANHWEhU
p0WnFggQOFsocgI9QeM7+FjNgMYcvu6iZr63sCNHDOOh859I77HXBnj5VNKr
LcBFCaPl3MWUK4LzN/NJkJTPJ12d33DVssjIASH0Ad0YqbOk3/Am4Cpfo2it
3EgFD4H1lKd+h2l8Zr9C2uD9jnvJr/kP8K4OO3SIj1BAuKpodYB0G+B2KX0Y
zob+M/CACYzwqdTeH61l8xTbY2uoAiwcxLIwVeokE1q2YsydvPyCt8P137yx
bgzBqvkpW2JoB9U3BU0xK5MouztBM7R84QBUrmO3Cwkfe+boCDb+1IiM8yTf
1uDKYPNsq+qhwAnfXsOAR5UFVgCJzk5LzULXYysXfzEcjOqoZspAClHeRXcs
J6DF/u3MNWcKL3ssiS6HBUaPhiihm3/xM+leKaz04j6DKi3lVRl/knp5N8X/
5pJ9cduv5dW6W705VycE9ECs0SCXDtqFXdh5WD8GJ1s0uTkq+MgHdLxT+Ndg
yOesxe3qHja2/GZdgpfu6HefWYfFZjd1XlfugjBkBHU1dYwwloZSlHpBhbxs
4Lrjp1Yf1ucLtpJCZ3uDlxk+yh04N2HqK1S1G+qcV6jbQa50La8AyXQGJ1Nm
g3lVkuVFGb1vwg6iGSnMZJIDtQIPNfmotvxEHayaBH31CAzXIsozc+m3rEmb
gwonA+V4BENfGwRH8ONIcj0xLtAPP2QklvdrX/KbBUA0aCcQXbVpk66DdTO/
KSry5v7iBhjX+WI/IRTTQI+h0Bwj/ee7UlD9KboLQxak7kx+UngH5RqylDjb
jcPbTWtY4THIUliX8Gn/7xPLEYRlj+rmeEGgbSDJwEbk0hiRhqy3lSPHEDVE
WLJJWTz8cWsJKRPtTnk4P7ygdS+r2P4SBtESNgMlGUdzTT18waX8EZ+qTG3b
7E1LB1P+4QdfAwwnGgc7Z/zhgXVL+982kh05h2hF1IJ3Lvs+iMK76FmDE3tB
+SVkpB9LTOiVYfHwaPYLbUkEoshRSGkjMTyq7N8+KQZofG1ov9R/zIYo43Lr
qHJXm7KRBKKBOenkHQYUwbHLQHGQ9dEiAk70p7twxLYk+/XVq3MzwsIQ+CNb
SgWCB65CRWn9AjN1m64ra9+kSTK4kvXwgUg0RjZ2LRSR2tf54VcVJSOjfvH0
VzrY5MeqEcwU+DnFC6Y4GziWv6bUiUU49SrcJ51OzkE7GUzvSSt7FYFpyYNC
SQ/4qjKT+4mdOOE3Z2+o9hrzLIiyGqUs3Bl+U87bl62W16f8tGtbxUH3P+eH
osP21Gtq0Zbi7c6B+OUbKs7+yqQmu1S1fog8L1cWHUH9ou34ytakA4oYgX99
BeTAeYaXenJypxiJ1B4RycGh6wNfxILBFvbNZBu2w2KcArATOmfPnJw03LVP
y/R1+Yfb/2oOxqI6FbanekAWGsrZi+YaUodAzUtT4mX35wzsa1tWINLSHEb1
2e4gCmb9oP3KJtVwE9GpAaVwSiJJ0tK3dfIoTylNgDFr4bDDvWVxLrkLJCM3
DtFZkqexWK+MyLGE7lNDX6AQqh7z/56dnhn4tGdkSrXbNfdVA5wCiPInzTLU
Bomf+rZivB34ql6C+0opFGM2/Z8OXalcgGCJ4g7X5xH4BuflIC2RXozwmoZe
srifL84BBrFCPNUsz3iH4eELMXucvKN+piP4bnpbcMsjskHY50px8Tn2usti
2eMhUXab+/cJIZzm9hULgSyVQh+gVjGCi3BqnTcMqDbVpaHH191+l+O4y7ou
hY1hIAroOk4D7f6UjA8e1TDEC5kGGi9zPP6FBJGKHsPvcMfs7AQgIlb9FMix
P7bU7gThy+4GErfHVd8zSyqKGAloZ1aLVkuvG8TZzrOTz5rGW3/VDQs6rJDV
BVhcxvg13D9WFb9IXdh8pqvutxDn0Oq3ixH9iXVOhxhhNMgEkAun7vMYnnGs
jWFBdI22BfTMZPYT/zX3KtaarSw3F3l9daiD/ZwXj9Pz8OBZcsymMNj09QK6
UV47ZWyPvjJZEx0Vw07AVuQGcrtWkreAyWXpscc1okECmp5Na6qVjFHWjaa+
qERxw+9fWjIs3H4IdlEObSMhJutp44rhc1vi5N22S7V91HeTX9Eg/GyO6pVs
3UZ4yIVhJtPSbnqG8z5sQHd2fs4VK9T3QMqva5jGKAWOmqJuRUQVPqWnT0st
eClPlwD1BlfHCBcbFM7YHapWIRgmw8QXm+Jrg6t0ElpKqGdjGtlv51mkw4gd
tbAjC6k2lrwdQVnJACR+6w8OoH7EwO5e4IayqPYA1b9aLFVCg0/yhyVpHShs
aYci18Qgt3rWLNhAVsHs2blMAQisvYR8Z447KCHlpw6/ZihxrCv97BifSE3D
luWRV0SNXnPriU4IYCizwjLuYS1Ew9UsE5D5+qHIs3EgKKj8BBwTUcqJR3aR
JtfQ2MQ0axhJcb5xPTKoTfYs5H5KzKpkk2u6oUi2K0f0sWCjHnMg8lch8lj8
qsLfSvWmtkSEnfEudPJn+mdA8r6zHJ9NxiYC1a6ksNDqVnICbOFrktzSNUXM
Kwl8eKNHRv42Z7bcwaSiQ3dXHL0gH4jsETVTghoar67zhJHKFSYxEqeB4plz
kC96PZOL4rADAjF6ZSa7QM2kFjARrvWSA5n/vwh3POL4bcpahBOeSYfbHx44
eVP2VMrN3u405pz36WR5dGHHUxdQvKVMcoD7u6J/qCuKIRUj1+XYpopSy1D/
sWwB2CHEs3DtwpSX0zFslVmh1dUtHPJ+/+JShJKBPvDxPIYBk5mBZXAkP4jX
1lgxVQa8ENIhL+tvikPRljIoeA8CuHAzaKRDeTdrJse5FQyq6iwQkgSeBVTC
fLZzb0VpZlq9tPLI4ixzRdQe+9GYUWa7tPcKzdrF4kOmYzzqL4I/NDO4VUx7
sB0kvW2LG0Wehlv/aLIQM9fFhQeLmENPnBW7ZIYa1Le0K/0VU7Ti4DmlAIpE
gCG07pQJdS/4xl7JEDeD87aRs1Id77zHizFHBE952uEzoRdPE1vs/gE3WB0w
/u91d8RyRcosJTAzv6P9yKpXH1EhWKEkjsoQD2y+g7+7LTjTMUdjfCvEdXiC
VjwC+AsDtCFn+tsvHultBMM/gM0Tycb2zEeT3kfDG7c3O/KQW3SVRwXDuswS
ZQv5+vdQCAMfYZkmyVJ9J99fCh+1bDFMWQOucQImwfjwf6jQd9jt3n2h1BdZ
f5lplAcn/G0/5DEmRoKqSYRpJd0pKNkDFtU6YCCjYRlLPuwHOB3+716qS5oO
ywTigHNnld6ZtLD7Wk6/WviQY5nUkNh2VWL48G0DbBZLRYdus+awSC6JFfjY
fwmnUln86ZZ+iXCnb8+DCrLW5bst2g1OM10MFl66qlZlERsOj32j3ZVQ+3Uw
fmqRTb9XMUgWB3Di/KLs6451e7XlzHHZiDHub25zvCLjkGiH/ASVROyGL2td
HigHt8UF+itRG3Y7LXCwROb453P+rxFW+dOIOO3UxsD70nO0nJnPG4F0SBtw
nSziZM7xOkMTCcmnv5w9npkLa/dz+rVLUBzE2oX+7Izic79SplPCn/dh23B1
8IS1clx3ocCZhCP4ypOJw3UK4fcsYDgmtONPTxm9PxWsbB+VIVPmzkmPUftY
9TJ+B/uItheIyigTIW5rRX4/AjuUXN+Fp35fktNSgzeP/9KKFryQOCWbmUyO
46hg4k0imABfqy7/9qllTFZdPN9txzAHAhAEHgP9ZHNT3Od/C9j83X0UpGc8
/C5M/1rSD8y4FNqGd+9C/3MWSpb/XkPmvjD5bV8Z1EXQP2U2EKCCahC+1vVs
XyU1Dn2JXK/zennpdyT+vgtzQtsBkfly9FtR9g40zmj3S+a4VdSHP0L/ZQte
r2S1sDcFd9pWy/0MyJNTR3VLKtkUCGYHPpEO9Jy/ZzHaVM6b/7YugRMdx69x
I2tVR7uCpUQKIDodVR+65JWvbtfgUwRccFyEFFISlHtUW1UdLeHtqyGYL1FS
GVivotE2Z3C0ob6DfKZNuqprt6MOxtWsRKQLBTHKms+2I+hl/YVFuTcvCagk
vjWU3/4fKkdt0ZPrskFpU5jQpJG1yiyzHikeDMwG1jt9SpvIlIoqL8yuaJ2P
/wGx4i/YlU1Hd/1BR/abAsbwDhoXiQFh3EDzIN/jhSlNkn0RsaVrSK7bx1Fg
BcVgtFkOrK0PpOg1n0Gb8IvlA5WI4q/hQWtISm9eH1lvekfpbkrrTtVqGtdj
S9DwI4I3HfBPe0xvpJyih/FBx7jV5cwuqj57r6TbpZM/eV/KxBq0tOgp0lhH
Ld3CJ/8TEG0Pcp5kfZeJVOvg2qcrLOZeAUYNFJVOg+suWAvniuY6CcFA1qtq
YDPhIuxIorIiwr11xGVWjZZD1VVEJxShLV2XXruPlntCyJ41n2FlRasG+NS8
xJVNTlJ8q6JurnMP8DHZgK+xG3PLgtRZ4oOvfYT/pgezy19Uyu0pm/CeGzm/
MHL1aKMyA8loKnwOIs1fmyHnFHPKtuId7JAI1Q9WQmyeFEFIG2K3N6usY/FR
+3D6HpT9jHEJB1Nlj02AiZoRidqy7LSOTHAmfUAxqwBd9uzcb52iT7FavgyV
mNYwsWRp57yArng+bLm5uGwONmEawmy4cM78E2GNtBk3bNl9gI6sb3rjtbEg
XyGvqhW1LNuQLf0j7WVPnB3vfFspJkA6I4yqpHnuyHRcGMWPzOFI8Q1/vxYh
dXB9s58tnvTbl9Mq7iFEXllwlbOtCbPSjdAMUv6/Sd2VYs/cty72Jt13sto7
E2kFzbD64PL7Y0UcHttnOpKn4s7dy3x2byf1nNcId33vkZAeKLxS3HyTmZNm
l+XARY8vCe4L3/6BGVien9m2pJgSvQaAQs0YovyPcDnCIkbCt1bEATO30ABd
U5tixfa+iDNtmyScY9BjGw2tuTOAShStImb6UV814sApJFLGYoGq0fdhBVPq
6dMdSKsgjCAm5gA9OBJeshwibvSiwGNNvzvj5pgPnpSsMjMvDZQdeHAHBg0l
3vPftivsK6eZgAPzjmfUz6iJVdwcQg4zTKX+411eYAnLCnDJWub1smhc200B
S17HtKHVtn6fVGPxu0iCVYxHqzTOC68nhIn5AM56lun381pA29MHrEQafrKG
/z8CV0M/2UdH05JGQssf72QkV4pe1cdR3URDLVqlQTsmRhY8jB9QzOZu/VNi
B9q6JnBmgRoJlW+OwCNEwKQ3dyMmudaFFPbRtTkblYv7hS5cyC55xyvoaUDP
IqGliCg2eheDycIscahJv7rOqZtkc5lwxkaDfz13GTKZM4wFtqa4iA/ymnBA
wZCej5tqdKzIGCoqP4F2P25mgND1JJYWe40h3vV8J3+mB18dz7wnafYN+uDi
eDsye3PdQU8lXEmt0XrR9pL22YRO5YotW1tXSyfqjQyY+uSD8/cVq+HygbbJ
CgDshMtnOt196fi12DZ8IMiwQVsRb4JibZDMo0+D5IBwkdYxlPcW6y4/grlN
/sZTaLr5+hdLHvJv2PFX9wuchZbswjPSP1XEE4DI5UL/nfcwUugA9rgoKMxJ
zpFCCeBm+BmjRxcAoDvLLVL30vH0t9QpzSbp7mYU77GcG/OLgXoJj4m+f92c
kY7GjPnkcwTLni0dTwd5YEqbbYecNsXxGSb6s61Pc1qh0U6+EBN/E4toEGAo
i+PWSm73W6UEDs0iPPQxo8/85T7HZiv3mZyXjW6nbMS1ymtV4kGnlbcU13FI
iAscMl3CEHT8OZvBPaPd1yRLkq5iBCDJDJUJloVvoAwnvrbaRbmQlNo0IMRK
zjV2R02JMvpEGKk7wb49CESzfYYf051j8pYwuTYfy6ogLBD7oSovnKWplUOL
URzNyPZ+EO7bPuzTBLHyM5ksmtd3ErhUoOTSv+q4oQGz6fsLWS8US6YbEvHp
Je/hdqv5GqUM6UTchj6CkwqhWnzWx7v7U90DafHXvCTMC8nRXwJcmqocDzmC
OQKWFqD9wOhlt5lpsAl7xKyIqyiJ75AmtX6KORTRMoSW9LKVQUNFEyFC2SvK
vb9DbwryJeJdOHQvUYTpB20REfQAeEH9ECtvJmJiKlDcU1whcKIx3SXZ5blT
LLcBSxbCwFtfPaTNsg+Q05DPRN3rLTKH7fg4gYzKSxYgZKrrlq1r3Om/Tqrz
xXCv2AwmN/5vanzbMNkhiUmwf7DlNXZXKYlFXa73JvAW2lNlaMiC8nKXJTmL
5sFN4gzF9O65vaqfW0JLC+UwYvPxL03ASB+G3sZrDLrB5al1ZaM41V8lhxfB
osBEWBKR2/rHto9znbnAn8HmkVh6EcZMaq3/vxPIbIBaBJSPpdOecUun2qer
bQ/0/pvjFSVLHnXmeUXAKpIuZB5PxgexIcWXNC+uNtu4vpxGu56f9U92E0y8
UAa9FDIjjTAMP0XSw7/sZTDsWCf0aIjWIpqyP8CxDByWuyqn3n/QTkHr7nTc
tzB8u6qTAgqrdx7Vpo5JS/bL0Lwb2LodN4cPBfvdgBz7pGM8ZxXB7WvP63j2
gSMHRRz5VHL6rGKNmoTyah7Zv2WxzG1ceySDoVqnGSwPqhP8jQeOaOS85kT5
UuXRJielxUX1hEtoVClMiWW5ndp5AQFVCEBMkIYtDjOx/weS3OtEy011A1l+
1eiS/TOHiogywQaTWzNz4+Z3N5lHPUcqdodF0MKqzwINeuYncKgml7/skBH+
3jkzX4y3Ba3xA2M38YKXcgpd5bnPVbI57n8Nsv49oTo65uvipcMttDzQCX/7
WL6cdrrQ62mGHtKb2uSyBL9CCJu7PrEvlPx00ud7Gy3VWOBHyQjMKOXeMANv
sEu+zAqNoVeADdydx80pxDjqfuEIRwCB5yrRPL63smzv2p9WRi4sVQtNLXyE
yeanVK7Sm3gsR4ARpxkqPPahfzrp48wWMEZwdWMzHm3s8OYdpQsYHnEYzgxS
Oje+XBFqcDOGkZU2+pq0qngYUeGhrwAE1iVAxMcDW0uilNdYxvJAPCQqIpwi
Rxb9IMFGKPZjXuI6mdtrrqtJqAQFug3M5aiOrevd48QE2UQeO/YlkLF3UT+L
Nj2B0OHUwXV8SrHGC1+ZuNTn4S29Rzpf08DMtUXU9+rxOAVEy3BXUeEt9dk8
L+/cr256X/AYNwuMnkt9ajKgJarHKyIiW+EUUkO9NRHtBTGgHZOVQMmoQOLR
qubUCYMRhA0017One2V+veLdWG7fa2qVIj07GjtC3ovAq3mIwqP8McFYuMo1
hyHM4l7ECCiFchTLSaCe0OTv7byZEfmi5ET/GFE+OgdITzV2+jzZtyfh9VYm
PqVq2JHIOk6PyOhpOtvUCHMl3atgs4n4SbaAy89g4DJGQAUKDdvemkX1YbYp
PK2sUfKbFjfIl8eahubLhMW+zG37iD3oVpMBjpVAuDlyz1ADm6mRjnrPEMWU
qfAKr35Qno9YvCPEDKmWtmb8JXp0hAPvaRotk++PVCgdvxZRoVkC0eAtALGV
HRIEnRu8puONw+3JvHX9G1+TlkQ9e3HHqchND/DKimUueygydzrB6hD75dDQ
yCUEArV/v+gLpBsli9yb5sEcmdv8DD1iLFe22tWLZzkzG3tXmmGYZrYYrKqI
3dNS83oanbhecNlmKcpTJpk2EV1pIHkXY2261QCmIAebpAOjwYdqYd6r/xV8
QZvkMHhNyJFG3KIVAUFaybj4/6HAv7f1sGvw3coQRFPDuaan5JpU56TgNOxl
sCh1ivx3nn96afnH+v/Yq7dVv/s2URseeRbTChM/6s+vdpT/7bgb8QucOS0n
sFbugVBGHv+bTz/zU5floAAPN+oCazKefr57kwneI1w4OeE8Q7JRqhY7hycK
PhMPSqUzeELQ97FWZzMcRicZ+Id5JMnzuW7RVs84ETGNxq8FdjMrIiDeD88s
kKJAmgW0RPEvlDOvEWAW5TYYrumzYhTn1ziIxMH7eAKsZJswulAMaV7gs+zl
c4Frf/j1Q0H0cI++gECRODiFOf9EIoaIVSE9VvvcjQCixtITX3p1kwQnce3q
d3RdIHwhJdsuv4YBkrCeYpYQnI8PxGKqn34YzexN+K70QcxYvlFBO8ujrxtX
nG61P1EhdfKv4GmJCr/utpW3Ej+ZbB86A4RxJjyW1PCbhJeKNT/yXTwTxupT
osNVwh3/Yzj2Zs+1OhIoqBRFl1ImMPuWafOPtGL0XmiyuDLaZdglbLwhX4aS
guKYc13YXmECQYR/f8wnBOHUxkWhyGD7zVRsi4WaSr4uYPhnGMY/gsKuV4CK
2JzteDwz6GP71r0XAv3qn2yVMTxGUIR+MMQ1a11MX+cb6Bj16/ZJ1VHHs2f0
A3X/NSe9eeyGZdFMarXiAlykphLrzYZaMhRatF4AFi+Z59pKIe95Pd0mGSyL
StS/EPD0VWrH5bJ3t3ajZO9wqq7tZE6VzhHWL8F0+X7VwJHmGhTpwH/cNkJ9
fGxzi0YgWm90eItEebB5Ha1qYwQ+pI0tIxKB6JrbuA/WuEtncIhekPnNnyNU
DLx3K/UFFzXByfRJyB9qQ2KWtW7VIKdR7Pa4PiWrVxQN8iaDxtGoKXGJUPoW
lAl1Qm1jTwRrD0+5iHhKCdl9JR35XFEzDS92W4O964Z3o8qLJxceWHpwwStx
c8jZhmnzcYOZygLdzFKHMdkIlC5RDti/NJ7uUuSAPj4rUJ3LrNmPJjo3vcAg
ESeNHCWrFZxKEeZOXyVlF1H8EI9wRX7lH1Smd2PWFaS9cWyqhJT1CjHmCqlJ
bITaHRqzruZkbo2h4itINqT9eJS0j6U2xI6Dk/VLn2XxXs8B9sVRZuHZY9EF
4w5q27WyJaAVxPNcA9t4k0iDn/fqFbnJNxReA1igM91ZgG8hNOaNhgIE6Bet
CSLyX2qmTsws7TJ7VFmKEmHvIxgIHUmf0f1R1yq/2mngP1I3ar/ODWvBcxhD
XT3YsaoKWhZRcoOhiBZ2egAhk2VN9wokNCMj+Jdj1mMHD07A1J+N4/gKwAmD
UDbYeO+7ZxEYZGOmGYDXEWJVM2DPSJbMFx7kKvBHX4+EeinBfwBQwfGaY6te
hFkCTpH9U3ZXPHsA+z+B9OzlSMnAJqP5aldvnC2kYm9mZ97oaXK8TYwbZGrN
VbxBo69GVyXjabr06I658MwUgdTwL3D1De3qLyteECrUiVEVQwFOyAeWst9D
RMdh8hq7a6Hbccrf51L8OFqjqfCs5zeBsj0bG/E2aPvP+ydJ1eQVr19aLj1c
aip+ad95RbqEVYnpA6V83uBfwdVY7g4+7QGSWrFIESnmy7vhMdJfncDZbTIX
EakZ4emratcoOf3NHv1l1bCpWrdcz/jev7MJHG9GQcpCZcYglYyhmpyhNsuJ
CYsWzvyyyuCkupIEsJeMrhZIl0WWQ2pJnUbXcFJuvwyE5D1zxl2cNSylFhrS
dVB3iGd5qqfGrt1r0qg91d3HqV4tbcebU1WQ3glcIQY2c6EYx3Gf9AJG9KD+
6m/d1mFUT2RcIJTS3gZ109kcVkc9qGG/DXM0oJwqEUJcFPy6LNe4PE+BHIdA
dVrhSoX9GwzZpAX9KefXY9apo0uoQaFnRBs3WKODvx9dTG2URbiIuDdq+vpi
/zTl6s/IEMxv0nqzx7tCa40bhHXtYr67QKWk0FG71XqYnNDn/XihOXbv5+mh
fCm+bkxXms6b/dW+hlZmXuUT6gphbmKeROuRyfJbjX5Lah8sw+8qy5QLaTrR
4t1WHOeIW7RviP86pYHqWwf/Rq067/XkuwdCVRlVEPGRFrsbW2T1UpT0bkqF
j9f9RQF3wASxyqmImCLV0G9i/WWYzOdN1Q0yVdeXU1evXgQw3ZGOqDO+obAf
umn4VxQtgLfTcgKwCich4i5byK8gm2l+JVre9kS5v5P0udIF+NivWzhdnpuw
rmtRJ+mTAmmYW3jqeMefYPU2GnzwZYn1IVteSOtXQ3xk2IeqOIbtv/IYNlBm
DucsTRdR/287tpLP9XaJO2gUXA4VBmQhVP1HLcJ107tOWr2KZpm2YKImMoWf
++OyePQDP7LOfGBqw5WYrzFNFPDbTwHqKAtZJAPflzIrk7+ZVbPIc2kOEib/
9uuLgWq0Ib6jI3mPfaKoMWmR5OZau4k8r22DZ2Fi/EERVE7YgnnNUbEB/nY1
yvNuSDZRSnpIgZhrKwIrzLCVt6qwwQiwolJTbrZhYiqU3bM1TqoOQoaAURvs
JFhU/k+9DPFy/8tloW8kGijzmRYM70CoL/DNcPEzLP4hjahdRcxid8lqJDfb
DH6kG3KlYEubC4FhPWHrLj23ndhF2KAhlq0zNfrsr92TX0YEgZ6t19gNRxHL
eNebxHce7ekvKJi3xn1eRsJphoXSOgWLVx0SO6lyIKhrqrEL9mEw7rn072tm
b0ugC3D0lbevCjlEJKc08BXC0yPsFoZm9yNZOCYvr1iASgf2T6rBjF1cRA70
ZmyUd5lMMqbKsnU5jKsrUxCSEfEH0uGOHw7hjo8LJWdDyQvVQxq6Facc3VU3
JTZMssa3s9oaFYSj3DOBqRRaz7+fOc5DYaXLr5jYbvBS2YlSnE2UNnTyUSM8
qP3rTYu1klcJDHM9tPHFEEGy6SUTZpV+ZP8/RTq7R/Xa3dLNnSW6jdLBK8rG
NbRZP7o0f5Ul6kw/pj/xi18ypIY7J7yU3jSUV+hdztcT3xpbtcKtIlQJvYXy
FWyAwUemQekNVqNqyObHcGhXAXGyIugOE0AR5M3Gw/SV6lOeZSAyj7ZOUfMM
fJjaIGNlVHNRV6KpBWC8f6p0ltZFoLqisgE+wdF0Ru7dsHr4IAEEk746vWtl
B8UIg+nRZx7TDkQbZHhF2tbRywlM4XS1zHEBZHIaaKX8/QRDwQs6VZKX8rjr
dc9wTtQv2yUT/DYHly6GAcf1PFYtW/2rXNvOPUHr3dJq91UaLNJ7kbIVjEDR
H7SkJoZ6IdPmiPS7RnFCYUEeFz2zHMXTQYFnXYhozl1IIQbhcNIaN0e4vLob
4h/NHkje0h550ZhW+85xdvO5bBqhsrth1bTaCrzLIvN/cNr85kc5+1G7AxRI
BxFbYFZ9UtQwmhOvw0DeFV1nRju62PdGouKw7j8ZovDgp5URwoeYrSEMi5qQ
dRYs5mY1N8Yksk/T2v53lu7yHvz23pb+li95QJmaNEh0Sppd3YHhKb81Vjit
0Fki4I5Xi/jr0WdE7KT6aHRiY0lgpSJ835xuYlcoLb0xvezhO0SV+EwAJ7PZ
dIwzUwrhzgQJPoF1XbAsIFBcc+b73g6A+x/J9S4iJiQ3eMZvjFgPrFuY7qfR
4ZHVwBLhXF9B+AVOx8HdlH+lrrTf6ARjKZIERorj4BlI1CYODNLeqRROeb7I
3WAXjPZP7X7cmR5Oc0D5XfCokFvxsW0HTx8EG1HHSbZcQ30c2smg7Yrm5xEh
D6I7oF1Ut8vlIIt/HgbJVflliqutqvvIPG3oCJc4u0IA2mkMBiirvQnlCh9t
iFvlejPqQSs7kiIa1N8McpXKIyDZIZNQcmdAmPhyp4Iib/El5KIMghnTH9PE
m61qxDl3TYOSdlJHjauSe7RHs0WLcYrKj7GLoUWjG+eHIslsNqaFu7sH5DTo
W4KaIbaSUidrSVP4ajxMW3N8c6obks6fjPAMe8RuPP2Gl1x8vXY6c9sZZPlG
gAE5sJNb0fIUZPROEjnQvdFcOxjqcxHflqvMpHfCsOVgOr7cK3ftObhITrCd
lsUJAQriTFhoF/VAKcm2eihLRW/cnX41146XlDRC8Z+Semd6VUNCBzbE/aTy
URG2yWC/XT9Fi1tdlapym0KDBJeE842VswQnKX1xPnnKd2QPTGRQ35UCnzMd
2i9RtrZbitYYkUNypOUDHo0olLMOBfJ2UELX3sOkVttjzgaFaQS+fPbBALLf
JLEyH/vdUOlU0sjolop44E16tqhC7aRalW6BjxIjie/vLqUZeN0Lwad7YwaO
WPtp6n+1C+aN0NkIGxbxIdctoT7F0RcwKlEQPfN3Msx0qgJ6zytuO5HBHU/U
aOv/Vna0ZpOlX9trQYpW5J5eyhLOIBf8IoYqhHjBHP09NJRIqUKYP3mItHcU
rjrdJqFZJ97vCL25KBuFX006LTslFdETEerKOC3Bsc0tlOjG9lOnqHoVI/9/
3puxedfeOuYCKI2VFDjgYteqdmr2v7tjM4sT/GQmlE1re/6U05+QR1N93fS1
sx1NkhL8F05IWYVEDSo/E5K5YaI0F4Tt30Kl4oa05iib+nPtwioD4mQM1bjg
FRsf5Zo9AcBPVE3lNoB3csZWUDcXu/CMC5RpefZH++2jSPUmGmCstXw6QS2K
afnq5zfdsbEovjYH/ir9xn7FKIudf3IvV3vXjV/5/kgq/hdAN27S6sPJk5Lu
7Rn7kecmLMAvLNzaZdMuAOFP7HtDLFvOrF8j0Yn7npM3LELKQH4YoTIzB3c8
nHPzlGmAOlEiHBAbBlnpYipjWkns9CwCzD7ZQZe0uu0uKOCI8MJcRj4d2zwo
6kk+8sMxn++gOezO+CHMqO2P0qWIKV/ofdCv1LFJIPdj//Zv+Foa5j7GUpqo
f+91lJwaSVACPNFtzklVEDMwkfI8NxxvrFWNnZ2O0Ozk16iJY6JsmAVQcrry
phL4EyKAOdhC35awbzqsU0BFg6VQnL+FXV5dzUDgO6+sp4W7qjanq9SsGp6W
FtpHog1d655JiyVEbjaAlWx71JFwm1uWW9DxS2prqDdhTsFdBi2Yh/i49Ui5
cARhlaVXn6ADXFSqgOHnkXjJohn0FjOLPxVnG1x+PihGGlvSS914QrYQWREg
NG6SPkKEBA6Dq3OQoPkHUkyeOz16wyOrWPm43SNytJPslK6GFRbrCFEWr0xe
Y0ZF3ysjvuA77J+vBhCwCcy6JKDFM2NfuMRnHgDEWt4FPETXGCYvCAYGBOLY
tMhFji99wSvqXD/DTFl7GvYbtBuydmUay6+9m8tLBNIM9o3I9tlIOfkqTzjd
fwiCVHrHgqOpaUZ98WsLnd6XBN4EYP5oL5lWKTrG+MVC5l3rXiaJh4aYyqRk
gM6s/D5ZDdeT/IyWOu25wHB+X4Y9Lvs1Qe9kO/DTnLwiZzp9PZdpaJIeDewQ
cT6waw2BEvI9nF46J1mYPOoHxbad2Zjum2r+IRAno+hxEAi8F0vLBYDDrnMO
61DN90QcUtgvPL/8RqwTq+cCLj0egi1A6y7ps+E7pKw5bKbkVe2AUEU6pOpy
BDJsyUY3mpw3fr7rXtA1gFJk5gfC3lyAHWeIgnNvYiCercUn+hahuyibzaCn
i82TmbRlUIqDhbhhdXgtHKtCDVdehiPXI/mQ08Kpbzi1CDK2j8oqL5mW9aQI
DiUf5rPoeQ+yoa63Ka3WkoG4uOr3aFeKqDrv46Lce4UDjeIcIwrVJ7NFnu0p
iyw1B0afDBUulZ7O54QYR8wYxVEZG0hy6iL8b6E02Ixa7Xe+/YGkylinpdVt
uuesJL9l7C2q4F8oKI8sDrO5cHARbMCs3e94Qnl823T9gvzPpOz8HdBX7Nlj
HiH8rJO/oAnD40+ID3Pz4wQ1JCVzjHWoa0dWfujbWFk7JiUvR/3TWtr3tjmc
8fgvbhKFKlist48ADgqaf9+WGV3WtlKgywToNWZf6j5CO3eZsVcb/ldDy1RB
tyWkqRXlev4l/BbG4wzbh/LwGxwyXG1Rz0fPM+VsteGYCdmIR7+MkyiqbS9o
cHS2gEodN8tPWR920O5XG5pucejPJrUif7LpFQQGUaRU/PemkbehJlnkujlt
I0PXARnX+8zxZfy9kPxw89DZiWZiEbydssONCfjT5y158LyXob7dhLLG1Rel
iwFj5gsDg0HN8LzjAEytEskNCsKqSjLGOJS5RRE44h4OnjPuWh2Zd92xewFV
2TmZptydz2QCysVj7qppt0Pl98YFxCosSN1MviWj9G6CYl21ZJMOhvAZEIKM
AJcTqFHrqlCnN686PQEOARZ3eqqOdtVfqVRI1RX0Tkd+zlpzqUJ0BhaqztNQ
eqXTdM2gB1+NGKeEKfl9uLLsCD+qbiP8Y72IWbc+DfOgnuAmSgFZ5gAPo6MA
n5OrSQErTRgDQXqJjbDY5xQPEdwf1kEeqVhpHyx+jW/A030PkZtXlYMRC18H
KFADUJzKFFen3Hg8bT74sYbwDZqSjS4B+uyMKV0tMS8yhcwtf93XC9F9tDA1
gmOhIit/dSek5EdqCcpjW/Hju7c3GwhXJYu5+p7RpqK4n2CnvpA/3PcXmdoa
nZ3DJlhFZ/vbGFxN5bx79vcerN6sAJSvuh3JIPvbTNv4+tj+ZEXNdHkLNNUJ
ofhYsULGE6QvBLz+xJ441Djw533q8NduNfNI/KiaPcZyFfrj8QCKX9SzwySW
dMw5i87lb1U5y6HayzeD2Z/7zz5bmLC834UZFYAHKReqOhVDqOe6Jq4r4lIK
4GRgELiCSdYq6yfVvMwXxLLvdV1StfaUiAhopHOtHfv59P3FR/bIBQROmss0
xjoA24Rx6ckqoR/nxGSq8OmMIbIa9aL1Wu5+LM1TEbRa5i/OfkPlqYqyitNa
jkHBlbkoxkd+Lb2W6XIJUNGEso7f0mrMkwaafZanUYNqyIftQ7owwEUmeRhS
r6DTgXDgJTz+553sfkVbVjOGXYbxYGzVXhEuT9d+QaWe+5vdhLgddmZ7sZ43
DiK/bcWh+ipJnV0qdzNjhTzFOHDasHZb81ECHf81CWhObpAgECYap2Jhm9+S
CrsW+jgt4TJ+lpWxeS6R2Cx1Oy4KnKENMYcRKXrNpZDqmg8eqaqcQiowzhqy
zaf7IySOKZ1zQROmu7Fd+CeuExdZjQBoXe6zdbkkhjO4sm4e3expV8ztrv2m
AbrsZutkhjE6zn05FL27hvBisP27T3LRYrFAnMzI/BRXyC5EMSsI36bbLDOR
yBJU6VJnSujKhQyVcZf6+wQiJhdmB05ubYwxcFcwpakzy6IYpVZ0gXnyIFGQ
Ji3RSdzXv5jkQIqyaA4ezz1twzyDopUuaJcA/NWc1+v3id/Tpf6kSXzRQmlk
xUy8I4SJ/C47fGdMPaOjpxjgW/koC7OBPfR+i+r0PCj3G410E3Efy8C95IQh
oGIj85jlNJYKxwci2Qdf52XgjebdRKg77vu6L/q2tF+WTSZ2gQjEknZ47mpu
r+90OSogEISFY3EUGsFrcGWpH7t5xQjpaufm6YEaVdC+kPs+7pbauGp2CHum
1LRTmiqH+PFrD+q1zzZ6PNttHSh5dgXl4cqMN86Axi5pm/jZyJ1PxrZOmDgy
lpcPqnk7LxXw+kE2QXqRbFq8tgcnU+z4Qehd7uSNPBYvvVQDMUcYdq4CunGb
zTnY00mDFTy1KiUJLiqUB4xIlJC6QZNQkvQC4sqXHnaSqVibuPrk0GTPgP2X
+N5dSuIFVGtvVBahAi326r1+SfJFdJ015rZLn4sr1wV8OeQnnorMobf/B7wm
C2KY+O8j0/EHlZDYx7kWbl4Pprwi8q4FrnFF5ZMheNd/tf/HJWeIybv9wpRz
ciyuQd7Hlc+rXrhbdKKIR/+9LKnqYsF6RhegdzigvSYuh+SQZYZWHL/ziNYH
jpGSqtg7VcKD5zLmQmcAgN+LP0vdItoq9mMO/a/p53Y+82R3YkLOuenVIp1C
iEmsjws7HhxhmMX4v9EEKHoiVk7Oh8A4aA+AZjYflmQ10tcwT6O4DPTjCZGi
a/fZaApdTNPB5YDjm0UqTljiNHiDhRWm6BbDFSX5xBbz3NfHuag5Bf1dzupb
K+ohtylxG/kQY2/Xk/I5vFbkOYordULK8XuzJS1UwwLvEGJrT3uCZLaOa2OT
awzePbs2WpXJt0y+gwCJCvqEWznc9xbF6OBOXYiujbx7FPUkuo/+COgQcqkT
7asNRAQKRAT+0yDm76MJU4ysG3xM2fth/YM6eaMtidaMaaYcLUV01fcUZnRY
4+5opcaF0Jk2Ih5MUNWDVCG1CXK4QTyMWj8xH0f5q62oZz40YMZDE4IkKi7j
I0iJZfHEDAOjaur/PPDLsE/UUWVMl0FFqxjfi5vaJQGAFmp7ok8/E7jMpVtn
X/dDrNaOU906XvSPosG7fOGk6at91XObxZZOagxNkUcJmOmamheYvHe3Hly3
UEQxg0VHgud4pP9uu0530Eo8+zAon7hDEbUWJKtrXVELWWjibkAJ4p6n/CZ8
7MmJDiKAT5peImYRkdZZqxWS8ZqINXCI8xAtf5wO3UmEHCmpg4qKYtKNYofD
kEWyJjBtnrbcQHhNnodTfDcHeKeFMpcAVI8wb2tyeWzxg7XNVaFCsuUMxCWx
NljeHZdOuYeng2GFZClJLDBpiQQRqHOUgKEKNncg+UC2brkhohS9jFoOYn7K
nO+KTV37lHKqDxb4DixCh8Uu4V9O2bvZO+BW/3D/N3JgYMv1+8DvazljWv2K
vYsQ5yI8XpGMzdWPeIGFWFPA6Nm11i1J9zv9NygqV3ZU/jxF8C8y9CXNG5fK
oBUn5ZyVZbbpiT6N37TgkCdET2LVmfEXGa12mr3l/1GJO8CHO2mQwJm6s+uo
XYhSas0vAK40hHw7/xiDb2IJARTj0UnNAkp0n205NAwNr4aEakV3FIKyV4Cu
U3VVsmYqO8c7RKWNYiyTekLyTjlGyYDj0efRk4TPC/szVOAaKrU61F35J/63
EHDbUY9LcNsUCpj1jJrouaRJ4xRnjndwVXIcRTXfhkezYy2WkP5VM2saUznj
1+CMB4W6wApWrXk6Y66VANjWwwYAU1D+JhK2HWFGSXe4xBilG6OLW9cLeDYu
yk24ZySsq4GhTZCpTCT2ydfM0repkkMYp+sb04NcvARw0Sp4H3+b1uVttjmY
ElEl0DFqcFBbDhHRN8+iZhaGP2GsDFNHommNV9i9nxNSBt+vZtx93DCV78Ye
ejmpf5gqLcux27kDoPSXV9kDheuEheNicIGwxl4en2lEC2rhCzQTbIkCM4r+
e0tR9d21NlDszCllce600JfjpmRp2lZ/Mkl8aNl2pd/eFQ70uqlVk03mKrjd
dtPE3DnhDVK9dOarU0Ga3kb7RJCCW2xEniQcRJPsEFjUYCbla4O9g4PisFld
5AkSfB2/FQrba1Pnr/OtyhiXbvrJuOwJGnRaZOhGB9KNFVZ4Zhhi6SucvNpm
5OFjt51O5yqcwTdh3Wh9hamijVkFg3lCmKPGrtsOcMWqbXBmJOm/cankm8fR
8Iy19S1RaYdvk0ptEUaNZf3jqYVVT+bL+pptqC6Sbpex2ynpSd/wm+X9qTNa
/EJtFJ/hXLMuOkgYNW46IOih2R2wY1P6HJvdcHVWY+t4OVrg3q47PYpxlwcB
pIblDI9RYd7PeLFjb660skWgcKUaLLmYuQN27wiLN/PAIZjPLq+uymUjwwHC
8pCVCzL67eSTKmcgx2Cqkvbj48UNdfPcyOwdM7Xx7ceZVYW6sPGeJhzZHWU5
k4uMvUTgebYXbc5k5lP3H7wJqZEuTg91MVjwNrLjLiv/wd8Gu0Yt0uVeHVVs
nyF7QlVQYgNLd45SOBGluESG0E2fWjyrpimiHvu/HlgxsBlwDC46V84mheQ7
TakQ2HXXH+z6MDE2bGP3Qd4HWxuuoCdkIEtsCIes0rcihZ2DbzAqoNfJmDRc
SPknoM0UNlDeEWiNM1nQX54W+A1S8ytnoBU0Bw//J8/APcxYxGpKzgglcltB
sut4ptMuHSuLRsmuvv+RDDDFy3gpyn73boqcLrxUOAFrvSV4MJUAEBwDTtmm
2b8P/rTO7qAHA9w6vSSMXidhDcacUVrT95x9vesG4/skdybucEERbaKTNfAB
Kgmmnd2BhJOa8Rxgz1mqEAtt99MdhUict8dTqAF+2R1ytyo/sFHZSLdNO8ew
Iq2sITFO3wNzWRcESor47v9Fp6YyLUCOFCJkfkhKQKYc7/BpogHg/uWC/mgM
8TQidStkXJ2CxcjbtauYuOPUBnjXa39TwYlrhqLZ5f4UYg8L05pVC4Ch37FK
tTc+zy7ZWsL50+BPd61fnrtqec7VcFIhmfvJgcoouVZksdISGS7sgGV1bkrh
t9ctUgCRzpk302ESbcIq65/obaiF/PPrPzMM0qXrqFZ+ACh+mTgfMfVTUI29
OKeN+MsiS3qEY1vTjK9viFJbxJF/+qsJqMbcvhKTXp0uucfrfpppr01xgU2x
GvLMM/Y5OLuzp9e5erHcr0juYf6ln0fFnmgTih6uARu2gq+ZfReTgKV3NdJO
ewkVnf6l/QaDKC98zMnssd8UsCtPCs/kBrasi8ezhLDa2wYPNvLOwP/Ivs9j
JKqABKKEYR2oD2Y36xuxb/D/ZyXL3FF7nT9/B0x+ASbVk/IhU/xh/eOspg2Z
A737DvK6Y6Kr4rSzPcithHoosKgCR6wTjPcHK1cvszxZHQGwvMvZJnRkySJx
WQoAKDCdEVwfhS2KBtXvwT7sUqkHZ1AIXFaNf9qQQTe9IAHx6Bg3rkUmT1Yw
WW+ni4hbFVuc4MgwS6C9P9N5izt1yirZ+ejXqFb8VYvgWikuZvyv5MiSdGAW
KCNCKVRzce1M2PdTDrb88o+hOUURdF/pkDA48/o/2MBadplqBmCqnyUaIksu
IhvMzyAuW1toGHMQvxM2/W9U5B0HbQYdeF2HZ5Jd2V+XFrpaJxkYY/JqE1jf
1iXncoavUw0/nu+B8iyGB2T+jsvyi0bD1YCVoGq6CfFgouuAZOGsCgF0v2Pn
9ihlpxB9SYQE38Ek2Q3D1HKKNVW7nlRXTtVK4yD5EZZ+5ICQQJcWoX/aUQBd
1IN4OuVqyqXrDAOUEOU2bGinXE32NTlAfinaZyCU9L0Cswd4HPO4JzBxLuWi
Xx4faEz9sHz7/4BWEJBnxvII+lhxI+/rthFycW89tvV1NqLtHujlMNS9UBVd
b9kphFury8CjyhtRT5FQp4lyF6VySm3HOfFLQemDkSatwuYV1gPMAIgnepnu
Wpc2kZQ4SN6zsNjH5oJe6QJwdoLvO7Uf4FYnzWduh/NaKeh1vVcZJliEkDx0
1fzskw7jtY5TwszhpLYZujpGnWKFBofnwKKYeI/EOj3Kfpt1WUNJkiyUswz+
kvZ/XAjhf6CeSPOwV961zD8ZoXWOAdnbJWz0XIN9R1bdeE2lpNYaAMus6RDo
Z4gOtq8GnnH2uOtAqupo7JT8Z8mpEJXXU+aFqxrjipg6PAlZZljVqsr8ECvj
V9j5ny6E0p4swCEY3iU+rw9cKtW83uPU4KL+uQ71sv9AIP5wBhaG6IIDpxdV
aQMuLuyM4weYyIJ2JiUT46N89XAY3rChRQl7dhtIMcR1jhC4clbL3Lqfpn6j
KsPTvytyd5TJ3DG9R4E3QItXZVGb/KNlsj9bwWwMp66U8f7dLmt0wA4cNTUJ
0fd1f5PQe+YtF1DsRnZCLFDH+Z6glk9jVrF/OD0mZrzBMKIeEv3R/259ArY3
0tcmEyqcxLqwqrGhQ4zjGsO6K1qLbSUVoQEmh/LXoYmrIK2T+l+XgZn4nLpL
wau8Tc61sTHpW49HG4bQW6oVQ/CP+W+9dEtvzbSsdcMaEVdduODR0fWTRcPA
ZKtDQoXBZ2LgJjq+HEMC8l8pfGv6l0i+PncAtOi2SRnjJ/a/MrqmtA+tEYJB
mnTbox558VA5R4bwfXuvPMNSfetVcMty5LhSxiwwRrKiSD99Kdu71NThkhcG
71qqPaZX+utmdz+7VJfQx5FyA3CXX1pez4yFqhAEf3suJ+I0F+u2GdUIel3Z
VyBc9MeuSz/MhGIXbs5WH++/C8D0lx9gcvFIs0+Y8lgofyCbYJmA5dfcLQ2n
s13ws1G8E5Cd3L4MmYNN9lcZdOaG+NXh9jH8uS6+mQrHDGtN5xtbbN5pXZ+B
NZRFuzWBRIdFTbxUKs5YXvwvX/5+cs/jmHdpNMjIPgqlqT0uJnd3uagacm20
ocXjz9D0b7mVWEneGyeaEwAYuo/ZT8EbfU8Jvuc8FoXO0a9wVAIwBYpLMDhz
jP8XgfDptF2UJhR/A954jsnbZORM7vJ52MK6kAbZYg+3xOjH1eVucce3zKIV
ZOZOaOsfh2L+KVLcY9agsKgwfbFIrp7tDUoEy+E9wCRivksBpa3Fp8XCi11u
CbK6t13dXTGn9ZEf1dsgyphBsJWdjGCpbO/3GSAny4FekGeVYPSBsBO63DUt
pv6MO2k17UlBaJw5r07YpStQ9V/6H4Pp+uKGrcqeXCRvlJ//xfJNo9+Xi3uK
Cycx6bzAzEQzMYGsdfDztZ1ojgVmh8J4YRjWzdPzdjrxLbnVVnbuVZnQHYoW
IbnfUyTp4mOhGDxJOy6ovKwJm0gg/SsVrBSCeSCt+xGa8JR04cRFkbjOFW8G
7wRCWls/HnTxmtEvy4DBV6C+jS8sVjnQb2nZ4VmwQJteNAaJf45JUGWiO0Sm
/LPDhhNnjfFixBG2SRwJm5kkJiZHgdRkncK3H4AqmHh2MrfWyNNqRQWnJvHU
omHuQt15At8O1lot+thCl4N+vqJ898sW5lT3UDFLpxTId7rrcxW+zlKlPi7M
JGTCWcp+FKcFFMuX/bUfkkcjWIIEs8EtGqkKdV5uC7RO00JLb/MCyLtYoOpy
0SfWwYAgsf3+WPQR34Bn48tJJg628hBlVcgVdhoas+v39+s0xVAZOXUt2+cl
P8kZlWMp/VAg/vzYjSwdgnyizHDzHV8Xq8gmGhs/NBhYO6CHMvJ7JAWpTb/Z
e7YDUmxfY6mKbnjy7YPeECYzhSREQQ+WoA6+SewVnyuEzopISXYC3r6Brdow
UppILjdzbiJNVWX9KjtaN701KS9/YO5ezi3XsVEo479aRK+pB18/J2j5num+
bhRkyGMmYEtCjw70bsxIUxzE1QxMlTMCogIvOtbCbnVcY7m3UCUNVCi/ACsB
5/j8zyfxXCxxvoI2kRMZDvZxQhR0yVXN21PY2uBd+zt3o5JMAVA6Nl8x9NEl
MJhdZCkItorTwzMsIGeCei8r+5jXd6tqBr4F2TIIOfX3cmZHODIH7ZSPPh3T
/+8FZ/dU6O0iIcWASBKeTmz9NzAtUbSYRf12rZwvUqJ9iNm0SWwUzZBeUOTw
p87XIN56HLufgusyarL1SSRwnOn2uNHiP/zPsZBEodu6iTQLSBpuKWgXv0Zs
cmK8NifTgBP/WiUsGUD+MytRX/2+88C4xhcBjqojKPW5QedFwXS1r91rQ/iZ
5dGruDmr0yw2/7v4CcOPst/0g8Yt/wg2CTCjq+EK2nsxvTknMq/KW5fs4SHw
RtU7xeXDzDgEece5ZHl1buKqfV7BjMbJzarVWdKUvf6fKWaf2E0Jn6et3shI
YYuwJMfwhWr4mDwcuH/x28hV/NlxAobHFt0o3ZTW4OH4EWifsC1VBWwjQJ57
Oyqao3u/awPW61Z1GHOtT1vXfIGLSDk9AzWAmSRNe/BmIQY4YA777bIS5ssa
TFp/Wzw2XsQehDHX4BckTF7ZZtrVfX2L4i7gUvuU63DL8a4VBCbNgVawgyLN
K4CJzslAztOTFSNDrgpyBvDZocWHSR/lzOV0W+nexoZshQiaT4VdvvYK5eSm
DGTG/5zbl77CpuzmYP8mCB+uXo43nOUYgIZ+KEUSnMB8+K0QriHJ8qu6jloF
MehMTy5TeZzEgTAs2qzDnSy/GL1EnOC6iahn+UnivjV46EXDEuJfolQZX5dR
UmSONcwh9m8sPB+t1h3Z7pKgyqyK/Rj8xRcoynnsdAIBwtXT9d3T2tN0O3jf
+j1d64qer6uIdkeHxDeq5KuO3ndJV/eJPTc9cMlmOWwSd/JPfeS9EGDWYORB
vWObG9HIneY0Q63uv7yFWkEOqIPvGXWQb9SeWMZcDL0gHIRldvAxVCX+a52O
fO1hCIfIuapIWuNOSoIKO3DqO/KbBECESXjm1zKzlgwmUz37wCN/dm6hlHne
2VRd91/HQt094oSjLURNf2K2XkkYNrS38V1N2LiUNVqEdab4oQVr97q6yvoK
M4UYPHR2lnCOVC7ff1RofHuVvG8nrlRnS5/PY3mBhnd4/O6XQvfQHPn+srRU
7XnpKOWmNUK+BQ8iHMBoF64h0resKmmZVm3uFO1CJWg3sJxR21vcfEP56NFs
mzi7v3xW34aGgcyxlOWmPexriLOR4rap2spwuK8MVTNa2cD5rcZ6X/ylQ+cN
DamPb0wZcAd2TaYLYHltJvnfXTBkMEUNdkUudqXO9G1ODBSxyFqcTEgrSetH
8coI2wj+IgyHAoTuYxrZdjdrabXhIC6aa25fD1HhkvUqJP4Xxj7draVmC0ux
wMj9umgwOpyf8cmN+dZJ0m2ZzKEY1NFFxWQxAbdSGvvdk/unqv2nADZiFHpC
9fx7TB5FWhln5d81cjIKbUtyL+MMhe4o3WqcFRfxk9SZ4D/xUCk7fADthWx0
c4mqniKeqFQBpOBB6OkrtfATzuAEp0G5n+CyUtSOXUUTvqbNVuhBnfNgFM5e
k/KR1tkaIx8lXCIXAD1u9hGtDB3FGgwQixK7VzG+ghLYSmsrLtpMzxsCKtm6
rMYsAUtpGjaystqsOy/d+omMTRS+RAMsjrdDZJtRiLIIMXXc0xnAiD3ShbJC
QzIcv2mTGzUdm8SevvJmzUHXHoDTeyEEYwSexD5cTyfm59J0xmh5F9GoUKwz
oYgNqHha2rzRFRdO0LAUD7i3xqLVJ8kGyWAkg5A7S6KdeYjQPOoY3HzuGGXW
O949siwCo/DVPQldFnLFKLZaoMehWZjm0TJT4l1Wp95fUhdjK77+5Ubj4pl8
fufmntRn8HmGTcw/3h07+XkNhjEdJ7pVouYCswZVsXjSmZtaRfPw0k0EUoRG
7aZgpL6fffUkh9kwGLJsa/O0jVErJofh8L8PBUNgMI4nD1hemGXOo0MHbTEJ
DldRdmC4MwvWbUmdetHjXvl7Ga4nJMUBFkibv/fWqQ5yvcGgJZ/Uh9YYEl++
BKDGxMeoNLNvZhByPLl74oE2PRzITjhZa3Yg7JvVg0gbXdu6peoAYl+DCVOx
uiDoAyLjQ5Af09EmRG+I2pyrdKMJ40DQ8wN9OVu61SWMNmGJ9absSOrt/ZSa
A+/DNllL8Tyju23b6RKUOmeD1M8To7L/yME49So0VJ99QfNL71bt6pFE21mC
Fdb7BCkf1TQIZNdMBw4Yps5HYpMjDJYOVgV7g+hMMYl3mq8U994sK+QlgA19
pjEgxMeni+M7l2rov2hlfwCGq0IKM2TRMGUC+wjXKYsOgaw3c/wyQYzhHh1w
4gjPzl6fLe4DSqladOjdr8tQ4zfVrccNMv98at7sFjtN0yekf8WEaGKJp3CJ
HHZksUBMSbSs7dtc/zNG4yh3T/Jz/l+9LswXP59yudSCWZCl3/PFS/PtmZYB
mAenicLVsUcGoO8ghulvR0MSQwZoRq7kHVNye1cixWc8clZJMMwiAnQCBQNJ
1jHM2r2ZSEjMP6/ObrGeq+KQ/eH88iUFQn06rbxo8qHp6o/HtizV9vU4ft21
sWedJNHVBUsNeBI+xBLr3/7ao7O5Qucqflu6VJlwEwBeQ0iNi6tugRhUJnZp
1pkj4oR66oFBLyqVZ1crkV8gvgTzK3Ow0YyIlXQjreCLgZs26/6+fhxByG6/
NqY7dReEafKuMHYeeT/eDEuvrfeNVfZaNwS7LX2iNBgYcfXzdAVyjQR3Q15g
5KLni8K6fRkghZyCZ+ePt1r5NXQACmfhdyUOAC67qJYV11IQ6jR40/YxPSR2
L1LkcJCKKCALgOVxgP0mxfoBUQsIE5VVwhVsUzQIIB4uiDjOJr4Txb2GOGfD
qWCrmkDQSEXP5hmQLhbyZIXw7c+8xiKS6a/hqg34gBotYLR4YGFrFRUAnmS2
NsHocdlKFoGnodGchdjIEPKt7U2sipAo2+q+a3vXzoiQ8hDDIwjs+1BJKfrW
1Qri7sQONF1ZhJj/2f/KZnK41/YNYraj4JTVwulRyTCRtFBKnXqp09l4wVEB
FT/Paf18Uz5ZekO7lRJSfw3UnqN0auM9tIdHqQsrJ0zIvVIlpi1xlTGq3g+G
qpoIIA51FsUp34EfrjkuGhXFSyCPnasJ/9FZHja85YJHMc5DmEVRMBQEZT+q
5LZFO/s2ObA5RzL7jxGrpTnrGGrxGj9MQrzCRIJe5l/fxsUUe+jS8YdJqAeT
FdJql9WX7OSeBbhJwBJStEd8hkwT5jGheuVGj/NtQCVaBhq1yTTPwQuj9loU
x7PDB6NcnWxezpLpVHJ2j6jQ7arfEMqdY5vJ8Izgimq23dwJFY7NmSFdpLhC
eOMVkWq70x4UBo1EWsfLGT4h0zBpaQ/SKZfDIMmrHDhUsiDuKcm/ycTsXBw8
JFz0KEsjfU1VKewktFDSrVAjwlSd+FfhqUYAhClrCkb8NSLX57I7f4dISZgv
EVeaXDyQWcQN92hVGylVQIKgALccHSdAxZ6XfSjYr11MUV3pt7Ze+WyppIIq
5Pnpq6nPk/e9UyyweE+TsiXS/+H+bx8/0ljgdZQtKkUrZUOkvKw7lXVmlZtJ
Gna6UThO381L3CAUnR580cVuXew8cdfl3kB97agfGrwbfKuin9mKHapUfQ0I
Iv1no7KYagUmBzWtFLYIou0NFrdYaXu04gaDywA+AtG8FEjNClbTGlORAsDz
s0BSH74ZKTjTFToCHAOWs/m5zwa6v6tgYnPRZ48A56Lr8Ks2eHPnng28QoEB
e5PU4OUoqn4Ybjy4dYGbX0ivzIv3IVU4zMdNMu8mq+slGqaxM2MUoeB0rWWK
UggEJ8xiMelzgXuZE7ZGKYPUCjyOyWmvzMpUQr7HCOEhoaLLzV+ZldpXdovZ
ObiIZUH0sA9kV0zKeyYWbBEwlZgKJ3atLyr97yUsvg49OR0kRKh3FeQuw9ss
3as1XhNhl0YYjFb64bRtwasPf8gjMLJNYe0g9uE88t3yqXTrdD98nRDE4vn2
Q3gHCQyf3xFZKpaKzoPBBuDW7MaiuJFAMdVNY9L0TSuKli+Be1smgqw1YsQc
xqtJN0E2ah0eH0kg4TyBbo6O/jMzlxzzXTVMkEbB3NWv61A1fjP2ZQE353PE
3cE+t51oLB/axXfhs4lv0xZHRj0QH1UJw5EHVZ0uBDDXu7ReoTggdZWqCntg
KytLok7cHnlV/EOUyy8F2oay9nIslzvFCqilbdOmk9xfih//7l1xXTYPCWaw
icU2/Wj5qhmCfwbt8oSrnV1nle+p9nbliGabUGR1gUnvUE1qzoE8Fs5H7t+A
Teu11ImhsdTRh0DZ+9QwKpYCEp8YdaaiFKQ0mKfWzZYjebVk8FemT1FYd5Fr
heTAlZ/rNJ8xSCBr2GgO/e69Jq0Z4V/9B+K9LcBIvgal3PK1MuP7JApyua3Z
JaRwpqRvjadE5j7Y29wBQUaha6cl8xIKQ1hXoUgo/FKtwbRmNFbEPiPzxX9k
QSh14pxE6+zxBz/IXARmauMQ09uzbLVlQVkqeRWALJyCDkX4ME9AaSi1QM6N
AM28BSS7+Du2q7ynIhmGrNZpnxPIoNdp0LgJ8k/Kthkxbg5f/KJVi4QLNGb7
3a8BLBQWHIR7RMcudZooWFKogdyYXIpMA3X7bOphi1wvMm5I5Op1GbYazU1V
sCVS3Bu6mJiT9v3NWPhMYH7nTgLIl3EwVYWieWbXnSWKUbsbHJuVstx2n07x
4fe5RToFr8JDTd7ERxSyN0mramd/Laz2v7pniP6dhDGHNZ6PC5uQWnroMR7c
bmOguBZx1Vbi/eN5ajB/FxV+5GGC9HhZxwYELBL9Kh5p7wuJT5stT4P+6yQ8
a5vUnlUnI+xTq3o53ZMo/TW1SF1I2nEIPQprksyBrQcN2VQ1NRZ8lqsCRRbi
PURHjI8DwPqvQN+TTG9+AUqR1JU15zR85rsfrMf1Qq4WbZ9m83Qsoh/hcc65
tPP4U6E+3N98GhSVgKn9gmZu4EvyDljVwWWDiKB7m3kWcjIk7klbBCIbqVBU
y6QKO4zdxXDtH++TNx/wRD04E5ghMzayMre9ni1YPLbzj4lHC9M/L07rbebn
8xGYJdpIfPbN8EGQM6NnBbt3+XpqLH6RMQ4BnF6Dr22TtrWCtkSF5Gd6nwq2
/YlhnsZ7/bkNAzLyyHBCfvfd6nmSWoKASvFS8lFaEZ5iUD1hsHqO9Uck+aIW
M3QTjQqJ2W/P/oRlO7HoOhZw57OGBYM2Ykd7SdWxjQYy5nPGuxtVMhaalaiM
UGgiYMf18c1utiDukXNxLEZ5JG2QyzwsJBjhMvRD7vws87L7Mh8yzMnAxRZ1
zBbrn9TwH5cQ52VC2NC/taB0XlfreDTOeSZyb2pqdj9r39/Z4oFLcb2Bok9M
Klr8bkdVknWKmFGJ1y7rQ+WS05USWkVLR6NT9JZRuE87RXUa8BTXnF+9n6Hl
d6862qapje3LfUbBfRnd77Fv4foycmyztTe+UPr4+cbVnCMQSH+0RETpn1Zw
LB/SVqWwZOI2/Fsh5MAO4kK1ZSON7wedygy50lSbADEjyvf8QMmxTTeaGdoQ
XDTI/iNdxPOrDeI8yPusOqG7IPP0ETr615bdX0VG02rzI9zePIcl3lsg6fp+
5uukL+Jld2urIIYCkvmHlxaPtjn/xGbgVpidjYNw+xMCzUgY+jfM9iKx0UWf
/9nd8mJqqCPJPUClpTcMKvEUF3Ufs6Gcn65yL7XlOouEWED+s3sJWcjIueS4
fK9MwakPq6xFxYmAEI3wM/CCcun2RULdiyZsmdYL7T5zAg+sQgk35Lc/9oHR
Wc7Ej3CoFMHnhJIASR+xfoiUR3HN64z8NV9Imiglk5sztRImGCQ3UIVCaWm0
2Ev5lDZOnb+7ctm//MV06+3wknorc4ElzvuchrEjVQWbJycYWvDg/q4v+oqX
3qeREYdxLowlPjzqSfJD7BSLwEjjsAL55V8azR0++KbVZ3goMdw4XSnGo4KP
w4qUmGMFzuhFdTcVoEaKIbNlwTL73LepM1G+2d1ymm5OHlTuU4xU6R7L/7UJ
YUWYKI7vKw3ePtGaNbPIKiTUSbcCN2ZCttw/FPKo3FciKhDZIabGbmX22DQX
Wr+S8O6LP61i9RdAvFe72Gbrrg7Fgq621jCeBoR8JBZYA25IkFfUPGjASgc/
Op3t5CE59H9kOJmT62Yd8dErlbA/JCEdVGpEqBJgnIiTlhT1UDnE0lIloxij
c6FCZHwoBTsxiM86+VvBDfNADwxU3uASZkWYFXOLPcaz1ApcoEb7BQ7pZgjF
9AuMtCEE9GA5QiPtsZoL33I4od7Fo2vWkRwc/4oE5adNdfBOVi1VMUOnqyVx
ewUsRI79+XrDwN69Ivacqm5GjcBhCnuc9PbjNkaQP+rjdsKjAH60b8te/cf2
7wEsvPSLlb8GCfcLlCHZj+xW4JeK9CG0Y5Grzgs9idTHd3LzvCFAmcQHgCjG
4japII5ytPNURopEUhgQdUhTU3g9iIzqtwH9KLhSmp+6VKp2H9bV8IlSvna5
3r9G1YmHs5JFl1Jr0i7Kimy5SpMllcxvslOuFNtIigPDQmW6eB8zsDxTSTJE
4J6f1t9Pv2a5T+6CuUr9aRbO4L2r7dEGpPMKC7pi1CaK2ODPOd6lgXINlpgu
dVTj1RL/OiinudLuse9h+4Cyra0uFzPY86GVvhzHg40QabIT5hBJi0uZ4sDa
P9VGj0OZj0TXLjol5SK0US3hIAoMbld5FSJ0fsSQlyYiIPm9mVV825N13xMT
EFY23ZImEh24kzN7rubm0D05qET2/dsu7BXIu0MLUpsbpphyS2leE13xYf+q
AmeKXYj9sLV7KiO9w6pAHoMYPYJWdqjukAUgDsakOhMG0dUnLXRm9yUw2Gk5
zDkyCdaSnYbRYQ/gWmur1Ys7NMIg3kphQqDG2r4FLxKKh4z8jigiw2dzeuYy
9hNhO6uYuq0hXpws5JNJf0KTjxz0FhUyKcRjps9D/F0KOxV9XYSrpBg0osJR
ZhsuPpuc19rDUKfL/IFgo6xCABIBfSBBx0oGxesyHeas87yRvID1Wj3e8r2F
BOMpO5DNot6bs4HEJGZFdCmGHwKem49CC66DiTdPX8o9DuQrV+Upv6s97g/Z
Oz1MDM9baiXsS+IKQnzYo5xFBq4FFtNRpUvIlF3mNabd4QnRhwKyQIefHikN
+FLUS6AW6uzR/l4HH0owd6llB2xjMCJaBgRfeoYMM6+CrqdeptLsGTGbV4Pk
xkaUbQOeMBImG07Mz50EkvhLE+L0Y6IuY3kZIL0ms0Ron+AbBRJ9dUQ65nbI
2oOnR8KwfApu7v8OziOfRclme35djyDh4yi/kQMNXx8wNmd05d3GBYCQHHX9
3jUnzJSdPrOowJttxUYek+sTRWTH6MshVhG9z6doFxembIpQXfHvNA/DT/tk
XFcP/JsA8E9i+bzNxVTIG1NKC/sQJ4lFL3zD0ibisFeU/Ync3oplDdQ7jcuT
Y/DFajAFlg2JxWwWitlq/4BmYwoj4WZ5duzWyZaY60s/KRhfSI56BdLYbVyV
poJ2QGpSrafnp8nzIJ62HamjH0LsBg/iq9p3zU+3Adeqv2HREJOYWZTXsvvj
5WZrwttiRbEGJMSjPQXlrnP9h4CmxDB9v+2Lw/gmjbHkF3Wj51Q4fPR2sqrL
vnq6Y9IC0+CzMoAQdDYup1o3JJMNfImAOUPerq2PLtpEpGADZidGvi/9ZV15
vMjex/PeOGm/BenDW77XqC4A7rrhTfjGigiwD9hhI5w/rMshhgFrQBgSL3vn
cq0UjSzPVyCv7ZkKiH7vElLIW7A69Buq/Izl2DKUsPB3fVBe7pB292rPsyw4
tyh1XKwb1N4F6HwFXtTOUBNdsGz2WVWp1GJb4WBedn5OxxYHwkTRtWsGaMLN
d6g3ghQ1fUTbR1cB0WzX6f49EMtIloo6Im2gAM8LoRERvWlMB3nEV2qRF/lv
dZIvSSpf7bk+n3oxh8DjDMt5VziIQxzOfGkz+fTGtNgy2AAACi/BdDU09oc9
bUdZWBx0xCx9uHOr3G1pmz+uA5mSwCZ8qX++G9mo+Rz4SGa0FpLpjZzEZco6
MgR9bCubkN3/hO3HRUzzBjHlRtowyW+J9mqeCr6UjSdyoj5hE+V3gCQiKio+
zUQKa6XCBJavuJtUKFFX3+4ibbgAom3/q6QGcHngRynt7jf2sWkGE5A8XeXz
/Trwyh2hkHIrhJgtb/GtJA4PmeOxromXL0rvoYMYT2bt+LoTLUyVKh2Ehjzr
774JgebmadUxf1ScSL56wNEn+JnpcAR2lrJaNIHMqcVj0gwThqKhbNjycgof
Rxu+PYyBXLyKnbn5tiBxozAtwb7Kyqz4UEIllPR07qARxjNckut9IlAbCAzk
rVUROruv73oxOLZcqeXtJu4Q9RXOJFXBPbQVorUHES+dxXudvSw8LqWvHP3g
4akTJ0xm8rdIPH4QJCS7+ggGEzLytAzeV3MO8+bAEd59SGJEsBB7atpxdQf9
FtjUQ0B4owUtweidXtyROSIQI/qQPYHFRwkeTK73b1vqK9IUQJoFPggZ3pwX
umygD46vQcsvjgsk0gNUZe3zdKut5V2Ifb+6laAMqT8oCTxzU/BT4TDwOvzz
D7sQOzqm/KvAJxJOClFQdWaswdi2md3pPeYjTZ+S0ECjhlUW/xWJnvpuvx9s
Zg58B9eAHujYhfBKG6WGPTDSET7n1O7XYb6X0EuPQXW2KTdJ0PDEfVqQAQCg
Oigy1TVh5lVZt/TQTU2PDl3l5St6N1Bj73l3RhaQTskRCJZ239MYYhxMqH9h
5fNFFNbvZIHpIm4B0a4HCSh51LX4y56ffZN/h8GDe5aUUIRiSiv8bRUQP2g2
wzj54jekyTH6ul4sgqgQXkTSUMu/IlSIK2D03rWRUreYoFE1CIWNUNzaZIgV
AAtcVcdNVJFegenxV3HKyD4SvTWbPuN5J+OU+I3tKFTrTqwaWbKtn7WYENNv
zqLSsIhDPwJsAETn6FbZIy3QfR6UnixlHIDe8EyAMSBq9YxLcthxkRdp2/As
wjxkqaboLFSZQlWEifjo2gZi5hKWuxjb7kJOz7Dh0PedihyWRPqQOlHUic99
V4U24ubZewvxTN8OSoqEFnVak7Pxhr72NFcibfwUuRkCLbrt3vVste/stCED
r2HisY0DBJp7rfM+aa+3G/N9FRCNJd0BtYvKOOSlBS4JJRY6rod5getSCUX2
GDfA887UJEFz0WXoDAd8oJS6TqSenE7c5qMXTEcq6x6JziP0zCMh8tDdkNz2
ufPSXpREibfzUs8C0ajwrhvcKEU7Odb20ePQNZZ/AvMBBOpY+SsvjyP0Tlvm
yo9iJBWVjA5b8hRyEOcMpPPdhSWtL2W8kS7rw1LMUBcnPV9kIf7sfzfh4/KO
B3rOcB75R6ot4hgO0x8P5+qAjTvLsq83MH/0TOoE6nwos2V4pa2oW/k5NkNZ
2WpRBmTn8APRwoO9TdiC414norABEw/D41DHyFrTbcYISd4HTRsm+LeBKoEV
LdbZWniltPWzBZilEEzDzVNamSFkM4e8PMRnddyT1fjjXsOQ70FCvJjPDtOY
1Fx3J8gKf58GHGFjA/8fGL48K392Tdg0UyqmWDpPAxMgUj0THgC+/eLgwJ2y
/rhvUdIqUyfzAJHckRMrXL/GILFC2WJ46tFpf9fd5bCHFUNkIeUXQ/QRGnTg
qAkche3GhAnnZYAmrS0QdmxuOuufFwhln2bP7aIMlXuKhy2c5K2JBXb6f7Hv
XKGHOhCG++oeIQkddrKoZdS9MnCcqYtqdsijWKE0q4v1SMNYKR8YYlkLFkQZ
MuTakufdfj71we8EV8LsVvcI7bvQHEWUlWKcc14csXWq06xJ31QVH5EspIvV
QDcFtYyTaqcxr6nd9WFSo7bPcN4A5wKloGUDhB3ac4VHtlnZ+7Ex4e2urtUg
HzKlzELXHdiZYfNr7VMnfNP1DVzbC2SidmWmOp5/7kPyxbdG1NIQjjyP8S5Y
R8/etr3M31dH4cQ8CTl4D2mZAKUpsfsrBn001OF96E2rhhSL0ngx248QRfQG
oyGr4bYfi1saetMWYQ298wD7I3Bmoj+dt45x7zJ2iULZqu0sTxc417KsX8jl
pNWQDDZpAPotCdK6atcc9KMgwsm248+ieanf3wfUaBQduvcyC3wSyyrNkvc2
I+P2vR0GnDxlJ5ZCyFKIB34A0JPbtW7TpxNvAJXpxFczZLdiq0xGxsd+2vPt
iYnMQYNhHHtCjc9EkSfFMRXyNZExee4sfgrYsYC7paJGTExpOO+K1qCU8TBR
q9JFN8Y2PWMJHTlbUFy3gwsTEV5HvudV+RygmiJsn427b/vGJGEpn36G8+up
L7Gjs5CLYdTjWwQCv9CNdnCwmMrU2Nw5KBvhG36RFSnZ5pZBi9HEEQT19Rk/
89iCqvItrtMOqHf4eRYdRNHwJSWUMmcpMLN6Z8pA+rJr5IksLQCFPoGlOL4j
q0yUzWEBzC6zp0AGP382X8dvDqao7Dg8BvCnqkMArhn4fXRm9dU75Gz3fhwj
ayhpWVgEQRDzOF5sMRfs2e8I6C7/4FxK16bqt3YFxL+Xl3T3SO6A22eY6nTx
rmNVOn4nuLK7JdqQ3zAkuyM/5hDSWscmKuzJse3w+CO6vQwUzgHEe0uQgqHu
9sq3ic8uks0qQ3bPm/yYiZ5S9ptT8w5Xpx8A7MbopHwpt6S+moCBmBN4Tu7u
t04F2XnH0DLWSOkFpp0HukAdGhEQNqeeEfKLqFaekNHWtdg/jGWJMC53UJnh
q7RfrJO+eGEaDCk+P6RIJvyCcjM9Ls1ZT8KjvOIHXtRZNFnjQ42n84k/ebRQ
O+OorP4vpxwhadXM/Gfaos1R7OBpM3+r3Yn0uZ/cdEQErac5J1Z70dW7rLFa
AvuhOooyjGMx3A7Nmio2NeWq1K1sv07pTQQgajQBqNjG2ekuEHYQcMfqjNdK
ODGomwrIh2aBfE182vWuciq4y0GKCyjz5gto0pkvK9NbOSrDOc/UOJLOaTi5
csxHkKYijJ1ncO29mjMcTKg1Y0/I7lHtKs0T54aSxoCqC9jKys/ozQcG8EGl
w9y/1DQhVxW5PYLUB3Wy01yDmtCjAepz/zW/yUf+qzrp5VC9kfzGcsW5Gche
+UMfMCJW8q5kwSqkKisZtyMG+nXD42ZfrVXC2cNj+LNGKA1sTBtkp/9tN0mm
JtBQiRkD/Cg/DKPFqPFmQtsUy2kmufSl2oKahcFM/u5titNwiWWB0d/P6bJR
5bjZlYgRhKA5oK41pdScJJMTqKsR/7rxNJ64uod+bxGMgxRS00BQ6aJ8j2Zh
k8drKbRXUL4chBCVongOnmAG5tHaxsrniyvDMxw/uhhB/21St6k+Tx8TEROU
ho4qcnwliaMr6HgHQ6CoOIpdVwTZ1HrEAZO1Xm8FZXrLp9lsv5ooiFrMwnAD
n4EA6Hty3Gj3qriIJysrNZVASoQdAOFiq1h7aYdU4tzFXV/z1adnkYyB/Kfj
ryvNk5VvYFNbEn0g1A8bk5rNb4AFPs330Agf1nr4q4tYyhf/klSgoKcaR9io
1vxc7I5E8OH6BTBkD50vk9RpvZJeH1o8rTu2Kmf5qCUrLbkhkF/VCEpvOFwR
Yad0n8MVYyaZVH88LK+ePNKnjKTsOS5wKbBJ1OBn6tvyvDDnpuJ6n+J6/eki
gebwKXpsOja+6VzXyJPWlnkRg4DdRUKqz6Mnl13VOZRQ8d2qTTw8Di3ZNF1+
9AgCykoi1MlKXBR2PPWCOBvz4tl4OIeZJD8B7vb/7CI6ccaS2ox3+scg9bI0
IMBnYNqX7HVHh5/hazdxVq3hL9JSU1bLTorBBJ9hLhiokhe8HOTvI3YOx389
OHmlkHt0wCaZcKrDvNIakIR4lvSE7DSknyQFihKNR96wVwDBoozuJfyBPER9
hBd7PR0uESKogvx/a3tNmJosmKrmSYRgBy5ms4GPbu7JTQQPH10qtuDQ6Jph
mCaY6zC9C57zi3EpCLTDXSk5vb2q8hn6WOQdIlDgLhYLxPpXArXQlsaHCzBz
DaCGsdh/dBlu3fFylP2YuOrOmRT8wQchFddR4weYl6b5KhonnGW0t4Wjel8u
JAJKoY8fl2Q0XjnLA/wgsoKKEv70EbpChLJ8WZu1H9D2GFaBSOJmQq2BJucX
lgMVy363P/PnaCHwQPRa2mOSkJTI1aG4AbOJCDn8jvQe8APPNgIXHTLtxuQG
v5qtTkv2RjVYZ51v31BHDPgzG6wWgZOW1SP23Q+CbcSrKeccf23CT271f9MY
5w09K5YRqsMi6ZnUdhUyOUf2AX7cxByHcdgaxyzbVQYZ6IKLs3SqQBf6NnN+
4ErFZrYTumu8NxXV8TWPR1mLkBcf6PfRxGywsMp77gZfjOil+GU9mNZjHsVl
eSFLhsF69k1VHOrAv2xHrV8eSicXFzbTpu7jWs40RanKMccj+3/Nw4Lk5XXW
FJKDsFydvqslIXFxyEE8LWnYv6e4XIpPiTiBqruc/9hicVhEfjwinynvBN/v
9ex6E9HmdcXwNPAQRvMjFywYTexJwWlYbFLdle0F2kUTjTzFbTHS76orwga4
kZXf1xqeUDvHClzkwZa1LFqkzwY/vzeTI9Mv3VbNmTyVpKkBeA//1c9nZXPT
OgDv2LX1m6+gsI41p3rjqmfvQEIZPmH7IKw0Atfj44hDfa0/+dqGyIyo7jTy
Z1szy0mEJ/3lina81yT6eHvQm1jwEvGicWkQXOyNphD/jq6G0YQzfxqJn9fr
3lp1MmzLpW+1fKCh9YaMpU4f6eMNhD8O1LN78dmrG5N3V4isQbqd+BiEzcwF
JJQybtJqjqaJlnPklAkCbe1U7PDmvoMiNmi/IrhmCOZWovbNRXR13WGdIGQ/
fU64QV88luWXBhG71rvzYWX/mKsG6BQNsnLuPnt4demuoMxEFi41uPrOEXN1
ndqRi0KVUnk5S2uNsQqfJ3t6jBICkVE/PQdrE548dnrR4MDOHwd9rrgTJJRE
IBRaGfHIOyJwjbBMP3zizusZ0eIb+ipQq1g4XuRRgHFPf7ThNqaNHt6i3pNy
ZAcxZOJZo9xsB6zIJVPmLRuBzCU9YCBOVaCWx6kn134XFBiHkN1J2yrr8rLb
n13e7If3H9b+TyFJWe3LzwUu77SrE+kMd5EAu47wrQDj+BeJwK1RxJzKQWKk
1xJLbi+cocjqlY6N9kfL2tdcgAb8GeHeKPusRUTPiFTk8Rm/qaslM0uq3y1X
rfQhn5NuSDvZd9ksHmsKgD7v/ze1O3Rq9gzHHhtVndQtt+D0Dr4GlHyWKWMM
ZA4BjkMBi2WLodoo69kANFyM0tLkmbUUensslAG5kG0H78e+vt9FOHwVzNO9
CHh8S190E4Quj2Hr//nf6C4qhpIVi67f2zgS6RtRWFhGhoGk5Ok2VH+w/+2d
1korfBhokSzEQK015jyjoWb1qJo5UGPhQIslNk6lRIMUMxTFC1+DkDpFxo1d
DTdC9S2LqjR+r1SDqcQkoGSr98+TbwsPO+At3Ad+pSmRV6QJkQdEFZ1m8CQF
F0YKC0oa7rgH/9Uy22E4EjQYOHe4sHAaw6Xph3jUkzrsjRv7QcVOJGGDQsVv
fL3LIW1Bo/0gaZNECEnRVQwWIcdCRu0btAhOxdAEjW6WzTiAx6Hn5QhmZN5S
j64Sh118uhAXR7OWCSVVaNeoAFLuWS/0mbI6WAPH7+taHfuzuMuRajvqzj4j
K6cJZT1D5nMqQKXEWmRmMusvw7SziiZ1J6WLCV39WIHSxTGvpxaJlmfvFeGF
KelTCaBmwZLrYSjjCo9Wa6lwLUFUl9h90oF0k50pOLkFT6avpVWCayYhpMk7
smDcfPOzKT2m8RcmZrUlOyM3D/QU06mNzoPtwDylDLpdWBe+IE3ZZ9VSUB3C
iFIOSUEx04PUnLklr6ukc3m0bWlpH4nFMz8nFZ8dngob2lHxJUfXf1LweoIu
52HUxGGmozJhOUW4eP5mZsCta3Yt31FC7SZHq94HhN8XMdRfMTcJj1hCFqAJ
l9nCpddx39XJRtE4VWXFaL4pCGvGGHhVoU4FV54/QvdQg96MYXT5f8b6qQgz
bIWjP1Iib5ao+UlMynuRduYqBu5cp8LPpeXjUf1U+i3fyXpdgGsTS1fY8RZc
l5WnOR2amZJ3j8DobFi/ZLkJERsU/wq0NVbvzPw6u134nWbnC3V8+2Ssq3cT
NNnw2brKCpBQtZPQYjLgE8T3ixZxdLoZ/YnZe3cPDYtJWeWVjYWmde4uGHOf
8jIMrsda6syZAHfF5hOUsjm6QHrQhViYSxlJmyyFA+07vaxAjci1fhAc+EjB
IO/0THvJX3jBOMngIGztNOhe5nIYKh/jAqf84MdticvJJNH1CHo3/vZ95NHz
fml/sQu2AtKHqXD6dBSEmpgQ1ohvpcJLyE8EipUOwnLwGeQ7VmTUxg/ToyBd
Iq/Xua9ESvVvnDX7UDXOPitMF4TWx904kD1TXIIuw+gRkUtObbMRlum8rcEY
OKFgwrnHTsjsB7S7y9WPWkCmOzeQEVRt/dYjErHW95bmqPLTFuiC0mMjRn8o
8cJiD6uLRzBqUo+kTyAhd5LF02xXQPq8Ah7h15hLtUXEHPtBi5MK8gk8HPo6
OOvajMDJ4WqRbTP6f8jF562KKZyGL9PIwntRiMAeSoRaJ7x5WL0SGErGfcaV
GxS/yGsX2/eRDINfDNNyYn1NJZdqVkUDkUuoMVFUAy7dvJfAygdA3iRpVZyE
VcuhS1+gO1OC3C6HE15KPozgFrkp7tQB9/TuGlfI1TwJiphnIUD0C3EExGhB
H7KCvzc3wy4JQIs/nOIVqouYaNau8stOHKbc1k1303pvDebEmjMIpLswL7B0
gR7Ro5qwsPDfsOXx1HUBVsOxrUcwom5TFq29AnlRxhgaVgIsfLbdgqJ8h05n
C6ljgYNzsOkhoQs1JP249igL3yZ79b4Lxujur3qYKt7xzD3dj8BrIiKXOsIF
IRb+hyDtj+OiA3wg1YpMHtNJg5+tN0YI5+CL8N/SBdMctf80sJxFcoK6vG2I
q8X5AwfKr+9azs9pGr3fOwjMpP2SZ+rj+GqOOQETbntFYHTiaXh86H/e3efM
+nLVgtRCIQfxWdwAYI4m+sB6GgreWCLj9DtpSAlkhw1N/g6dMAeEuz6Pr7Oz
pGzUDW0cMWhaHpoEjH9dlP9wJpNGRsrLs1/YDa8139K6BBoeslpvbl3Atpzr
IDSSrvNlXzgXeh7w32c7r1oMNdK+yHR7gmPSKukuO9rfypX+BWHyZ+HuL/gT
pTftMaWma7gWxhgosvS9uWaXVH6mqOOrO+AN4n8kyJz2x4Fv0c0AjmQnola3
CbUVGRdka+XQV5ZK058ScSazpPBIC3uNbsDRAqqzh4fYrgXJFJuZX2VB9xbg
6n1NJec6guOFWfpXqVc86bMBryWKTm4PSjQHpEIussgJwXavOVff5AKl7wzi
lEoYUAr5MXnIae5l4ljBXnwt9nJFjhScOBI2iVmqA1s0sjz9OwyUbudK07wb
eRCgvYFdevEOtlJRnBqGxg/9juZsOqcfQIRbGtyqdHUFp+6rth4J44xJS9Ei
lY3dwpH5rNp76jR4EAlUdzp3PXzOBkLnz+csiYynK18LhxpZMHSzNozz/DJ0
nWm/E5+19OEoqyp2SSMK2UzGbVxv83U8JK7X58+3piJ+TT45YPA8jX/sM0Yu
MT7JpgEVg1BnHomnjmeQk3ICeE/Dd3FsN8qoMEGQSNzwPB2IpoYe50BbLFKA
+RlvhuAx6PE1cgAbQ4xXj0o1DK+Qe1EVzhWSvdr0GCvqIz3p7kNLIUxS6PKh
B9Q07LyFU1xfVgunHu0BT+dSN42Gj6MTYJR7d5yMAnS453YoGtNJuDPf32rq
rqUBoIO+/z9DB7EtT0msTG4Y1orkXCLaVTSwji3w0uJHYpctwG9qGNC3+HGR
KGCw+G55yBODfUupsA2tQVUNfbRR9F/+Sewp0R/mVh41H+nOnKJNcvJKeVPQ
DkkiJtU4fPnyTCxnqSJt5hvcEHhzL49sNudqVapUOix8+H3Ny+FNdCtt3rT8
i6rMzJIGFUVHP5V0NjAPIn254wwY3f1voNHzrylBSkTc64KzqL2qXPT11J82
dmzecfx2yeY6cJCNZ80cGkCtaWSRPb23AyIkMh/5XJJVjFJ7kkQj5+fdEpE3
N96fsEk+Z2yY2wggyFBgbE95WVTiXYXNlclvzvC9f8MkHEcJJQl/rttM5bpu
vneJDfHLLw0CO6lPhGOjxNMaTszJB5CwqjVZl1W4CrsdZts+Zm1T14iO3a35
0l0wo6LPIlrjraIx+SPBachatjMXrXoawjQrJ0Vs9o/VvWxBuyV44Zev7ovr
EZHNioCt/zoFzkpiTX4rHaJGJNdCTCSPcfGjg0P0y4RBbg7ojLqV5weCfbOe
OREJI1qkwndUbMB+xd0lJU+yZuoOhen/8T90LsL04+zdwGzU0Xs67GUconhq
574IZCJCGWaImRKywUgpPQe1Y4OOZspDr3eppaVdypZNZ8tzJUR+RlKx8lYX
b8o56NzpKJxDIukw2UOKLdLgXwOhohTyd617zXP4q9XSU7+58l3iSqPLrdjD
yU5FKPMuzRro1mJpT++SnqmkNK0v9RApf4WkCMlsPTZnno+6XRx8s9HLL1JY
stWEIWLM6E3SCEbSPqcfPiNQhn1eeHERzGYIjAbD6LKA8yVyTJtlNnbUCnXc
j7y/ZOgshuYy0AGy+Xm3SRZb3rZrM9xJYD9eNqVgeF1XHW3b4iRr4A3T8Iw6
XA5+qpLEs1ZQwlOHB4qexa5Mr8aS3jXR/DtVyVrrLmet+OSLJs2CTFAv/gXV
K3R7RiViOFGi/x1P6OMTdIJF9kGsQLY3o19hic9+XJ4IC+31DU5uQ6S/gOuo
uZ3JYXDjgiAsU6RAp4Sw4THhaFsMaHXave6BAmq0479bxqN48CY1jlYjdqbg
c72iER67Mx7ELqd/Rx8L8t0IKG5CzCuhej/M64p4RzRHAKM2nnQ+LnxGCshV
2Ad7tLk2oy7N8S/e8vLKboNDnijvR/Z3xpwEY7ZqV0Lu3fazbGC4Qf9PkDnC
nikJJ0nCXpFOhYGZx7jwU8qI0ISMt5mj0VoakEqmPasQp9Ej9HmAGsJciGth
XqRvc74zrHhMJcs95owrZAQVyygQjK7pSJPaDBTTEOtZgDGxYUqys+YHhFc4
B/RfzU62KwU6Nv3bIojcrpJ9cPkHuaTMY8o/wqqUu93yWMg/mxFqfAnnQLSW
UQjNas1asjUVDkYmNVUrycskJb5IBtDvmmpqsGV1zk9xvJU2HwXWFpy6mZ/2
QRjFomBV0+g3g31l/eVbCTJAum5Skja8lYNYC4gI3Do/Dr9WyIbt9bGrv23s
Zip1ICbzifDDOVduzt9yawWOBHZ9W5/yfV+ht1MBABRlwkAus8F9EH4DunwJ
gJdabl3sgiXnNGl3NXiW2eYcxtTk3ZFGW1KKSS+qmsL4oUoHBsaq2kldgZFt
nFW+H5tjRRwT4cPuewsdZ99G418J/xvXC4WeTPXGJBE7IBvHxUxe1AEHunAw
cITnIekTbGQyS4+yz0hLkyvJTH6wKVek2u0kMacmSgi4AAXOQF950mOFcklm
IBi5AQzctZjAJSaHDM7yZ42tE5H5nOUOThcK/HQPykBGCDJhULV7GiFSKIRo
Q3jpmG/ugtokaXzLx4unXwY1rMAUIc7+PsgOB0hgEiPmmyyS1U5luOJlkYbt
rtG+KzTld+z1tkTRWECNs1HiidSHzJRn+7kA+DXYjlHTHlv3yr14JL9JTAM/
dbZrpzCBKH6epHZrtzvy7eU5AJpYWWNRV9jDGQaB4p7bxf82KuLDsTwO4D/q
Gb8OirrPf8Jsmc+w6csHWbebEmZZ1OlF/UonYiIRXuKHpmICIyNSmmSZICkg
3Z9efmr6LHZbuRcYQNHES3v98yqXb0n+0prGCDgizaAAIcJxLesZQEFElkdX
GpgWQvek89adlayhmf3XPscbLE+JysdZWEGeSlRa2iRIe9Wld6PKZfVFR1gg
qMXLnIh+2DHCc/pcpmhBpu9mhFlcRwVW0jq/7hKr1SYP6UyJqlD7sxGqGoqa
HEd4SVb3DmjKHhbPOtxXj3dsQtjIVasR4nZsxUhRGzP4/08NhyFGbM02XKn6
udZzU9XN9oPCyH5weJEoRD+hgfKK9IZAFPY5OUmrrLMWjYyfE/5hVNn8vn6D
CVeK8fOPeUvr7z4wqQn9pfGzukwTGloNhbhfL5Z4SyVWhqjgby8EikC6OL2P
iqgHxFMpqppa3aHlPo+bJ75XMt3FW3c0CM9MkHxVUQ2e0Qxd2UUpbg3Zs/0M
GfuTx4y6wrV05EcA6r9D11SfQre/NR316aod/Lecnk2Jff9w1NcA9kVLpVdX
6Y9T2IpO3ZMIgPdGfOZY9j04zTeQIQ8/x1ebnB9X1K6hE05uutWEo+veCnyp
P+9aDH1FJHfTSYt+9uWx6a2j3r9/S+s5FRZBEwxNT6RJEZKu7pawHOR3umor
g4BkbsSIJXY0xJEpEK5ateA1BnFfAz8phusePEp5xRDIkdILMA/+krTMZhJg
7go6FDZT6k8n/IiOEFOr39+oqkXMNPD3nktrsi7vBDLZsxNMM+HNLXVfSqHi
jUd893v25GetXTS4vuNpA72rkzfHDUF0yahICyQN2r3mK8AEvwxLAxApj2JG
oCnngLlg1AzXDrbf8oKxih+nn5ENuJ+rFXgnS+IFT0mtspmiZclQqzGwuzTv
0kvbcyU4UX6byatTR7G5huoe2hq7eY4KqpJl2EVvP2eOMbQpfmR/Deh5IKXP
0X7553SVpaVWkS8Kb768FXhIjt69R+QCFuNnBIhTLG+wKfHGF9sYwflFGam8
kt6ZvDA/1IJJuT1NCKrEDqS6c2kODeUwiE9AkPO4pN3j1iUNftheqanxQYMF
1hmKG2yxgDMuQFaT/afPw/KyCi6sgKfJX5WGgEpGLiTnah73obuEd4uWqBoJ
m9wjhriwV7qI22d4JnhOaXPo7jKdaYxsMEm/RBFXnSZIo+o2fGk7pt9MbV8k
gqV4NzxiHH+LgL7gLzYD8Jn41AplzbfuhkQar88BplaGudHWkLI+fO2cQDEr
LY+zSj0jK9C5PmVSm5+iVMml17N9qpDABJzgVn6iiQ1Ww94qYBDYLxO9iI1S
0IYYSrXIXjFkqoeJa2b5TmOZm4o60jMeJ84obHD9ec6nK7/L+tgF9VHxZ/5M
cGJLL3PajSFiayJO2VUKXoLrzFoCn0NgN6+VxYKvwWau1YK7jyu7hdBWiMpd
A1b6kG7XXGS2wBh1F2Hnf3zWW97JYhou43yXoNwkStmCBVddQLWCuYqBpUWs
Zc0xuxPq1Cz0LlHJvpOqLnHaGuVvNbhcH+q6xSF+KOasovcUjWsTZMMyU3n7
M+4LnVuqV0F8yBjH32E1S4zfOMAORwfYtgskbj3HKJyQ0QPuQsCeuGWUmjoE
o5CMOTzXh+ebMW+EgiGPLXo3ZTdEmaG46OOJobaoYYlnjYzakYvLuEMA8I+t
SJZIxKsgwQPGly5tEyMpfc2E9Hj3XHn8ZrMY45qPYnt09uXYnM5KmLMeuUCZ
7JQ6EfNdhCBbIDlsMSNDA0HCFTcOOxa5MJkVQbjTx9J0ZH+KDHtpnmgMohGG
l3I8c/Cxg0eGx0/ij99TcwaV8wh9nxVPzDkEBOsf+j4ICYjVWPbt5Y3N105P
zsbxO6tdUmh4KU1HK0dkDFSEbdhB8p2GER/mDiA4Khyxm3Azn/nSwSApler0
EhM5AqADz0mZ36V0UaBF3dYjz+ZPi2/fRAHcj5lksx9/8voCuLylKyBjXMjI
t/f0h3J/SDv7vxmepCtxz4tHlMd1g7U3PoT7xqMocTh4AMPlAqN/54fRsd4L
hB/u1fMKDRYOsV3G+AcXYe1PNmuuUMuEoW/DpfBfVFjE2XVXh8+JB+xuZEZm
aeuImjivWBMjgn3woxUKe9fQFEAel/0DreuudfQCg1n8d6+fLvF1VbiDhEOE
bbAXlnK56zmmTO5ozE31YW+pE9JPwXr5mAjJWGzQgYbF9HIGIJv7s3ZUaFSr
RuzofW2J2Fesbjsmo1AG4nFXOretIPBNioTMw0xTzcxSS6EiGpmb6U/9/kX5
BBjiXR+a4z0wH0XGIL7O2i+XWkvXs0mqORyjNWpS1Znp+kE066s/kD5BIEQz
xJJHIlYDfBZLUWFSaWYJX/pBv6i4QyQ6cO9XJrlnmctHMemYi57GEKjrrjdl
XwVCw0+Yv3y66MkCyzRgKz8tbhM0HklS5YUU5EIuyIT9ddcCc7HcnxiokcMy
8a1YjNaBFqnPG/K8LqUTu9n9xv7kETfsyXBMiHg5E5kxWBTnV+9thdkyVLq+
iKXfERcBDjfygVauRJvCMCpiUfAKGVrdvufVl7EbBSp0rKQTU++1vXaihIpr
/z5SY7fsW3+TGoR5QtXkHTfwxFMGSkgIAe/thujBB7ITrYxSgWMTqm1PI3is
8aEB8zHwQMLHbYDBJEV6XiTKQhnyfxWmflQVr6/DcJNNC5wxiuaWkbpQw8Hs
IZby90wwj1grICkW8bLrXzBBkdcFKSadNX8zfTpSri00rdzx/h4o3Zfa5OV/
6CeuuI8M6WxClT7jBMlZo5mMNLVygp264w38BHmjQwYMwUttj8ze8qgIoy9w
Hzaps0ae7Oijns3HE76fXAMhRZyUNezeL13IN3Lqfn+pdhxcOQgm+tlgzvYj
T35036AwKAo+9VkJz4HEiGA59nVC1VkClU99tci7+YGmKkmTCKjgE9C12wOD
Q09lchTiJ7lqiNk54Ya5G55PkDANkZDx0kPCdCyW1SdQZPxoqofdIR+xKx1c
JypYuRy3+T5mvuWUOlpNaE1XXb1rzP6as34oWSEcfn/yvuTx8t6hf+xL5nHd
Pgs2G4GRZN4+cXck/ngO74BtiW3rl7b3oUWBI0HdhYyQk0URWnTM+kgS7l5E
8BXXpI6959QWINuIIiZbte3P8V65n0raynFtHfm2RfqmQJX73a6D4bLzAKjt
Lf63biAaonMTy6heHusHW6faaChDbZr3i1B4EiDDY8e02arAt4BbB14fzJRI
2jmM5UZITT0PFee0EHqHee9sNLhdyYWsSLZEHJzGSzbM8Aa6agzY4nx2GIDW
R6/FVuvnwp4kAgyoTzBCNRDYADIk+BPznKBRFBiUhjdIFDucGveew5RnzIjs
L1ppZkSQWMbw3jDzEf12yId88xSVHBa5wTPkOTUE+wOGx8u/fj9vs6N4zIj2
L6XS+JqT4h1pvhl09dSGRo5s82p5/W+A0uEkQVNTnKeaBHc5s0jRpnwZ8fsR
gE63gcfHqz5YwfJSAkQug2ism4Bmg+HL5l9hKBmVq26nKJ7h41fdfFdlT9/w
mhwJGM6grgDKY592w3Y3yEPlrEo70778OGo5YFObKpNjyS1LGA0w3czBUrZD
Zw1Bki6Q3CRwWxAuKvg5oith76H9Ds2NNJIrdc+42FsBy2t4wgLFBTJSzsEy
J25+e+YHZX8DioHUiq3gBJEAejzSNtqdN5uTQqCIKC3W7kjfrt2bw1EyZ5oA
EEX/3CqUF7oYfuaQ7ND/+l6vkbiSRZt5IeN8PIviMZ5Lwbt4ov0XLIQl7/bP
5xAsEPmM6MeyFRFPQC6R2Iy4Y3+ukkLTIq/zux8++GC3tpEdlI8DjKGbzf86
LdrIpdWnNJ8kC0+R+yNydnmNJjgyWkXuLSGkNwqUkSXsD2oPx1tWodJyx2My
thCKaMd/D3g0UC77Zw0uS7cALMyWF22DoOkhHEQTflyrGQvSEuDZBhHBryy9
BG1zBZP6f3ornoyxFH4bN89VAewZm8ctNoKuL7sF2j4SdZ2YNH3yq82ScQl/
C276cBaW6GEV7Z+O3gqbx0YsdKgvPYiaVk7UoOH9SW/5gcBbXWe7ILVi1NEE
SrYHm650RacYJ9c7mCn6JzBRj78K0LAQMVRp+M2BtwaOdCNILbDdI+fqACOt
lYQx6sU8xJrPBZOXhoH9am3khi3xDqlt760v/qvjdn+007LhTNrprPTz9ON/
abOsljSagSnQd3w2qdxTVSDHfpj5nYUS4cMFfBkjVJn1e2uU6fmS7ngwKypv
SmA2lHciSGuDQxprUGHaua3NQdSMSrJa1J3sdYwY6WRFqStGFnQfVBzSxB5n
8P4XEtBhDdyb3zw6682wh44WdfNyRXVKoLCEUs3BXjD737uKSYX2GkJ0j+Of
EYBJkemB8BNtLAoXg+4BgjT6Jfz4hw/3ToZM2ZY3RWYjZtfrv6mdxELJeg4V
lG1kgt9nmddcQkQ9ExNO7UJiE7wB7jg9quBwBvNwiNHXxmjE1NUQdFoHmtP9
SzKCxHiQDSxLhl4oKcuiJ/ym4W5mhg5R5X1iEdKCpYMNqUQiQuuGWPtqf7T+
nRkYVjkY2WmxYoCGIT8qrLp7iwKFsu6oQCDtw+Wqw5Mm7s5zLZyVi11AN++q
gGGfUNweRztMwE97X1YH5zE1hxP6U7vmnQaH+sBSj693qrtsBBgyeyqPfSI+
rW7oi/dIFAMVP7zL4S7hFr56e2/y1z1Woq78xdwZnShwYe08W5Y1pa9Tm7b5
ns7G5sTDURFaE38NAyUAkilUWeptX8D+6THuvqAP7XBFM1ib99dKDCo5IA/V
ODFqRj6J8ATYPM/VQTOqzItrIT8lr/NC5gFPJUwHxz+8ZZ3qBjAfdUIfmLZd
r/3urmAzwpsP0Dmi2Q5CnSyPiJnrp2i5pKeupr3XQQIuK/mZD6+0zcC8myZr
lVzfsjg7Q0Gmv1SvRiExeP4IKGVNLbh9Ew5DsqyALG83lUJtCD1zK2mQTMAV
jRReZvAr3couqlDl/5gJp5MTLBVkU9jpiI+hYCEVnjwWs4kaP001B1KjgM68
uPzuJ/KyJCh6Lzo3jQH43ykOEoaPAh8NRP1dlJYsogEYN0s6SIu7K6YMZLpS
mTUhal9ZZGrJJK2rQ4jsenjegGPKyGGMk/iFXWPvNkVZbhENG7uglBG9Pnda
vQUbApwkJgSIte0I6KOQDsW2lKVWt5jzhjknmzW7NEc3NXO1aKQxYOxkv6yK
oF5pQ4XSH3rK/wdJy/43Tt7O6l8u0AFoAlHVK/yNwvmC77K+PW6CwVHbw/X5
HlVnAY7+N8Vbh1zDwBZDDlI0gHt+0tWkI+ivBMQITwIV0L1xjva6B/5HiEvD
73t1kpcxAiFAaVcisXwSq7GoiM5iZWTyCeYyCv05CYdOpsFqPVo56zYQCSls
2gVOn7zLrpes66XJ2xYvphYpZwbb++S38EDdzLZbSOUhobLM+RYBYfMgcAy9
AyYn3UEFxIHjVNUDCN2a9H+kjxsP8K3ckckRrJI3KkguHZhUyiZhmEXDB22D
I/JgE20n4YA38zKz3zc7nz4ot9ldRmBaOeOj+eDgvGVDXL7yXnP1bjMms7no
6wX5H5Hj8CW4elS4jTFYcgUeKsUEu18pmcOo9psQjg/dV25kTj8hmCjmj5co
ks8EXBgD6vE/u6jzPDyKZ0PX527wKcFAGSz+uhRLmm4+ZfwfnOTtsBH1/3+e
QZG9aO1Ptga3M6pwVfqiEcl4ID0LurN7ujO/Uzt3irvp7oa/yXnKrkndzYVp
USHLbfUnN/uOAKey503wMWL2h8JmotWBTG5Mr+L/o28qu7aKFOYPfmxRcVoY
MHwpyKtDVOblSzJEVK/BqfZyuPsBOjprKTOpkCzayaKmBT6hqFVQUzp0KsRS
wN3EDCat9feoio7B9d7Je7r/09mt9i1Hdz9Wb2T0Kz5DtS2FiPsdBM9hymFB
NsERF8PeJJwgGUSvFgCoVvZVU1HyfPHI17BHgOxNCLPsQLLilglThsz/O5yB
G9lhZNHz/dmKVNg6jFatxB18beAfT6DaPbMG/X+PiUWDC5LnfwJtV0PxKVSf
D5Iq78jrf1ENbhzLmqqikEKx4i333lvACXJad+ceTQBcPlOYxXK1mxmwmfL+
N9IDWnLXz4ABjPwA+yr3nP7evH56XDYySRiBXR+1KjlbgDxXaxzLjyfkkRVl
QgcwaWL+ztAzEeSCjxVhQdYwgy2PIfrPxR0erwQZ6Mii9U/NORMJ13cfWRpw
1dWaSxfAOiMyth+nLcOH3Jw3kwflvFinNx2ak5mlSwQzHvPWuFITpVlFkTqT
09HFLeO26INlf4DAEGEVKF32nyuUwiJ7H3APJLlb7Xlxgg6vTltaE2cY3fnX
re8P9jLaWsrEBPgMwzAaZ4fJiaiGDr/v27HNlzSNoS8HG+x1eYyyK6ErhpN5
SHRYLUvlz+kZTpOZB5KD3brqHMWbkNF+ROkgEvaFlMl7JCnNnNRFpaEw0h8u
KynkISY6UqYCThH0iuejZtheYowArl8S6g3NzhRLMt9JEMi23C3Fr8G/k/LB
rkXnRownFOEdgB7uACocRFoTpKzcyg+GVn/sPQNAeUdyd3jBhkIuUcezSKN7
kZcuq4kD8chFjILXbILoS2BpO2mnSsfwAzU044xmjySIuGSADK/bNNCxcrSs
j5tSakZ7G2oxfDtHHyhsgyH2w7XffVDZUkgOf5aGiqlTCVREXJ1qPKF/szm4
QP/ukcbMoZvpEqaInVCBGeI5w7iQOyrCoHjXXUjNJ1WhzU/rSWs3nARsRboB
hxH4cIinIj6mB+8vHOv2dl+2OrJrYEZravev3I+MqIc+V3kLzC6RqBPIbRhN
Eruls696ychwf0ks01ZZVHeUfoeedvl8p/P63RHK1uNhPs47HJulMTUuncaj
zj3iL6l1b7xnXrRH8ZTXcrp8Be8K21Aw/jLZEmgf9TFRZUHgLOEBNNWkbkUS
kw2E+Pomb7e2BlPmdMFP/aJxqPMoXyiOacAflkTaJ/DXj9USG2bKo8ZikaGz
fZ5PKNLDgfelZuDK2kbQqYjixvF7NR5Hfraz0omakgqPOORDB6wVMbcqaeyH
MUz33Vq8nhEM6Aygim5Y/Rrtvi0ItVmp6YJ8WcDN/Udz6qiV8VSKUow3NU/e
QMRh9yGbrSA1s0bT13KZn1vvbyDKjl/1AiYxZW9jnV4i8HCrJXYP0Ctsffsv
88esYxJnKRkgyLlWf/zyBmE33WajGml2GKsfNhSXZjmI7X1xZphWZAa3tQrk
oYFNV6QsAapmvs7//gHtqSB6rv6bgtPwVrQo8rvs/7yoEQ0ifUDEVo+jpI68
OjxAn4VnLjFKxyqzEMSesvEQD8gXc51szJc8HlMGM/D1o4YvkPvVWkG+vjrP
RkY8A+sIZK+4sSIK1qq2krtGm5vVbRXuRzx5Ttsaor+Z8Ro9fvX3e/0oBCKA
ty6/r1TIhs9SS4+N4kkT/zdV3PjHW76yzhDdTLLfOXVFXiCzf1d5jmHGXC8C
c0vKBwSdNUY/+hzslG3jaEJj37vh6mpMaXnoaMZ6PWCvE7YjVzaEc1eoS8H9
7wilaKGk2PiludAJLulPvZvle3c11yKopHzjXeeU9F3r3JggfPhc//wQDcEu
ACxgMTbxWRTvt9XmSOIMz8wiCw6kXjPoAeF9A3mOSpDTOlLzg4mOq4Ul0lJ9
6JhspT7a0WI5VHlyoMtlJJoT30ylQk8/nGk8HlTUQ39enYBJyflwuedClQSd
AyZ26w27p+J+DGuDomtVsSyTz1oyCi3lQaJWERf0BtYxxpwKc6rTJAMgPYS7
wLELMQcWhSY7umiWUQRTYqpNMbgr5rNYqSYmn+0ww6XfgYnKMLW0HJ/xn3fx
ctjQnGZa97FzFbPo+1dMnLeopxArS24sRWUsPsSCf1R/EGXfnOm+M6m94CJH
+nnZZ3yL3wmq95r8+f5B6aUWPQV3bZ20qVMdBQiNppKmXQY5tWVZE0psWtAC
bJAztxNEI3Ctj3Q9Loo7Rp8jUDaDHdYQEC0Pob6/ywEWLs2K7wTBBP60BaOQ
pwK7lQPlFnywHKk+OE2YHk9CadlxaIBDxEzxQVfIcvf3ieU5A7JGK0vR81SM
gb7hgbZ+Gkd6LAsLGQGXNqr5CsagPsC7fFSpofJ/YSKUHq9EMGU/8zYSnxLS
+T7sKNGTuTfe4UWXcwXS4QdjDeomuKNf4QFYvBtQJY8OmeohnqjZbBUNTbCv
Yxd6zcEfKdxN/m+1BLUoEkA6x5eaGbFwOvoTRJbFK7S/l7M4fc/QTew4VenL
QAhvArpkS4tmHlP/FITZrvHlAo1lW5Rl3d7f2Usm27nK1hldpSppbhZcuk7W
jbB90wayF0dZBttGsb2H0HqVYbbV3nUV8cQN8IFVUyqC+S4U5f9FysNAJHRM
TypBl43DS49XVkGvRt2wOlFl6OvTNN6JpIBdfG/2PM+XjuMutaqRtzPH/UWt
E11ZcoGqxhBvHExqKxFkMVukPsM/Na37ax9eGHRuhpCoQrLvYb2st3bXfcWN
aWCx06ALqKyFbnixJLtriI+y21zavJSoGHfshZJDK91Fl3nd6pPFq1ckYmy8
cIruTiJTG7n6ZyTKZXlOYQKmGWS8/ZLvhsg1MUId8iSU3k2AneXiSXTiOocp
wMtA0HrGdfQqhS+n5BQyspm5UmkGe8BqtkvTfTCM9Dh7QjmwhTHbqsu0ymKd
5tJ8oEgy4tNTO25ZjmcPpuleVQOZqFDNVBpMatqAs20tzsOal3cp7EnIj2Eh
TG2Y8Mc7nau/EzblRUWTT5ulDI9I2TLKBguPpNVscEiY3b704/JEDstOgtM6
y+jjx1ZmuCCIr8AUj0hdH72Qnd+b7KhL9P2CqWrV0XPJ0xOXnnoqiQ32fgfJ
cPRPHIn9OyUFV8AhGf4Um+DAL5DnaL6d+rJ6tiHkNW0UUWOIOIufvmEMRezY
gaBEJHADFD/ofKcb4Kmp5RtmwNG/UqWmLh3BI1c3Zg/vTlcDbvZ8K69dtA1f
9yZSV+xvaNOebA2Eg8Q6hfK2DPYReh0uWnRxSwkGGgNKBWtegWX3DsQM2jai
8RthLq6+THDifuCw5JvUuM7iwCweRX9mYa/6bsX5HRGuZm1JeDY1STFKgTkR
yd2K8CDXsNaGwIJs5lcKswdv9CvfZfnM9oZOr/cHBguYRlrVFx66jrISR92j
j9X6OO0uq8XLY2qhqgrooo05x+jPQi77tEa9RNMJKEs+K3kUFcpdPvFKAKBr
3KHMD7NfehalrlsO6V2GD7XdZtVJnWViD64GIfpGJGt9JBEUEenfJAq792v6
F1lcj2ExvCBfYrhyeXg24S3Vpgq9B7eGzJ5v1p8yk9P1BFJujuueCrUp4mzm
jqikPf/TxlsOYKNXdqEWeToP3dJw4PF9hn5HN+W+dM2/MyXk4x7WRUxTfDm/
eMFUSER7W3U89LRq5pa+am4+MhZOeGZcMo08Y9mcW+nXiiBzXFTn4xYA7Rzq
MBUhBJlPKSF7xLRPEoShDjeGEFxP+iRFTo4rtb6/Jof7b/tLpY5hpiflg6B+
RqFD9hmrLMgBEYPgTNV4uiLRt6N4FspaqvTuZyKGifLqhaZP4FPIVyJ007E+
UzCVksFauWZb2yQ56hXem78ni3F6rWcjIIMMDYe9kymoNxP947bCilNaY9Wv
d3BCu7HSdq3hA9Fkk9mwVQEdpw2D9EtwR4tpslPDQvFuf3KAYvb17kERZ1mZ
PznVCigzx3XrJHbdoChtBMeoVxqoAUD3a5i/jQzqQF0q7fQk1/zR6FsNIuuA
ZIj38qygWScyhbQDdodLW+AUN2GVZbtxIZJ4vb9HBWrSQYwbFBqtySL3/PXl
4crG1/upt4k4jF4Z6TuCDCcqQatdbc2sy7n021S3fiMqCIebXFckH46Ocbab
UUIeIfDjMuiIQJkiQnyVa5jn7hlO6KB9noNxoQWuEn6994ZyGkd7g3fSYyp7
TjxfT281BYwtFgEsvjxCv90Jo0Xpjdp/d7d0eKbTN8AapA2nXpWihXkD2D4S
yceHW69YRLwqpRxtDff4l1SRvmSxCMahR8i94WnYwkHCJWgMneGCuf/nXmue
6nSqtCS43uzPV+z2O5g8S/L8ECvYnm7F8GwIYPENQL8hTiSusP/VwlEdM4IE
hJHDfTP0HAsRKnlsDSNb8PeKxIqLYsF1hFXrvSFm4knjBUt8NovKDIA8vyyp
b1r+j3mS/TJn7ZCm7zZM7zYBY0iCxl2/yNRluUn5nu3UzgN/T+pyPpuGl5yh
uOgrdTV/STh5PkuzbgQkjPPe3NtSbhHBNu+sDvo7JKnWu1oQl4xYqRW0MPzv
ZZwfWr0aL4InvvIL+LczTkbI8nQt5qyjyV8DNbiK0mYwYKlqVvUzoOkkRc4z
zLR3Ieqyfx25HXtHDupXlzn1OKbZkVfasnDcDImbnSfYWi8TdbxP09HVolTI
J/cWrtXCHWrIxqn+bfrQG0qn2BebwZJ3SksckACNYJSbe7usE4kg+kGPpZdX
QR39XhJkLIvu5gcmKXEH4xEgyiZqGrFf+waShKYjnxZM8Xo3WGEzazDDMsQi
4moYDpnAQ5+PBHUA+6cuQKoL8+CI/QZW1B3mXpspXH6JQAlPLznegwMak8T7
sIa/bf2TNbr6UAM8ao9cI6EmeDdEsXRp5SkO5zuQp55jxqv9ml1xbQtZ5OYJ
sK5OVsfN5VLtm6N4LaaZq8Jo4Vs/bOs+juqvJnPnNoy24sXQNCfFdYvTerWh
Ldrruftk4kCiamTdcsFu4bFqYe2lfIVhrG2qrvBYCBr9X01BB4Lhqi7Mowgf
AAeqG3a3k7CIwiX+wJNO4/RkKELMdPNM9JIjZAKLkRTuq52r95si9m7d/EXX
OcGUJcmTHmzM0qlUb5nIEwbi6+khBehJldgJ8s974Vcpul8lPj4ZbsMWD9UT
QJyJ/aDxJyu4aa+ZNwz7E8yCdBV9NCNsreOd8PYYME47EW3hNlZS+Er2CtLi
0rRHmXpjxncgI/EqDUUon3WTila1j0GI0upN8a2wx+4i1TTK/06voObGM8ac
mhEoGn7DOD/nCyYKRWg6+PmVjq0IeRQVERbYegSivTo5jlK9mKI8NYgaxyAK
BYfsTazuyOYdWzhJVik3oZgOhHlbFhGSr2gPi351vjL5s9pn1T9bbAgrJA4x
Uj2RhTvWqLgLX4ndDn8URHt691fV1gBB+ppSqojThtrsQ38y0njj57e5zi9R
XtTpN8r3mfyOvdoUzVoMWTc3VozuLqgh+6HYam5Zptg2/RWLB/i73U7UV2iC
/wlEmI7x9+DHDFO4A2SsHt840Sn0f1BeE50ySiV3WtLG7A59OY8PkB7EiuKF
C85fZakQAFmmYERg9jW1tHi86saRXw6XmIbmDNOEWrmdpel/4vzYqlxjpFbO
3xbNkFS/Qwl7qCWoTkLAH0MtPrGEnlNkJhHeQGZqmuv2KQOVR8cQhGFlNx2L
Fk99q3S6lWWH09+YPr7bzJoi+yfM8fWXOqz/ZU70wxc/BT44bP4myIQrpnVT
4JBV2enacWMtOBx5R5PiV5DW4tbe4JbEFyAyEB9I9SEoVdDFVvaUyHHcd3s6
sV+NrseNQ39ZiGKWEFML5Wqh6NLZI+2is3DI1XJeylI5u9PFskdJCM+OXvqX
qXPAW9cEwNvllKbKIjg9NpPjwRAiq3+qWbz2Jba4Wtm7rg1lyAPJIpgTFR+m
SNqi+5leujo2kdYdILWLjNa2OHUbpVrxsrHm+/pEGbtCt1+jpwCtc3hZWJFu
XRMLY0u/ky1770D1p2NJ2jpLQ/xTkz9zbMtlUkAtn/K4v3pQnsAYal3ZcWht
bzP8tnCtka2TFtKM97Mf2vvO+UYk6u71/U3wjU9RV/4d97pyEiopvLdyiobk
fbvu90tY7xGnITZ+PRhD5InbUDiVhHwCmzDS9S2HzAPg0doC7+wREGnLBvkp
5unrPeOq7TDcNGKNULSk8hdVcNsxgkQBG67IGvX+SopyxtwgwYD7rqb4iK/C
Ur0Ta8I9xRwgNiG2fjk2BFNCuga9whyQp2z9C5APV23jRZVSsbcQkIft/rSV
cwVrFuFvJNLyBDK9h3za1avDc6HhgtLJGKN7VB0RSoB2Cz1KeVFf9AbARyUc
1hf21pvYuV+wTxSMFF6smJ1GHl4aT6XMuGj1OoV8GQWypVcfDGa9NnxTzpNg
fPnBAHeYKUi6aMXQ5wKQ22mfrBumipjvWceDVxwdMNJPjZ0uCooPV2KDktzi
UuZivdEvhBdqIxGQ0Q/8yyyr1vImZUnNl822Knk9XYJ55h6x0Piu3k2/XX9A
d6jIpB2H+5tehvcsaLoWForK+H2zGR7Dpv1wqwY3bhNjO+ZB78aHJCDjwZcY
7A4BcoExsKAfr9QlIroxjRQ9D5u/qP8Qf1pHxFH2OmYvaHTbqM9eXCPjea0S
qQyO7nBW3lC8YCISTlpXC72E1dMZEnyOZvcVc/Ld7KVK/bGHEEUpEbDvMcoU
VQCNunErVjAjz8b1suBhNi0aZz7QMq8lgK3TMfiRTt0Lql6Ka091QQ3bjeS5
Iv3fa+5YUUDgSSwg9vXQCD89ZH6rDjGRngBqUftxw6jwP2VH4NIPynCNPGZi
38O3cJJBMRB4+2Bcqj02+jR3kaRKTVJWTNZ/iyxUT+KW5tQBmb9kp63i2Adb
9Z1CaYEID2fQPAy6kbe4QXy0EwLpz/ZLLK6ZxO4iA/P6yWiLeee6fI6RQd15
V/0zFTwLdbKcN64Tck+sGrmElhJ6lUvWzPytoiWsLmXznIjIKwSDSyo8EfJ7
F9AOPgsuwoPfsWeTiRbuOHspIh8bZC6e8Zb6yOM0WW8L02Revuek9KNKuHYU
0vWbw6/yDuSRz4ilUEtGCxlmCdwUEZs+AvczqIYGn8S0BBj2uWCAn3BVaoNC
5bzqbmEl6VUTaWHGq25hT4TNBvodBvTUwUIQSzcSzdTtPAxNyXvHmozWSr8U
G8qvUqDWVoSEIkqxtC8SjX4odhQ58T75tsxPXCvT8yPLJYO88hOtX0dtfygb
teWpK9HTwyYEEEyTaV7JS3uuUNzRlH+vNtvWXfixalnelZQ6R0eVLMd6ImRu
f5Cv8M2yhl5o1FnZw343qYkBWMoUj/enOGxkuxtAfZ192mSQIa121St4LF7q
PpBa+ud2N99e5RO81yuL4jYagD1lnmzX50HobFkODFm9pnKj4bV+vmgedQ6N
9s7VLthGtyK40xcawUpCmSm+T4sI3MzGBOoX3rD+AzYcS0sF/q6Qq6AssJGR
LxgFPrHPUNI+R09chl9i31t1J3ZIbpnLM82yxdMrZJa0JpDr6+UWqwbodjen
fzKWdrZ1pjDzfPiTNMYdxGncBe0jRYth/5RrlbhK7ohEFfZRWE2rW5CkZYNE
w6VbLRAtILXDfBEmmtt1hOxc/7lWlF8sqgqumnqic2QLCfXGoKrm4V6Nyl4r
sXcrNPNau8RjK+69OTEfasRubQqFzv1mXpeV0nwiutqAFkdAhaHPy1da3Y+z
VoU8B4Dr0uCW5YCptvYjLxQPyJ/aTBt6qLLCN8lPPFNHW3Npe5H6kFqpEsHB
nGDnGi3Vu5m3jJUi+KMcs5UIoEmbuNrlR/EMPBs4LKfD5N9ei7vrivyNL6Vs
zq3UbdjsbQ+P5N2jp530vNcld7I8oM9gejGx2oduw12Cqe2OGKUaIUTWv2pD
8k28+qo222kt95WTmc8hER0zIdCF8iGGEuY9mSihRB3RoJhMhI6kbWGKEjF0
LFdxqk/fxLxd6DVnqX34Y3PwMERvTqOHObQW+4hMubr2Rp9iKBBsHjVcwPag
8GW6SRdf46VjcmvmxYUOfDQydLOjapV+3XRi+6S2QWnMxF1tn+OZuE+2vvRy
8500if/xna65+0sChGFXX0tNIRr9z9AQkHwrG02nK7UT++qtcTvE/WfYPcE5
12+BfLXwJ6QBHq1rlFYiy3iQtLuJHaevUiRgVPyFYOT5hMnXaEg9MzFGLSuR
Am3unON8TePwiI6Pvg7dDokFxARzEjsD0cAIPlS0DqHqTzA7K0ou9i79Saq9
EOrpVTRt0Q4iDH0ztoFqMCKnVmazhb+NncaK9UYsHmz7+8OM38BGA76GflLf
dhH3thwGx6LiQ3FersLkJ+aWR5s1N2e8L6G5dBoMzSMRmF1Qwitu1pe4TdHz
cO2VXpDC9fx0Hi9KjJL27GTh7AAoiRulQ158QzEiZLnd5DmuCMHQxaLGdyGV
+h6CXRoRQh6fsU1PQCFUVlrO+ybyoQWjatmV0As6v7SdCbvoeet6slms3cWp
VblYOpJc94PQjsJf/TniycjzucVl+KFbQ96a9Q/lrVwcovQqxvTfjkYL6ZHO
f7N3kzBPnVDciS7U+RrbW+Q/sA5BGBvYJdTFHBrBizbWnJkyS244k4mKhxD9
EQmzgL7Bs1LKm/LJOLWTnSiAscpnnjFYWnmBWCekN+xQlXIAkzc5H8U/8X7u
g4tX0MK2DwBtnNLngPiAUzf789BuacKscYVI392uPgOnJvtkcfB8x3ciruuZ
u8Hnarbp1Gd1LoImfvwbhfrz7B8Pe8DohZxq9LYgcMoHJ9up5LevAnGEb5ZM
j+xUxzmyiqzsZyG8uwvhnKbq9tt04pvxQ7TG1JM5RdPrYj09M0YsOEyj+XqA
RXdVXa76S0FFzMBPty46rYzeie9bDV3tEgFTbwaBkr2vQzxib+vBkv/OF/xO
9Nurnl7BbZ122OmFNhr0gm+0cBIKLo91+tfolsAiwGaCtHuaR8xsvT6Kc1Ix
t/eVw8RASf7g2FTvqFUS4ufu+ih1bSiK/zaHcu4nvNRwaYupALNmPrXoBUeY
e58KgKY1FUBsU9bXUj6VvPjuuWTNzJIGhIP67dklEJ8DkN5S7c/tvq/tIuK+
KcXOWfSxguG4tlMzrrjuDgP3e0Oz2g27KfaVKszzc7J/P6U9XrcGC7IsSl7T
1RohCdoF27e1cPxqAA5Sez7YLGpZdVnp/CdrgM2vhtIc3n9RQOQFNfpLddZH
1SCyzBbP9nm5KnRsE3kghLH/8EhooTp9IQgKvXw3JJk7L2dURMv7yF/1ulSN
cDSBrZacDlcDGsWzblUqzzg4PBVz9TAm9JybRTlbVT4i02hPlWshPt8uRiy8
DNz/1eBmf3AtWzxTgMBijAXKxGwMpyyuJSTzCZ3I+T+dQ++D4ZzCufWHS65j
A/tV6kCxS8sIFGOfnv9WGYaPaTZutN/nJmg/MAdrbqfuEmi/DS8rMZDhITZ7
gBnVZYs7YNbAyuVekVBSMJvfvORzmo7gfCys6XsD4yNVLFEzqqfdZcYD3o8T
VRy19YH8/DPrRUC+VaHPs2BEgkOhsndBJGlw8QIEQbskigOdzzUOgyBmtjYf
LE2nJUM0JLnlIT3mGhu7K97kjdoTWZyVC3XvYrdvm9JmCW3Mypg3sGKgGs3r
bcPqgD0r+MUtOhWVQ04xbvAijbqBktu5eV00bOCLrLC8K1sTUP1FGzfZh+Hb
QXc4KvxPPa7FowQ9HDLEaskEigqNwM6z6qpUEUfeyzuAp1kT6QRV/gVoKI+W
66Vus8UulgbJlPlHflZHWvWWX0Wkpn5f2CVcR6yWVMQkAanmtJ8TRRfqL9UP
K74achCwghK8KE+Xvwl+VcWlKVQxD01czMZ2/YQ6kJLP7NJE/Tera0I82C9b
P+oJpUB4cRP0t2fEHS61vz0W3Fx6GCTvoJt2IEeBJ9iCChZFAPlAw9ejQorh
gidY/hLzG8PhzrD9PlBs4pXqLfC0xaQWw8YYIshev32zePuqSb26vVYKR6ae
e8n2Nw6sBidDXxR8/r23uVorJ7tLrtM7Vcc91BQMO4SUiUafhYG47frLchZ2
OT3Aj4qnLd6nMwrVRNpsid8iFOVEb/5lnnGTXm4FNoFqVCk5bqMHzuwIbG7I
Sk/ah23JJusy9IyOU6da51x9aNNRO8PQ6HTC2Fjihq6r5cJTr789XJkpAbpe
4y+xeKh/ZgdPg3O+ravqoNwOkFaoqfCHEA6L13frIQ8Z6uCPpKAn403pvRgc
6HqXZ9xJN0TaZ6CYypI+CpkarY5lgT52Tmcvyc0DGsePiUmFc5S0lhAVMg+E
+bj9XX/5Ad7rrkwYsItIAtbFCKO8m9kUtXqbd4B4whOYbE6Td0cQ0X4irprB
bQ5iBGA7FEdz9+hWTxV6LkK7xlePD6zw+9RjBQ60dYMpWydh+XxXXtVw1YFd
U4e+/+R1+IB2EscsKzwDWLLFO0g7FDt4Bci/Lyjs+8ex4VkFVZRZ8S7TLzJ8
7Qd0htBklEPI4uPnNv6VtS+gBwGKy4h/7zR1tT5XMoio6K/NvipS26hgSdW8
hPJ2lD4romVEq0f01Zzqx6YX41FHTjRFWHLsY9UpTSM9bopWW/r+tA4iXAo+
pksNoXRKjgVDB6EZvRT5wlTLLlkO9P8Yq2guflJxoqpGhbHDFlNX0sxQ3GgP
WExdaRXuC+3VdY30egXWmCksv7AGmUMwm6tYCBJOAdjXzE508DqlYbRe15yR
Tx9hSwryW044ihKp8w7Cs38ZJ9JhDDyobQ68+19Q7PcYa5uymSUIb8IvibbL
OpaM+2glvHtnE+K/W1qDTeT6RRmpGiKX+aOWwrAWP+3J9XiD9+CFZ/CiY30R
DjrVoOBbzPGQsEnHMCrx9HOYg49VRN0y5zkCg2jxth79FByQROen/Lqn0znd
cof/+Yz4RSr3CmuK0nF/8SpVm/iXTJRJWZcxLPEsCpWIbYg087GI1PsSBBtf
jCNOFhGAYy62bZEXAqzrEWppxCPfNXU+MgiNRW20zKHaQ+w1aYbXDZn9pG5V
qrXidRiyDLTYBrFmRxtoThiUiihnCUxSfmidMdBIPl3LjaUqCB81xYpS98Ps
h+/ui5I8t4UQ+tGJJYpU5T+VvzZybYnmCVN5z5z77nRz8actjW/x/pMXFXcX
pfY9oMw4Qou+IqLjqgaH0iZuAX5yEIVL4GoHyEQvdb2kIAGaigVVYXIl3spc
S0tQWfZNgegPeBZw6V7Sj2DYCh6XgEdmO523yTJOlRTn2mjbJHKNHr3TPpV1
mvUj5id86J+AssxWICaIlkfBEHegMXo4dFjxmRqq4HGQ3WsXeejUWcXgy1yt
u1038llWwfY1MtFLiLIkotkUiv/LoOxhShsieDB2q1ca5PfqQOF+k+TMgNdW
SD+9xQCpRTlLgp0To9YfniVkt6fgPU/V6vpB/Xcm+TIdSoVp9TVt2HiGOjkq
Op+pqoNVq3r+S0yukMf1ZdV8fm/F1BQM16Mv+t+lNMcCuaRutyXQCQxVo0rE
1d+P14l6jHgeFGFybOYbsZH0tYN5yjn60Ws9A4TDNGbC6jQUFcSYPwSJAuS1
V7C4/Vqn7Jo0ohu83LRDdr/Of9+sreya5G/qfvo0K+RrIQiEZmNmV/fndvKr
6p0zvnE4R3osq2u7jTd/kRjk2kVmxRRFJUgRPvMwxvWHNzJUgwO5cR8einnA
r860wYmFtCGApG6FWjz+pxzXKJMrVCzRizBSpjpTAoiVX8yyqaB3ZVElDaki
0y/t9ro+GkeelpDIcikR6c6dEiFFIJeIVxBZddR9qpucjSEgSaD13yrYz5yN
ZaSL30FLZmx/M90wEx/ekRGNu6hKH4Nm06a5DE/ylYpB0BsKifFb0Ft9xUf6
WXoVdbJ1gaAafIyizYSH3HlR+MRka1YoqywM6r/o1oPLkYL9mCYIoXD5uWuf
DzVp6Toc/E5Ay+80v7I59wWECwgr699az6UmQdiYAzgFIq4p+/UjvT1Jv609
O+hSjOKO5ixyTWKr/NEq4eWFtDyB9baeqqZzlz1ZfDzSQYhtre699P172XfB
H5C8k8JioaO5kpmwm5LakUL5OY9SHrgDtif8iI9f0zwuEneTBZ5e38HRwm1m
B0mppLvmxdcPCpNPCGCqSCKv7X4+LdbyxfThskWtER2GB5YwJ5uzLUtBg2qP
B2+7YUGczAsToNs11jpNXry+7/qVx51Ab9fNyjcOBTh/rPc+I32bHFgov952
JWuYHP7beBU8Jw4Q6TVCTIQqS+y35kRA23poZwzDj0K41bQyXZNPgspTZvMM
LI4OEWzcSPYBQBkBouXqhUeA+nRzpRCa6Os6oGxMENFExYyov211NAAwgWri
MNDbZrC7CAY5YkVnhHXziKZZkuAV+bqfSNFg0ZNRZ07rdxMWat/CT6nTRnLh
RA54KAPGG4T67Cdn6yW0q1/kvVp48QBK4Av5hW1hckNueMazGD/o/XnMpL0O
bdCCVAwwnJn1y3eg3+JOlb7y0B+lS6EfPHxol1nwvHpGku3eN+z3CetwUAyG
Oj/pffkrDhh5P8u8YsK7SvLKj47+DJCEaEqsB1JN7Zw8gSplKhV6jHA50MdW
74qSfzmunm5KagO2HPtg69l8RWvm7iULUg61mP+CZe9BUSJ0mnlfAsN078EJ
wx4WrFGGAHjG/zRZDDH5w3LWYP97jvcpk6uhVtAM7o3WD0dzJez8Wnt1mwyT
XvG4TnMSnDCYTAHeV8z/aU8TsS8bim1ouqSMmwlRMiJgs0Qc9p5CR+0wzlko
T5XK3TbyB7pi37C/xpq6FjWkk4lUd37ickKuiNORjfx/rVGTwtLRwLgWEwk7
YWFSSGtUdOetWBoLAqNukhjKrirlomT5ZCmLZzNfa9N9LRUh+1wA4T6XFopV
+JUOzlyZ644ao9+/Bg7TeEkFgUqD/teNyR/lneL6g6/owAyTwpcZn/A+aT9X
er9HnTUw2FfSxRNtes3RK3dKJmibn3SRWnbVufDp2T98G6bYpDPc1buDWFPc
RTDcuV0mWz+GCiIC6qdTczurmQbVRfukQ0k/SL3CdtlUx7K9i/wdrhfl0HU+
w0eYAAj/W9eR+PGHvQjMeAUlV7k8o2xXLbJsJPOwbzLic8heiZ5y44ymXWIC
+pX2KGdJJkHE4HOJblFoBhXxYB0ZeT7KEsx1TyULBQgfR9Y1Kpej5D9P1+4d
LAfShkPlnSWKssdYFrPXv00yhQa6oErauBVpCQLTwog+KLWuC6FEb9ixTcas
PAZSjZhYE2yvc9TB98Cifco5N+8UbmxzZHs0QY9XXz+5xYEH7iSZGHxgq5OP
17KBuG8q55zT7JOCU3G4r5TopvUl1rNoHLeBp1oG7rr1eXq0saqytOusnAG2
HWk6ii+/QWmAUrcGNjEK8sqNj9n9utz1F815Reg0Z0Oe2dh8CwzgnDzRtkgR
hNoBAMqEbZDk6x5jzyaLDbTJ6U8eqle/JOwdVm2y4XvO5le3SegKdrvFiaZ8
gK8lSuTfk9sBxiX9Ai886tOXjpyWRxMYVM2vdUuy25H9fy8JAgSyNQBzHXCB
nRsugFCqWpTUSMgJYWqii8YagjT+9QLvEns1lwfM2axBxYqrYyzZVzNf3ifr
Yl7lx2aAxJYFOeBM4Ri4B8yMKYd9qIw/ExkTTJ/97kspgmpS2lBVZXRqLPgd
r142a5EXdNnY6aTlQyHXA6AT8tBcTpIeru9r4XgupHEDHQP1SRVrcC0P8L/J
gsEfFVRY3uNA7ps+/od6xW6I8XFjEcTewOGCJSoNfLsNIH5quAnjSxGE+dxu
HMhxQ4VQC5W1up9vCH+xxPtuiBCfXoZjjJVhMX+csdTz4qXGdiHhr2ZFXVJy
NW4AiioT/RQaeEmrkTY0d8dlJkl5/M/ibFSOkA+4uW+ThsL6kRKfaTV98Ehy
tD/puls2wKalBaUmipCLLvis5/xd5PL5O7XJO9fUkqrRvvH5fifVkaGnoYzr
OGKF4/rsCKQRNviecDyn/n5CFehT5IQdPUMz4Uzbg8nUbaGA6+gPZjr/Ztj5
dCnJxL9aBM7SCP3CTNgYazaV4OY6cAMdZqFVJX6mXuvMUQqLQQq+bWXNkHNh
5mHcG+uDmIPJNRr3dvXQ2EPV/onNHyi6eg4jB3Y/H2uLQ/VOIKyDIxxGZczt
oAY6hUu2u9CaS11B7az6g4vJSPqB9x/QrAUB6D5bEIx7UqpkA5tEotNi9x1H
v9pbQhHF9GH8lCdf1gJxCL9JIW0d92ms/nsMWxqwTiEVGGX38QMbB2HzsFuA
kdwLKtc3WQ26n1LPsm4NRmqTU5b5rvVGKFAzy4mvqN0cys5IJu9I+YcnBFly
Tcj1qNvfOCbNw+zJayCWcDA4QxJWcJsVzCauTN5i4rsay+T7nw7unveqdKim
d7PCRCl8FptydR2EN0xMD/3ApMJYupUdbOhDb2rYVLBVeaAU7JrewY2tgDqh
oZ4Ao7nlodXUTP9Tn24qiHhXQ+yxLIyjAafai4GDfw0MRlRdE7ay8tYaS3hR
TfHhXDDqgGCIdIel827f+UixwWktgD1GkhPb5XfcF2Gs5cQ/+AqE+m9NIYIh
2jN2YM0jGaIaiAKSMqDSJaAlXK8PutLEiQCLBurfqe6b1d4xzrmrs0/qOy9X
OS7lAnsPYCngtd4XVfj9GxyG2VwNU8WlqUEsM7PYJO+n8ycPED9Yl/y+SPk7
av5c/6rcsDN3k51iwKWxp6RYZLwkB2YVEF4QbtMeEq+0x6WS2Y3htJoNJKUQ
v/kcPo4Fec4TxCE8LP9L6+txUetCWr4bj+sJGjjYIGi2jvclslYTrkQs4lRz
EbEAOqR3ltjKEG3kLwtQJ67a3t8T7XuUxkwWBTPrUtQJpC4xwBMyPVCNV2yF
X0U/Kyazwn7hVq0KSdJo32yD/fYv4TJTyNEKRlEle/XeoqDNfrktK8aJy+N9
sUKrtJtHz0k9rSv8Zs9GfsWzM6YMbKljnkAeKbM0uhhEmvAi31emt1KMg4Uh
huPi97Dp1WHJKzrSfOSkenFScgGmnTH1p+mELlsypaXhsz/o77fn0akSZY6P
PksYtKIGWU6LbMzGVZWqIPCQqqdvJT4wAZ4trVhTO+mcE4sW4Jy4u95h5xtF
cACX8sP7ti4czLalLryZwiAJ+ydx4X9WoDhSY6bpdmpQiVIPL4BLYx1vIXpI
hi1ahJHY3X36G8mEeBHrs/okF8Y4V/+HxRVN9MJKENH1vkIm/NArYp+gJ2Rs
FwjP76mwQ7peNeo6HbS99HkAFLInqhG7k9FhNsWKNEL46C+PxBebgsFBE9nd
zi/2QDOifg3eO5VpVU5OtCt4KUXrONLO+OEUgL1jGbse+4cvCgnEO2MjwKZl
nbyMspAsID4jIi3+GYSYo7EBBQ4QI+X9MMWvMY1AskxeBnAalgp6otTtyjel
YM15zUfL5CmD5+8tr9dQOLWtbnyWMr8GxVBR9qxSsEIlnT8pmPguLvjFp8AO
4PsPC1TOaBVwuUwyMcHDmRrCKPdnStLsmwDG2mJ6dAynwGcTECq75/iEjcRb
qZNE8pZP149JBVRPAP5Mf7SxX3tLgCAASoM70shB9eKd8AYJAyLTjz4SQR3F
J3qHV49bAq6+ZWjz7ExmArplmRGZBNEfACCUAfLdiAYilSiEpGSoQxYTu1y+
s86qg7vhJYGhxzceJPp98o3dhz46XAUdUqwTR2dM4SELSIHpzYGhLwQFIn8x
p1JoNwkS+lb18QjA1LLdXjEKzq/fuDzhyn0xYkZvNb2dP9pb9n28pJs0R1Cb
TZeImfRjP0tCvH2wcBArCr4ZldXqd0TvtAh6odjvtQseg9ph6j9sqwY09plf
lp6Ifm1pVpjdUOjmW6DKNCKaV9Hdm6fDnwyXIJBplykm7E+ESfBlG2Gp1EsJ
Z0wS2LnQxQuidRpvqtFqnGD+/u9uug8IykJPfz7Y93AqHuomcT0DzdW8l74V
iXDFhbywOnBqrE+nvYuHnIMhMKgY/aSM0j6FPubV9zWPJEM3BDg2NEsIPibf
M+yKDJ2eAjcGAZbhaCndbAtk/SVowYEbL838DjwCKIO66e9poGRlsU8Rz1bX
5DueG9C8DV3lyZ+dAlsQBOhIbR5vIBI1mEsK9aL847WMvemkR0YLxJQkJwNF
8gmwZKELXuNVimUV+t1CRGVG8sar+YpgHsBxfmV836moNKLe0U4lrm0h+VFS
n3aJ31ldJfyPuk8zXubjt8UE9QT39+eWeaclzOjog9EHgUqrdIRv4sU5+7h+
b173SoNBB+9AI3F/OuRiWLxk5IL4vddGpj9HIY5yZ3QqEXKuTOuRPANOq+DZ
Id0tLxyS6Bjt3vGv8o4n4B8wGuGTW567ZPC391qXubx2JybMOFiVusDkH3OS
UTSsTI8UmNQdHOaCGGl+vP5dKHih+gJY2sGoa2g70mVfgoSW/BQgE6I/8VM0
8FbUHYUYhyvZ1/iMTJiizsaOuxDVU/3I+YBcwSsZWAzLeU9sQXnaGkmCGSJD
rWX4R9GNDA0CfH3cWvLE4ViTi/3ULL+SubhFhvErcSTgeikoFKHIlGWd1DTl
AiOVQaoBov3wb3d+9cgekoFgDrdHQEisXJolCNcRfy7q+xl9Um/MnLWhAilk
BxbEvAXY267RPibZ57av46oL7+RwX5ATh9XNxES1lSepYYGJ4bekq56alqt7
EjFRKnOBCddbXsOsr/o4JBjj+h4VCVxIleyqMzD5UBNZ8jE8KiEuq6XkTrYu
htPP48XSzf7YntU9unljfuKPQdAyhyjCnPN8XPjpulBbs4tLhtl5Ax94IT0b
5QER0iASM34J0By7h+k0VH+5yw31Tc7Y6knovSdwveUfihcI4/UDE6+jPk+9
zaOktiPLDSIOu3QXFsITNV0ESeIJt9cvdPeOPFDwx5HyxAO2ycgFa+R7lwTG
89nscgvs5e94aa7pPG3UoxnxyHA3073KDuY2orUdLamhq0p2SY2DkS5iFC63
z5TRqkffJgeUnHVknpnTH9cJvXbXUPFWm8Ei6tj4nBo2vtddAqgklrCewJfv
dDqyBdl9Ueha7Ickff5ie2q61M6vD+3KiUhCoOPmW3n0Kg/zhCw3jykRZ+cU
RBvCMjaaiw9tBlWJJj93P4HZs0SiWQBUMRU8jSQvzDmtVLeXap+8mMkesF+s
HY41HEvLuOBY+T1mkygBKMY2PH4WFsaQYOATEuk2hiwf/0uyj2k3OywVNz90
HkANiH2NvbiQ5tOHOIN05jcVoT8fXmM2Az3ggxevZo79jppg8z9nCBZfwEt1
OxnLQLG0f2z3TY5uPWaEoz7szpfrqug0DqOysC1zw+kBtcPajKnFG4e/2+2T
0p6GJppEaR5Jr9U2lhDOc44saBCUEiDT2DED0vK40/i7w9wJjzbQnzIJR7QB
J+n+e2QQ1ZtWksq7BmFTl28cGuKBLIRK6offEMQWFDbvzSIPoUC3nETNEBSb
Sa0LEbEQ3K0ghQQANvlM/TXzZbCADABu2zv9ZpML6YTT7/NJgiUbRSKW/SKO
6PPAl8dgMyyiJaMk/ZAgjMEBTxsYf+uhpLkm8o4kPPZrpFVp7pfnnKV9WXpB
vWltY2EARwhVVcrDQF4/AWcko5ew0edOflxO2cTU2KAnT/oplW6Zu6KTHhKH
Tyf7ZVEC3nFMzuLncJ+T2ofQOuhUnadZR/1RKjX3c2TDdsMBhWd+awSi5i0e
OcQ3iydIJiNUIf6f5KYH/HFIH1WPB2M4BZ9FR3gV8xR36OsVqNof0kDKKy+I
Z4X8r01x4NHcFjyjNyoQ41RMgCZxJiZTOTrZ+VQmeXPyberqgEKmnUD8/BSO
MQD/zGX0j6HdgTsZ6pK+xOA1lSvmjN4VgNW0wYqxmZQEdntWqbRSYoZkF5AH
k+kAkcVGDwynLlPzI7l1gLhA5nnCXb8oLPS9gaOp85rO33qzV+HYquUuby9+
tRkun5wLnt+wgpx4WEMYQaP5yFMtq+a11jOlnDk15EnvuXELMNHYaEQo2IPl
mFo18epBN2DhOh+D8w15chhN1oX+AYMJ3PylmNOxlL3tGYKLF94yjChEbZqO
VB2VHg04Bl03+/i9XcEA5C93gwEe0f2fHKfLKlINRuYreQdKm0DpOmBImD05
FKsalSY3lnbckXCVn1oHugqdzDeg1lEgC1jyiuNZsxx18j9NCBqUWELUUhCV
V7RggcV4103+pJaGZzJUBMh1RuWUvt0k5Xv6k0qWrYfOG5Ue6auATWBM5O8J
QFfC6EdTzAAeC4sSj2ct4Medinbh5RIl5Lg3cqSf8Ak6ACCzaXjDP+YLNdwf
Yx6M62WSz/BXDd8eqRpbO7vfV6BrdLAz7g9c3RTnk6bzu+aafHQVgb2s3s8C
oQfMyqf/zCdd2sFyecQcutHlPRYqPnnb5w372dkb8hCbrUU/ceLS7hMukWXK
kNF1b8r+2R4a4ZiyXPAh7pySZzJtYnqd7ndP8o9va0eVrW3Z7//BH+yp9MQJ
MXabp3B19T4/tiqUv+BzHmBnotzFmSC4REyd9Z6kex+60dfmC3uJXzAv1uOW
nsXzGUlF6updjOEsIsP+jWIq7n0wsQamzH4Ca20F+Ph+nQtT3JCgjW0YD8lk
x0an+V10Bo0C/WwqDPcCUJsZdyMz3xMEGy45gS9WYroCIDwy5EGx3ZnI7eEa
WynmPa8Km11GLDsjDjH16/PV3xuWsVBC+vLfNDkJXRx1wyEbp5uvT8T7cMAQ
g/zNjCibkkUKcpRL+TG/NtvoJLxgwO1D7OtkARvYaK3N5x6jLlfjOlztdAMq
1TO1AGllYszbzWoFxEjpjrCuwrqsdjG6ye4jP6j07VUycKEPV/qoEtkRG5C7
LyU7pLg9qWlmHCqQ2xaRRYaKVBd85+RnqW/fdgwESxq2kTC5tlHR1ZRiqYqp
rqzvW4qHKV5CioG+A3PPAcSvklNFbBa9BdzMUmJbYj79OSo9NeALn+wGiiyG
8jV0neq8orQLUpFAV/Z8tTogsYGWVxS0joN1vRRFOaiIFX7/tRcQTw+gVFKC
b8NulF+rhOqoLXLxiYzEbFIUykkG2zCArE0lezg8PfDLAqWbSv7eMzf6kM+Q
lvEoYHe+t5GMIt7XXJAw52tYSIpnHQ2ebIxRNRRZxbp6xQev1aRgIZ0h/WXN
qT2uSqybEM3stZHRy+NgF5RGleYibObmhSkYZXemTRZXXPZcCYnkzwDmXjdU
KxafSiExwN1dxGM8Aucuqg1muoaDzmpL2FSdM5X/kKXnD+PbhFnoz9WDR8fX
4cDd6VOjo2KXjrpWSc31SGpq2YsdF5KSzS4sxbqPaJcEkGQxwyv6rMtHERaG
dXFmbtx8QTuh/HeuhtR7ZpQKaNUgPyI3cvIcb2ajaObD/KemfbPTNrRBV2Hm
lMy2vjzwiS94DQ+w7r6C5iG2W5Hjn/viggH7TbpYUexXVeZgdYSyzaoHa1xM
PdtCYHgNc2JBl8yxRcJzDbN2kdNoRHM2qpDBr/zSDuQ2XFqOjA2Uul9OvfF7
kCl2tZEYgLfhfuX6WVvO+3kbbovNFzO9y2Hwzzrego682Ro+HKLJjunhwp92
Cb//i+4c9KeREP3TY2ituosvmTwCk0FZ2/xKCJqjNrnc9ZTzflLahmDDCmSJ
OrvFPYUuUTrNdoMmbL7mV16uEApGixIkqpfrciUvXwm3ufKnsp4cS3zQpfKj
7wNlzt+xJVleJMaA7JSfeFqSxPND/04Knq5LrH8gE68Qv/dFa8bykg2KIuVx
rQNwntw8H7GgLL6DSGIaONq0TYcWcR/hYgPEkKoWuT44kZu9qJmN4j/vMbXv
YXFoHZmrfuukyodFU1xoF8inaCxC1WgRAqBXpGVhr4iQJU9nLMKFwptCy4cx
sU1HHru83x+ps34hz9HQbrJgK2zLOk6mPZYvjoqvK7knrP+3WhNDPDV5KMy3
88BQVDS631H1V2nTcXHZWFueWW01ptaUxLvS23nZ2KvFl6fOeWR7hpdpfWEB
TFK07JSh9v+PPKT1ybUrL/VtyoKyJjLhpxsTxWCStq97PMAZFF9XT7AXzhVe
uHtaMRcigHb5izJ7hX1hNb5IN9Pw0bWrXPMi7zUecWBeeAx0mp6eHKifNt1h
xxoEzvS/r6AwX65rnXFx7LqZ1Kt0+f2OLWvvhnA04gB/HidLu3tBvMpi6463
t/53Nl53Qio09jYvaQQBH+DEjEfPDd4lYocWRuqjWSLCK8sWu0zdlO7bYrnj
3dnln4qWzRD7bPwuXfvRUTx35OMuQ+71no7hmIwPn8Oljt+RAcDc8O+ePiiZ
ieriymNGGlAt5pEDI74RFHlAM6BFgW/1HKEcfK4MML/7lGJx44TlNuLzzlwZ
WhOJ6DN5smEfE5n6aIDtmPtVT+CWLKtuHY9yUI+b6Iq9c5LjsHWJ5y2JUryu
TOo4uzAUKHRzoV8xqZEzuHi8KU5HRnb6GC3N1/OB3sdoQ/ZUH8wvdW8UfO4v
vaVVNJ3GFuKC4ztXlu/vRVWo/wqVEkl5d/NwgJoxHtvDekuyz9h0qer6ZVKJ
mspq4FXbF+lb8X17rWmXeEubWWOAHiSz677a0FSwNq74aCPj6PXAzwvnQoc1
fh3WuvfAKNI8ubWbK1V0oS3KNLClQT8hxQ59LHrcg4w79QpBgcLPiI7KOFi1
XYvFVegR7uJtqRelIsD4TQqBSzKcfREggO1K0TyjNpCjHcllyh5RoTdyWb+x
LUBc9C2T7fiCRZ6eGm9JoDIlEuZ88F4Yqi1/zIg1ulq4wIRP+AYVAJCJm9wm
7Ldh6pggRS0zLa4f6bN2dWFcjj31C94c5tmGcTX5Gqmr8OEUN3A3PZCNTyoj
8iUfZN8BSJU7pcar11TjU9yMu6EB8vaeEngwcamGbtDFysqsXLxFHXeIs1iU
AuaILUjZEaV6CNnQoEShyM4Odwkf1BsvV1hMW0Utq0jClfRWaVGKITJ0RvZ6
YNr7/1LR2yFj/X2K5CXT5K28d3GPBZjuAQDeV4n9/ZRogR6fcmAFzVrEJ2/0
eHu94wG2DHUAsZIZvG2nn6ZZ4wMM5DmOzlufiWuhgO5mfjMFr+fFnY0FX6K0
gPhRcU48tPk8m2E+ds6Ikoo0Ir015CzWQxzFtujPubjP6H+nLMHn0YKIE/9d
Fzf1HtJ7A6WnjeG72DIWZ4VWYLtWCVyrrCdGCq9EwACH0Iwv2qL8Cvhkd9z9
Lp/pvWroQAwAPDYwZ4LRNAwbsdt6gMQeMleCfaLFrBfiGnrWSyfvz8n1A93O
lIkC9aCZoLOWvEcH1akQojmmh8FF+xc/ukTs+t5XyoR/OrR8ClBVEWYeTtD8
exYwaN7/RDWIoZczcGQWMLkoGUXmCyUvS3kWFgDraBrcFdthx9gBNLhaR4kw
eMaT7m41vzDwjYU0DUgtYo65BklQAn23gqMopjrBdClG0Pc3+1zN9KSBYC/q
UE/34YyohouBP+7Z9/xRWDRZB0uLXmuU96LKsRXUIX0nFU9AxvW/rJ6oX47E
TBxmaOX81q5gEMoHOJiSdHEdY60DZpK6WcH6TGAOGo6DpBnZTj30BxB9gNOC
a5HyMUqfBxJH+VZ3uwGS5hFFqNytG5CbH/619LKeD07EhnW4/wjMOXVzbxta
0XE62xId0krKsKBQyWPkUhLkyqipKi5sjlfvTn45yszIPus8sk1by26gn0e4
2GnlJKlREKPqa/mZi8BxcAR/sxGC/hyypE+l40zVGjCaOiEV+xOH9O8i7pLf
z6bP6xH1NSB4tGNz+LbXDTtbPVF4J1hi0n564WtKM7ZHvK53Y9fPzhlxsCSn
Th+St0PIcefk8V89sLreer8UZfhkhA/AA+L/fZzsgGSrx5iVD3byz5yKjU85
apJg7w/gcBVikwf7CIjXzMDJ8Q0QMmswva3BeCvJtE5MOcckG0paQ3H00Jo6
NpFVVU8oGXdCy32ogYxfKogGjUbNbhoPW/pxHJN72x9kdhIPUsfsItP/K6lb
HMwZmxXU1Dq7bgdgrx/q77STL/tHcHU8QyKpg83aO4WCgS6viyyEUVzXiRzY
A+r+rTITL9D35aVItdvuXDvhcwjOmliBtm3+Ivv1qWbCgqWqPI93o02MgyxG
9zAfHjZV+PXeKRwJorkNRK9XwLf67iU52/EuyY6N11oQTTmy2ET1uXaP7Vci
w8Y+t+wpir6C9tNs+rc6Rvsiw4tp28n78OHEPrifZFOeCncf3KmQLwDpSP2K
i1S38JQAeWfttiMUVBht/dJ0Ye/f3uVvTUwhxaf+4PaRnkALHz92IaFcexun
sU8fTNqtz1yz5ReAhcYM6gWbb1fj1S3LgAgyu8mSjx5HBqBWhHB5WfIAlaxx
mmRIyRiJK3G1UcmpCQwFUgM5H+HERJLIORDKk3yAYTZ5sS1eaWlJRU8nBhGv
IPco/BPkSGbQn9hzOFFLAPWpBPCxpGgvKjD/BTdg8laJRSJ6xbbG27CPvK2X
hU41xlrM/pDcY2wOx6U8fUpCVj1GHj2RUIJTJGjzI7Chwf/Y4FhW6Ri6WAD4
hhxiwE0TzZ6HuH90p9B9B59RJkkhfz/Riicv/YdhEqQIF/Qql/ecp8eY89Vb
S1wz7lnnh2SwHFxgUsAq5AyQ0EBb3/HkMDNZEnP9bSQRcgxt02yDGeZdIFgV
sQpboe0oOgycSKwu43oM32CPB/G48MMrvcMizAdkoYUeZd+VaObJd5mp5+F5
53E+D43frZwS6aUKf+usthrQFtVnn3yynfMjA3VVi86vgrZJjSSel7VORj0K
Ea7P98C9uBUpN5fp520062QLeC/5/ElaCIutBmM5vB+mWxp8zdc6/cr8l1uS
ctn5aCP++waNaSAqdTwVNKbPhLGxIcDYhZ6lHJ3hR7UvRGFXaHFIdKq/kKjX
j+0OoVVUeQnATIBaCfrhc0lMCi2ow2QCGttqFkTV114/H3OhtnKgOIcTIMb/
Ky7UHq6Wx9Zj2hZ/GOcln/3VMV3ke9K/+FLeR20DYXAZdMOkER/ItJC1bFLd
LXth2g6fXR5imEYtxrFBr1SXK8TSy4WfaWrTiQUZQmKzJgWnYzNOSS21pl/6
smODy/29XQx4Tbu3c91YkXR45+3H6GgH9bm/r74S+6CCKqhJhYQqYvMB+C4w
4F5m+1kQa9NLnVTxjRZStHLwuBHBMjCUS5V6G1mmTKgfT3kO+8xXZgBWQ51l
3gALSPR9IhEcdaS9/ImEEUVmy7a6z5XAXjfJEbj5jm9Kxuv1AYHTAO01pwGj
k4Y+e2gzANJlZR8dt+qR5lMMlXl67U3jc5dc+Bm5W1YplpbSSLcO7sqyQc4L
1gohy6kocAXulrxudJAjZgPVnyazYUS4/bUfoL7426Pxds0pYxI/vjT+fWYX
wPlCi4/KqacyH+32uSBTDSoVmkSeMhdAecYbPH5yxJgcENuqWrxeYEi48QLw
6npxwBno2hbDXhQD/9d0fksmZMvcdzJVHOStbxM7yGIkxxh65lCymd4KuSDY
0J1r+e8UOwh+/dWU0J84tsX5jf+hl/wDtE/CWxOzkSeAI4QI+kPvzBO9agm1
uRLeAUzb6flWfctwETJSZnN7UvARW/l5gDhJJxRutRJKWM0Ff9oltSNyMR96
YHc7pi7rBD/wQuH5oxa3f1RuknmbjoXTQh3JNArkEKWBSfaF616sybStpFNy
4kr9xnZXHAhASbtRF+MrvkGzwUsYZMcYwNIZQRpBb+vPR/ePTejnOFIW0zE9
BH4rgGNYE+o4iJ5JpR7bPnP9140n4mBIQYwxdA8u/J/rHq51iiI8TizvhwXR
xlybo3G0gTJg9iDAc0Q/jb4BblIvxsWc9mLm0r5Ad/rs2BUZri0ccLyXdq2I
Kqg0HbV3XPcSK/Lx8KXeDmGl7UZAWiZ8ljOoHD6ZF4gL6wwrRWlxjrZigEy+
iDLeQFsQbvGrFGF3lMzwY0YmlhMVR12enC8nmceJu8RXGtxrAIqsNLTspT2c
h7J0AVppcuF891u5DMwhsIuhadOZF3NDPioD7lRqZMAKNqnL6SV6RVxAv59W
Hnv/HJofRkQRNZvkjtBYjGDQInY5TiiPQ2ZYNjiFoMJ3k5Cqv0DZyT7HPbE/
AIgvRBYn/R7UKB0dz0T4Zs/Ek4xIrrW+bktONfggDLlzuY+6t7aeJMCmKNMf
zPssgQ/MXPSpD3Wfv7Psr7IpH/+b69nXuCBxwzbiagKfzQ8vH03C33ZBthcE
qLNKw8b38QcacevhfPf1KjLZe5o2kfRiPakymiiV+TQHcOuaN3svK/n503SS
pvV7e/LeJniRCQrku0F/oMCIb8e7USQKQfMk9leDQYhxAlE1U+/soAr63MEE
lmoF1178LvBpO9asVA2b0b1/Phr9Sx1Ow2b+1JorBapZC3Evtb/uqtvwd/tU
wKot0dlpEVea8dv9KO62KIbO3x3QafoE8Ty9EseiKYa2tIKfzazMnJ7qSNtD
hQAjJQl7px9CUOSSNHwJT0yLfzLoKf0Ons3PoOleiE9Zur61kOCKF7+eAmBQ
JG2uC8YYvvi8ZHMMXZFMkNNaD1CrUIT+qLAX0MHi4uRrmQlQhfQmG9lQHafx
ZGAr0ofM9KLHUXVrO/PhHXps7ZOruZvG46P7wbUIZriuIbMqSRzOREtMsZz2
zq0/ZHluuvJOBJGZXwfh3u7jZoHc6U3A+Xc2if9bV3JLKyd5VnQXJ7NFEtCR
ZPpBTkB1+SkGghaW2JMV1IXi0XfJOhYl2YUj+GAKpxe99Lyc/4hWlusVBNsR
FfI7yDU9TyePmCpmE7i1CvoAANj+HsPG835wtYxEENAyjmZ4FU3NrzzntAXq
oJ/fP01qlVUj+s3zPd1NMTqc5GuEi6MOw+2eh+jo/yF49mYSHMygXruKrOW1
UBIrraXZEa8mCfUa3PGkmucyergM+BDXfnld/Sp+O1f0QGNUItMEP8AM89pB
D0i5x1Y7GEII1hEeDKBBhe9E0FyeWRpLj19Pgc4AkV9DdFVw3pqeNraXon8y
UwsTXgI2+uMHPdGYxSzszSXbQRzJZ4qehluDY2uRvFaWGhS9u8O3G4Nbt+3a
4gZuOXpPK5wpjFj0OK7CJQLECo2jE66X43iC2P+N+xai8wiv73k5TQLZXU3y
+BwnTp2ElSZVaZjy3pPxU0M5Znu2qzzkSAJMe8dhB+s6ErgnKfoWTPBxWr1t
ofmq1yHJxzY0/Pasb8bz8YXt8PFfNYSbyotPDAP6FynDFgEMY8unO7V8B7RT
kVoPrDKXDpgoE39sCBIBodZjZw6Trf2wE8jXf3nOkqN9noq1vsAe9lcQWl2X
AmRnQV0BXrcqAyuh8RUq7HH1YChUVzgsKUx+gm2fPa6+4BjmdojhY7xjp4/X
oDSaF4XfkpQ9S2F5oS8JQUDIdaZcq7f9uJbiLUd/XH+b4TsJ4lYq4GxuiScf
3c/PY3UsILXV3HkvCdmm5wsKXQ5vQw9jAqasB8kEWEIIr2qEozv/CGDnHCEI
+4wAAjIxErRha/g+K56nQy0DNciV7tmN0A8dQA6Avsui/l5jBg/CZsdtBjkS
CvLcGG5dkCnuwbiT+oCljeryUoJVgSzV9a1m1KYr1GPkO4bBcJlsjvSjwZV+
gCeo77uIgJ5+rY7CXriTmLENUr12Hu9pfZUjr7LezmnvxgVrgnmeFJtVffhN
beRqs2W2UOc/92m58e0kJQm43qWX/iOw1hWoz+vtxKIyFGwNZo4nnN3hg/AU
nPCrvv/BRcbiIWaUHyqv75mwExGA6R/ckKhz5PUKarBb38G4kPfJlHA0ku8K
teWcO57xeFbxyJX13swTyRkkaUPz+IhUDCzfcs9bJogLue2rcyGXjhGJKo7o
bOphOfQSFKcQsn4x0KKXlfPNdRO4phCpZF3GV8+4j/U7vueHTwJgk2MdaV70
600Gp1KLm54Ak5H4ovyyy4VkrPAAVxap0Djkv1HIveWl6ZxtIY21TNOJLibj
hG4lTx22GJKWxUIGrT5lj+TerMSCNf4z+Le6tMQzO5PHrjxVqtGoLj3wj5gT
Y0HGxIUAoE0Q0kIvpzFBhr7JEJjODlY5LN9NAEjOEERrZogQAitSxe2QXvUK
jSdMZXV2M4myWy3O5uArsMWTu8TS29RrZfebwmMQ74jLu6WxZRuLuqIZcp3D
0obmYFSTEP8ciFn8Eh/NrAZKNy3pb2L0vk/fKvjq8GGFb6L+G+jKFKhiZsYn
6jOCWisrkttj42JRqV+em2QEEup+e7srq7pKomqcHrMJzZnIBGJXbpYsg69X
fBkQVRlm1YI8QvDuU2+KhqxhS7CQXWSw7WhEGQbqZWjmiJ8c2oMmieZKkwqi
9cu1f5MvIMcdN73ziKaOygYi/FaeHJ+P8cg3JL4t9qqs2aDu7e1gAmwcrYyB
82yayBDLd6r8iNWQwXyIZLlqVlHjl5fvoJT0mHvWFOZ0dO3KM0qIKcm5rJfp
meux7TZpeyrf5D3Vy4EXH9J6e+lUlJuVZ5owDgDb9/nvLsdQVtoPylunYbrx
dHdhAhXmDIa2W1Vmapj1b7R2+iTD9NmCsZH3hsudq1dDQ2vyRUpE53/byucx
Ox5D9xG8ex3XcxwxPAgZrKwJhMap5+r2R/jEqZq5iyekG13dVTWrrZcrfrbV
bvnkPs5kuMBYj1c9TWjPbDu6vIiTXsQSGXCP0FL7iXRn3hlVUv7jaff1gCBD
7MMCwwY7II2+gN7sZHbafaFl61u+zBgcTN9hQkxKdE47VkLY4nQgzbKb1lk0
EpGh/f2eKGFRXkmG1WnjTk3Pl1Rp28TDRRqfPDGUYW0Dlaqw58nPKzmvbyLh
hUhtuILEDwNTtA1J/4KH9mafOiedDlSvZb4Ib16lyRzUAbwlTBBkoRcwhoh1
hYjj2ujp8TIkH+7NzdsCZeDtqmYZFaPkbhxh2mydS9e/gfGRyADNjdXb9yms
WL70grKLn8FHF9O4a4O9bovEyyVKFjAt183tWAUr2fxPBbnc6nuitOobJ1FB
udjKup1dNCQ6x8PlC/rCv+4dY7KzbXvChb+xObcLkoMRKBHs4t72OUuuB7Z4
PS71YD1jncmWO+S/SDn8v3/sm4nGMx2ZdvyF7I46gEl2wcCEXs7XVKDqDxXd
7m+pvA4gyGY8zhaPHXNrYZgIJzLXwhM8UpKxskWoNTJHe36+51n8AJ5Fuelh
7UYHhZfdrMs1S5/yRVy+0vc4w1y6z8NYCnMsKPpt4JZYdeGU/eJ6I+gUVx+6
8fAEIGqRxq+8C/TKoSblNJJDHMi+6vZWzM3hV+gyLAVkKj6QtccMvNFfWadf
btG3m40UtEHUti2M8UqgBRoJMgSQQLT//j+QE2KrDVsUeUv2phkcOkFrUuz7
ItP/nN0HNTghM/vL26b1c/WXpbEf+zG2/vQDpL7UaFhWQQ920ofSmiZuSorC
PdRgGBT0hxptWMfgd3CAs2v/lOwLl0ysjrSxQNrnHir5QzAeZhoTDT88bJ+y
faU1C2ZZOY/yAf/o29zvJ3wvt+mV/U+xWb7um/79ozQuHTyRp1ZdSRe0PKQu
YNAZzvu1hny0AEMjdr5TLkiXJtwW0H7h6vZYo+uplwCugm71jfTfYwuH+LSC
7at62Lyw3NdobUZljYLVdbE7VRBZs+8TsnHt0hkuzNgqt67DgSFZ+IRxJCEp
2SPdQa7IWauuiQNxQpZuwMNz/c214MPcPcHT5mT0u9AL0H4pAl6w9+elfnif
J+iAL2cSKeoXAuMMsqQmkUsKqSPLcZ02ixgfB7C+k+XrQt4Nif1bgv1EddDa
9HV1GImCcTkynWjjOQyVqdupuDTmL4fbmcGyGbm2AKmddUqaYK4WaatDI3mI
Plzmf/mOPV/omibDb4DK/RHFhhvzpolJJKX7wJc57wY2EntgtShrEIAfmZ2R
hGqoyvg//CHlo3FO5e7RWu32qmsVH9Kk/FiHAdqR6dCIBthjISHsmA3p1CmK
RjT27CpwOHIbQfDGwzTQZaldxAl6Nq6ID5uTiNf6R5mcJy2zAzz9+gDzXOf4
vAYqP/VKvdLT46syMLhUspCyKI1doNHCWerWypF9s6v/JVUHODGB85YR3WTj
HZ/KWO+C+mHR8EVy+kiy3SVahPlfn6seNrnNBDL0KY74OY2jgWURb+badiqI
uE8r/TKbF36hWd2YKjihpDszpalLplIjYqC/kj0OPQDO8YmCx3TgS23XSWRp
xaybrMMz2aYyR4dAwKtfJuA7OZpzd/ufkXdPSPsB9gf2Xm3HL3TQapTSx8Z3
HDroP10lU99trR6K/MdzKDxA2wRCAvrwo1I83y8NLVXSRGNjygyLwoHQDwnu
Gju7+YuW9eYgCH+HiXV3s7s72D0estttKNewFEarzXYy8Vzs4QvFsBrs/84G
7PLSUPGir5TzItikdNeDSTIjuXpHNX2v8pvFFMWGmScT59jvEMnX/ANm67zA
2Dwcz0VcihtI2aeJf+Ln4kZ2REnjrwtSYlgMC0xnpdIc6RW/uqE412SdpFeq
DUoQrRaPqjRa6UKR60qzwpZuO9X397W5Y1lRthAkc8o3ymQTjhfPsa/Pqsjo
JizqyM9NhMSkYPKWoNtDI3+/285Fy8PCL+mT//2I6Y3SYFtawRf1ZkhE99Im
KyZjh1/qpS4v06NxCl17cVFALFIMImRWJO7eG4H7fKhH/Cgn/vISwEgP4/1q
WzcMnXLndyWprLIvzwSS60f7RMn7Gx8+uJi7QEGiOAX5FPHhbchZJBZcktM5
ngCmdJlnkN9PT6jzYG+98CYUeLyVtbcTBVAsNv4yia39vHV9k2N9w2V9TyHg
JA7jQFDCgeSX9r7kpoyV2H8AlhIwra0A1vax6d8Rl7VkxH3tGlXTlD4DZWoR
EkWv+b8dhlVTS874CxYtX5ND9EcY0pZ4+GFldBRiGLxKWvvCMCDJizknJ169
NL6oI4ryhoE43BGS8XqtNGlV0XAIbqJ0OIDyf6aT0a8ptRO4rsMNvr8Ce0K4
wO0pM+RvZVY99twClcS8P1dUz/sU14178MEOIbpDVh9pZ2QaLQdpvlgWcqn4
wkvQyjTOH16HJWvS4DEQquOpOenM0F5woY8PLCw682IV82TNI6C0TYckZKsS
KaMXrbMXzgcWiidk7tvcWyMzMBtItmB8C/3+M2kUX/FKbT2UbAgMXQRugKRS
aie3UewoUO79UZtpV2CtQEjuuby9eLPRJnPsG5wnuKfYlUrTb8hpsFHNYTGm
488L8UWbRg8izjoFqoaQLc6rooYUi3rTy9wr7eNZKATsmbuGL2Vt2S4rtAzm
kuASLVPY3YqX9HzgFfp/nsXOAKLZlDnFwd36Fgc9QMCnXqHyxjt5KJzD4dU2
yVNnzaAIZslVoBqGflN+Pn+O1ACzHdZOF5fySSjA/PcA96gA2woEwmJ3lOwn
o2EuqOgDyJcZdHNO95X0EMhZVYwqR2yfpc6JE+9NlqthjMS7EYm+XyKk3cZi
A/yDUUyfMej5a4qUJ8Hw9ZgmAFjEPPxYbYTbyII5521Rd4/pbD83IBaq4oWD
jeldVW/R2u95doWpQA1OI0RXM8mDF24nylWHMm6qqsd6y2GBVijKlMdz45Ft
gwHG45UJtttE5yKRF16yHRi4qmjD2+he1WA3V1YM96IMYvYf8UVILDC2ZrV9
rb3ihgv84C5Zd0CmuKUG8w8sTYtrUwul59xzd7q1aGwSSnp39CM4iWwwN2/L
IkEKfD1zzX0SroDhpuVHf6YYvVTY8E52wDz24TKKpL/YC+MHE+v1J2DmBipF
yPmCJW1QYuqC37SJRuJFgxaB1CfvnEyn5eal/4/FpZhT3KczADhCTcVPSJAV
roE4pQhUs8Chu8QWTp4UTxZcxFmkOjCb8hDcfbxMfWL1+joEtWnWH6ywnaK/
R/V/jZyVv5Y5XPE3KxphOK4NSUZ2KSJqFrI+zLTml0hVcDhjdP9YM6UFDMEa
EOFyMtMVPdJbX0xj3DAaei6jG2/CSe2Qx4REcJqdp7Nz3KRFKgWLxm8DvXXG
G2ufv9YdvxA4mfRFRJjQ/r0NyeRnl8AiS2K6ScV1lkAmcepLact8RGXV3vDc
C4xWnVbfBns7fQSng137RC86ZXVOtne442iHsbRdupUmG+nbYzdjFpD0DxXm
nX6Jn0tCp/QySxh3BQ2bpCjQvize5NjF4xhpwHkdWx0dbulKrivdFo6nszi9
OKmKqPue1P4bE7RzRfdcgNOAItoPP3vGMlZ+4Zn07lYta/X+8+xim9iKXVu+
mCm9/qemmmACs4M8HMTDaBeDN/Lg+cpSL/4EtI6jwp+PybvRPbwvwdBqTVlE
fU9UzqbE+iZFsSwYtWN9ma7gm+vsPZ1L2QTIsd62sgMW+ha8r4Rrp8HMF1Fr
4Hj6BXxbf28xoFzABdZlXNU3ZCvVEi1zK1MSYcgLYG9zD+s+Km8h7mympysy
Q3JrKFpXw+id05oGH+uehNSUAaWLMqn7SZEh/48jNkp2xRrIPMB8/FQT9Qtk
tEUV3ekLAxuLqhETtvgVCL78YruxiTXDHI1kxpqjptXFAv/2k4rpJaZgADzr
k/dItbVcbO+myM8Z21vmS9whzC/A+rCRFlQKHB87EeMNLx5Kcq1I6WEr5A2u
GLLn91TZaB6iLzvzA+Y6Si0BV6yK6EW24No+FFoLvryQ0b8b9c2HFZCCRELr
0BYvSe2UYvoMQEvQYsP3dV4GIn5K+GhAFhIUipr9zwBmajs5DMCazkH/pVlP
48YwiSnDqIZYOfniqP7Cw+XcG0S7OJaRaEmXjEjBgRZXl7MemrmuV6BpNYo3
NKd4DtYWH/mFabldameMMK1ZHUQZ+VcMoHpLZqhTNXz6DZ8n2wMaDw4bV7A5
vSJ3FI70py4usxqXGVy4TLIqtFDD0xgR6W1jf6YueIIVZRPayZjgx0QDBBMr
g+HpM2+aurjBRKW2O65fiDiC9FTImfgWKdiOIapXGoyCQxan41Fp+MKw6fya
nxiMUlIrJpv/3VZ8BJPczdRXhXwrTVI+J7DExnSoHfcKwlUYRsP9HvbhebGj
gNFfJ8hXqlw9CyCsvMXVGpwUR6bDVjTDbx+yu3mOLUy1wFXCgY5Y0ZdWQewO
x84ryfrsyUI/OqUW2ZvpAQICgzToaXQXMJUXI4ZRpssz4Jb+EyFE4cAbb4/M
Z5PK8qbuCOfjlowe1+WfdiFehbNajjudqltB8H77P+6w2H/LTajbNhcDm5Zi
fiG8QYtdG4MAH5TD546JSw8b8w4FquGxDmI2SCChsjALTe7u1VwK8S/iuAVW
WbZkdhQ/Ytqd5LPbmnXRWODXesLLPkp1w3wrj4dl65gMogkGt+5TY2O/DXDG
4WBIoQ6EA9lnhDXz2K1X/okiGtwNhpFKz/lc9cOxaXXalxJCokdk+9Uyf3fK
GBonGrKok/JtH2sqyyq/KQZsYYN2HAwZN4EIFoj7CJQ3l/DKbm90ev6julU3
JLFhk+6mVvITJrrRKNoumoctU+/qlFk6gipg/ndkHwVdpP0EbXq6L2NNC2WF
mtJuYDIvSl08/iwemYZ/p1AAC6Yztd/uh+WwyluXBg3BWvYRrFsR2OcOHPcL
QGlAaRWbLLWj9fbD1SxXYm71T8SpJimhupj8mfnsOiz3KaJ7pQMtSoZG2oo7
5hIuDojP8PuN6egrqcWiBIKXzMgJdBaZinSVAVnfauSRM52gU5bTWpa861wd
HglT3g1TLdNYS4ELhouqAmF3ZUmOgljqW72vahocqpw6jefoBvkYEZdKtMhB
h8SxeUMCTD/mD1TPA09IbmCG4rjoP7T4ZAEiMED+MBqlotX0QSEK7knwHbZO
dE0Qom/XXKXoRuS0QyejvB4Eq3LyKNG7n4mcwIJsro9vOAEYGHrLJYdoq36p
IL2GQzCasKWTqJut9Mh7H7DZ1Q4tdyjmYyZ4gW5LogGAkFbW6oiQD+dida+R
Pu6H9fCxY86+RZcc2J/whuzrY+oNRyZczajDJ1pQVt71tw2IGWL0A1jMxe2A
i1iR6Qz9teSocUDoTfCC/xDpfmR70bYMJv6s0ivARM3GLWQTSo1bEbPdQGSp
UwA7UN19TwRAw3U+FKSwXFJ0SiOyHhCsfAAAxq6ruGb9Wm6YbashVgIIsIGi
BWrfNDe0KglFZA+JI5q/kpD451jR6bAwyYS57Y7vhK8qfRwJrSKM66HTdLb+
2UDKixJw+1+5uFZQ2E2JuhVaRPbHd+Preifh/yfA94ggR0atwTfVuUYSFCn0
g7v8O1hRj27Q7mLI2wf5qNbgW38+0DMovEuN6k3Q+5/3SUIxAFIKddobv4wC
lY+Prqx6zTopMuRLvCEiKRTUWf2fQ3N0S490jfvr8rhK0ZaD9feE/+a5+bUw
87a/qTZI9tCokjFV90Zn3KdqgJGpeRrm3GviOoy3hkzgNBdJQTgRwrv0VQHf
0xRi+6Nu2GdBgPPSqhVxWMWcsu8KSp1qFUnc1Je8rCQA8e1SPluwOCQtmU9g
gIz8L9V+9ts/z3/XEiT04gH8Dv4MywQwfgNluZVA1+Rjev3b9vH1A0LatYQp
UTCeCpeHnFHm5rKVCIILjuyhRsAVPV7j7SOen3lj5b3IknnC5egZaqadp75z
6dkvDnbqfOFPCvnrhpMMsnMjoz3MgODxDfWA0cqfJ5nJuibVikeo9QSQHhBQ
zZeh11Ic920iHBrDP5wYBaTP63KF/b6F9qips8Le+Hc0W0b8mRYEoaZqTeZ7
4poC/M9XjeM7vUVUmisEJyjSrdVEBJEUjM12aygG1IDarZS41901dkg//RV4
R6U3f0UcSpayn4/WlJcWQ43NBpJGrMU+lHTm1hLXPtvyeKbSsgcEVop7PJIT
yHRXhQoA1VQxFsbVne0kzEIZnzhAOcFISt7mPb792lZ9W/4MMaX/RFmD/smR
feGgU2q99QRUtBrvn9C9kHejRklH9QrN6/I2Bxal77cnqHTSWZALiJkkFWPu
bMLsjsou1EwJcq1vuYA3hZtfBTcwQSEDEsfrriH2Wj47Nuok5P9fZ0EokH2S
v977dOFrni2irLuwAcuag2/E5g6HtdK/aVUtk3DO/IbTQsfGhtFk1RvzGP8u
rgJijZYLKTm2nAmM6OVz6+eo4axz/znQFUpZgnRpZiSfytFVmAL3m9P8E6sJ
RTCmjI1FdeCjZMXB+an4WlNeLN0zdN03GBGUoRD3ZRQhF+feNVXrWjA98OxX
jQuSre+/O4iyDsFE694yxffuxAu6nxm/02atEqaYNxkb9qrt7QMnKawDSarU
pmUoGHDc/0ui1LC2O2LAmLLOxsx2p2uagGIvopYlJU/rehZ0usCNElysg6pl
T+1eddJwwnkwwHWFUDOAJrbrZkqkwf14KygMtRFvxv8fOnTtyw024sJ2YVHc
SQOAVChfo6/3C+5czTzMXdhxdQha1HJ/AAU0ieWwkYjFRFC3SLORvePV3yiE
zPb4enYsBdBqtNMx0+te6TgF6Dw5I8AOf8Tq5rKZetSuijD/smasHdDAa2xb
SZ7SD9gfOHYFcD76GhqlXeAv8mhLKjeo7Kc9cojUHHDVRYnNDAB13IY6UuvD
tPvkGr+zUzXvVK1g7aS/Nx8z8D/CMBhCOvH+yMYQbaRHLc4a3WB4lc9YrjbG
ATe1KEJ2iYeAFRGg9rPePhUUAAMycTRWK5dJqBzZ1n9OViQaKbQWNTufd8Dw
67S/AksnSZ1R3CIk6WHdv1t7ugO5fjQEFqadr0u7PBuVNLZ579wOIDgW7T3Y
pI+Cr2HkLg88vPgqtv9ZCn4wMd33Vgat3B/vj+kATYruyfikcb/6I6f7RasP
RVYAFLMB+cpBzImjZsrh1RCH0GGOURRS7vl1dkVLcXImwV5Wwcqepsl0Lhcz
mCit8nELpelvp+FuNzgYGnsDweU8CupnAjtP/O6JhRov7gNyQCN3IUaQGcQ5
PedXMI9dPa1XdZ1Eg9PWK5JVI1X/8h9VFQE3nLb533VvmeO4YRrP+CF15Wil
mlnWGaeOv8XDtqT63/GX21ZGsPwmks198q1VDWMHdRmyOfIZRdP2vlhSf0vf
szeYPVeVZ+qsbG+/BWSLwhVzqRD6zyWaHv6B4/yR//rgi5VZlG2zn/2MpAM8
7qa9RC5CCQKs8e/YF2GsU1zA68M4rr00IhtaL/566q5cdqZk/+XeoJT5Jt1Y
vbwVipZ3wvJb3McTpS3ib+eVcxZ1Ty+MmlseArUVieax8g5qgyywnFs/vKoC
lVQTD3np8fgJdzKWNDSpM0ZouxXqx7sEYlV0RpuKQ6/RMeOTH6Vd0WVJk+OG
2mG/vRmxemD3d7AInYXIhmvNzQ095kYDD2kkMT7Or+UWfig8pHwd/4GreTu6
9HfBDu7bdZGY5OLapFN464C54gjH5uJkJ6r8d/ErXJNBjuhh4GpLCyPXFdW2
jYnORxNxFSJtTxIFo/M9dRk49mcb+GeTk7mD78f0gY7KO+KNBhTrPJOBiRbO
edmL0gfPG7RvI6umk3/IYsKOfTxo2kaPb7EPwBgNHV/Tx1hl3PEHpw0r3tmk
+hZvBwmkaUM+OES34DbY6pu5JU77f/bwErBlfnmH6uCUNaogfHVfm5Ya4xwC
2wOlnKsEBCznMEH5LNQ2YWoarJ9dpLCoKgM+jFj7+PXsOYYajNEHt9Kj4xb9
NvD3tLr4+Fd6CYmJ95vPwDvz6m7WF52IQ3A1fvjbSedDlAU1W/yMyu00kSUh
+0iRKxXZYsNpRCe5ZG3GDSz6bjD7Gfc750lLLi2Qyjk4sUYf+yRbieakcTh7
Lo4jVClHVfwU9nDqBCbVirSKrj49MOx0rvieDsFkV42Sy8vJ10RzfSr3dstO
gHr6LvPooHQNbpCS1UpZ+l667D45ouQ8fSyY4clEk84eXllQEwdmZCcoaZXn
9r8qWsNn7el5+JAkUj4ODi6sTFcJ3G9ZZ1y4jmZs9H+uZgg9aNNQkUm/wQWF
S8aSTTPqWVWWFQiUwCjnKV9+63L8QHr1kSZjD3zLSXEraqI8Xq8xbDe6Y3ZD
jnqKfIW8vOHVU5GTjYgcTLIMVwSey4x0/2XHVdhLxCWsQplZlCozz693lZPV
FnyRJUms1+aGpmWL/0/8rTIvXsMDuctSPJpNXV4yz4XYb1j6lw6O+E9Dts/H
or9AErxbLREiWaNvl/bBjKR81Nw/jm+x8uTwHi/MsvvYHFQYDYW13Y/Hq+EK
OxCBTYGab25ubX50P9b2Pqw5T5tOM6CsZlSLbuF7oYRntFQbSG9BPypcCC/S
AMNpxnZznqdOdfv9ki2HGRAJgQ7D3laLqT+UNgBnvHW6VWds3dU+eyv3mT+P
8KnNKkLYdhimpzI+YJ4FEEHaQP5sUhfbXNbJvEIM3g4DcxTgrk5ghQ/DKeFQ
xZ+cJxWxhW/YuKBkoZRURQz1TbsCOffHwXj9DIVPGTnpxPg/+A6cATooXLTn
PdSUWzmJSoaq9fRj6yNu8Pla2HmmBJdGlktVjV3Od4M8p5iEjY9/pbb6pkZr
BbqJL+3Q2kaDjKGrLyy+GOPOswjnCqecneZFm0Gj3DYLREBckmQieQOXUAbd
QDK/4PiG6YmZN58ZlCwe03zsA3PJDH7kjtbr21j0SEhqHIzt2VB9UTKr0kng
SjaurKi5HDrPqa0KrzORjfGXjuzkqQcSHMgVOHcTf6KlqB6ettvTMOg7wXZA
mbuPR/rpaCUEe/hWY2pk5OuASd5/WKSik3urqixXyJX1E9OJH5b7zEgov4Qf
Y9W6Nr0FQ2ejKYO22/v6EJaD4WSgMliAwmlK5sW/gdlZ8CgrY6OtbTj4fC0r
OtH7z/r7TzBALrazn3WTXEpqByzgzDzmYiDVN2s0SVZ7RAkZdSdzJabVx80z
KexDaO84DjRXV8uywFQ64K3XcdSMqtcITRbzkvuf3zNQ6rtEZdi3mZ91SbXe
6rDLzogay41WNw9r0+lwtBC/0hZNzyRdwLtSIoE5L4dVfYirCCTtBdUAmdNR
JTu2YxBCrxY/BimhQicXxpP5vIBLni2oZz571K9gPd7JY8awcAaltDtP77Bk
ZBAxc9dJK36GnZeE2gLnJRMrJVfj2CvBza8PN7FAfiexGEd6Ux71zFn52T54
pqy5SQCETmg+vE0WQLOQxyysCnzMfiJAdrj1oyfob9a4R+ShRraAfxboXRIC
q33jhJj9CknKSug0sAEQhBdlI2bz8fTrHIuIwrSVph7Pv139Wl/Hhu770q48
IxGqFaQBnOLjJKhnCHquzdp2fNBpqLfniqJN7Xq9/LzH958Msi/6SNbyIsTS
KEQq9kbaV6XUOImx48vrjQmVVzw2fy+quaO3bu6SRG+db02Ea+ikxhjX/029
Y7/B3X8lcnkn+wte5pNTC+oZvjlcyKvuR0HTeb7haqvd7HAgAmopKT9Blaz+
whBU8vBw+GH6xi5xXlK7SBf3DSmevZkCTJ3T/UZGMR14GvXXcf92yacJTgeV
qWkwsiOcihG+hH90wy9uvVrEPA0jiigONzopkCSSKvjfFmRYCER1mpQG24Ei
L+AJnRa02g7uE5XAw8duo7a/tZvItOIfw1yxSuYOpLGd9OWz8zvHnlWQMLre
e+2iFcOUVeOe17TaOFqQB5DX2pO3qBZASVEvNHh8S1HEhgjB5w/YEWbaY7xt
QdCN9hXPBnJriGsp8aZpS26oxO3+E7holHS6kqUPcwgiqQZCmK0qO2lev3ns
L/Ak7XC2PQ+TXDL0zsexaEoaLYx4O3Hqdpdt0anEENfmeFYgf4YVC1dHVCuH
kTX/G95Jis0ukoO79ECuaKL5JV384mId7W6Tcuh+3K79ZwowG0TRV76+tL9h
D9IbMlZNuEdcFwjakDnzBvBTGyTSpgCSM7VCtYaUWUDQOfs+Wy91FzvgFkST
9akKN3+p+NWjQDhP0ySroClu/DacbkZMsRtO59CHNB3K1NbkeWcDUh4NgOYk
JPjJC+s0t+w7gbAQqRA0wGQvcOU4o1pdGZXb++k9QIG3eHSJ4gIsuFp2bdO3
1/ALdxOdQq58YOMPeUpFhrSTjOc8h3DsiKaQOvm5o7B30xnAMD5GSjiNN5kF
3uR6F8SVGXG7cnTER9JocqIzqbOdCytziIgdGdWNzmqOBapRdUzBUjElitPq
HTXJs11l5QoJO1BA/tqBFB/ECJB1XF1CfdSLcI5X1012XBvqQPsVnZ2GJeDp
pgjnu5sIrFK8VkAGaNahlCZA2sqNCn3FXhFfvqkFn7Mi1HfOTZBKWw3++HUe
vUNKgMb9/Zt/hUrqJcvWjJnf612v92XtGp5AtFnyryF74bAkY2Nc1RukBxdy
+x6fRDqlPimIin3+9br28ppcVulQuDoJul5f89VnDwAr3pMbY2eNSylPixsk
2socETBMwgKPRrBCpX0bRfyjY0/H0jpEFheIZFhZk/V+8A1flkaqFyvbwtWd
5cfuIRR6nmUvrjl39d6B9kbDlrO7UXeqFE6S+oMvx070+CYMcdz6n/qE+nI8
j+3qD0TvBGUNsLN6uGJTxjB/omeuX1iJFV+fbVZlTMBT2eN64es616l9uMMC
Z4TDgwbtgsHNLy6oDX+Fbl88DsFv0BHODs3l4zYQlw4uB1/uRURTys3ONTob
qdgktgaE/v7+w1IIqj1Ei2sYrv6FK9/oyaM1Rr3CHnoORraNgOQ7J0y2M/z1
mXIfCosimk7KMym2AQ792+ho1X7GNuxlUvBGFjVizr7JR4vhZvy83NNvHfR3
m3rq1EAp3cBsBVDC3fRZf8/nnO3CwUFw/56vbpWWy5HbJA+AB68Ky5T7Ugjw
3etwc4d6vL1u8vAeZjCn9m3wvSYUXD3jDGG1yU2FOjncgfS8+gLoKqP83TIG
U2b/8Gh6SL/oR+z3ji9XXIGXtNP3M9C8MgJwSlItPLC5H9I7Gqu4LTAnF0EC
azv54uTZIW0orIQ7JCTQujOt6DLas6DTuQ/2vIAYp7v0yYfLRnxPAfqFYek0
kv2gcJ4m5p+8zirLJdm14ZRNFU/4WEKz/SaEKP7IL4GBH5+fw0RuPo4hXzBH
Mx/rnd1AKC5lTUch0Uk9vtoI100XFZmapuTS1nMuP+UiKEuBlVJhnA0c4795
RjLTCZBFByhlKC5KCNXMU46AZokerbvnedVdMDNHHtdAIwkHZ89268zYVWDd
AxitgXV15D2VJZh70JKhTkuMcIvLJQ7tnl+lLllIZa477Mhi1wP/yqado5VL
qeXIWt7+pn0yCPHIzuGhcXcuvEfzeZT1H6CZ3fDass52XSR5P+bZxgC+pwWR
owwS55qUmc2nrm25+ZTTDwjlkG0V9KpBK5s29+f2EAJu16rHNGloGWlIqFyU
nbG+42f8L3A5XTnVmty9aXo4mPDPjzIt7+jg+EqWxkXwU1Rb6SqY1pfuPIWi
nTM0kv4JWVe8gSJk4Z3jJuIqauPVR9FPPqTpACfonrqf7TFhyju8NTWIAK7e
exB5hqOKKueYarnqOAGoDMUWB6hqmizkfAJiN/qC6TZT2xsLT1oA6UCjQ4b4
3U1FWvIyErLgP33Mxwi3n0ZkNX6X/FudZ2Qg1x6bIN9U4EFzT2kZKvpQXSk1
V7HrJSTLAKsXsJ2345bYEWiafbGBXuvZSjXMKeJ6Eqdc9RXSoyJcLPCOjARV
u38uHecTxMv+4suaD2CdPFiOkgq6ePwI4Zp3m6OiytzKJMmRY78rdcUg6nMG
QtLu6MKcUf4G5BgNPgtnNLH14alYRAGvnABDGdHsNPC2p0IAlDV6FwKIa46c
jzEDgzjcb55vd5M6+sgYtKu/VKhBY8x2RtGtkoDZoN80t28zFHFinTH9pDrd
Lur6sQVvfWlyl1mpoqnnrZyLBc5RZnLtobtDTauHDUmBD6DiA7m/F2zvfL8w
Pv6nXYYUHsy0sDunGxSY+hqHYo1FcSIV9+Bqf59IH8W4Puj/Z36Cc+Bu4tkV
XRpG1cqXQVbHiNEnwynUSAoCbGv80MTfJblmNTgUTPizWgcE9tRFbR4dBB1w
QyEyvrhsYBKOnozROxmC1Mg8m4o8R45ssrl9ZvmILf4LwkH85IRErBDumXSQ
mIbpBODdVfiGOlWPXirSb4sl5L0sI/QZ9WULssaqcvHHwNfZyp4am2iFJ+bf
twVOYANJiA7RZtbtGBMdtxmiER787deodtdPlDL23M9qqHwXrXf3q4jSabQN
1eogUIXrGahycrBhLVxhUH7q/yS3YmncMeUovmq9V4qwvv2JlqSxpTIVZZC8
TOpk3xqnPzO7M/zqN/4AK1X/J56AklDIGNq9+gHIQu7g4KCpXhgB/KrsEOs1
g2SfQohYYH/hbx4mHtsr+GVMmGVMtaU6NXJIWcb3vdGIWGMaI23qUiekK1mO
dfoagmV5/9b3GboOuo1fGdSREvKMxTSnK3D6/ncKsDPtoXKdqf7KFNZOTzI7
ocplaJ9v2BxpnCBA4gfWg6cyCiXwV4TMZ9GBdKgPBMnfTSkzz2HI5TVhqZvy
0zxHoG1cqQar/pmDvlVgfI20zG007QK3toYC+R0Rdv4ZvpgJMCKS2tNTv8KC
6a8uhqucXKXK88NrwUYAiigYTan68yhk50yOOihvU6Rpk05FXTJfvkupPliT
gLUKwW0MTW92JZ/GPcgA0G3yzr/Qsl4j6KDvnBi84EnFpidVQ7ESMPEK9/JK
D74Nr7P4fJtQX+83i+MLt41aQmV/jcN9v0MR9UHP/8BUICtJvsSIQlsShsjT
ichOiyU+/c3MZp3zW5PcrJAWJOabjoNk+S4j5Bu0dMDP7hzGvAL3MLA++8qS
xe64COkL2z5Vu9KItZzyjeXaX3L2r9rBw5WFbot5lpzSR8bH1499gtxQHNOK
sf2eCC2L3cOa/g9CHCByI1PhXdmz9aOMg7Ofvm5GJAWY//CTHvxyT2Nz+pnw
+eyvlSwjwfEv7T/EhJA+faCi7Q6L33nbs6vRKjj6zozeWTgfpqUxvaK2Cs5C
2O9PZ3C0c4xNo0nkFjnID+VE0xM5vsguBmdctVWnNNPF7IFcJTSQosbHP8H+
hrA9kZAR0/id26sk7YyLUr8hk4uoVKagIw13Ztax6u5UsC7AkJtCfBGiEjgu
ECxm5fxSDRKuSpc3XT4yzSpXVGnPEc5W8JT30VDUxgmKaeo5bI/zNzkJQ7e0
MS4Nb7uW6YRhaIbo9ZerhHhvqJ/L4C4DiQrz9K3xuRZlpSJ3Y9KxUDZPFvam
gga39hhkHFeE8qJXxaPNG/e+rtf5fuCRyM/OK0RFSRNZDuTtd6iJNZc9Wl1l
3IGeQTOGSOtGIszSx8kbXSRQQhz4AD6JTfryd9N62YZta0QkO7vrRclM3LNO
ea+xRKL6HW8IXvVY4RnVwO+3xVIZ0ei4ndXcY5cmFnHcGxxnGYp3HsQeXOwJ
MAv9/mVKretHChqLAfSpZd6G0jiXTyodpTWaEamphX6mFzwO8PgkNJp6EbIT
NFdVYogbAxCQk6QI05HBlOy9YYdJb8OtfeKviqlmk+sowj3eSjXSQCytsjxk
8W/wFLV1uSZG3C1HHAEZLwFJEWwBbzQ3NH6mnd5fa6ZvbAYm4S7GE3NX/KL6
aR31VrG1VxnGDUYCXD/N6Tew7lWb396JGjTYSlNnHY8EDDCjUfIxP9QF9mVd
4SlgxxbiEzVi4APV0OGV8kgNrwM1Sf7gQFFiOHJ7vI8rgNfb+wYLgTYSGSxL
+YuGT11fSBKnsoZ2SEgX91r9QVjInN/fljZm4MxBTDuPDuAF2KOP7G7NqZvo
bPLUbt2r0qCHWhgJ1Z8pQ2xqVGSgaj61sCuADM7GNBOXknlVYRRvv3T4S9Oe
KZyYv2UdA0zN2Ps8lJnkrlTdWg3JwVjoYL2Gx4geF2x2tgzj18H5PeevheAK
A3k5G7pZ2oLSppKDGxyoHFk4TyMD/GV99YahZsi1bSCUQKdwR5cYSoG4GrK6
YZGqXIMyD7ixOZefChyf0fZCRPPIFriZAej3z62hm4+1AScHpzRY/fxH7qj1
fuB2+oH8/EKJavi2Rtl+MMw6VSLMOWzLk3iiosCkAeoanzRxdcWAsMlBZIX+
picf4OJvtNSaurX0js49WyAV0o+39qsqN+1jhommO2bH3aevVuDoXU9X/PaM
oSLld4B4qhPGbgEtoWhkt7aX2qRqiRCS3sJY/wBS9jPw9puFFZ38gA5Z3QSI
sC/DMRjYixCYAAMwrnLTdyqDEWE9WuyCX2Kh8B5jMcLOE0IKUAqqE0b0yhpn
pJF4jbbapqXm7AfGCDu+RoZWgPynybxzSOPLCV+lvHVmUSJ6Mxf40KkTstke
XPgLwFqcNMqrqwIKcuY/yzUoqOQz/bdUuo8hMgPg1bORkxC5ZNhPbcjp+/O1
bcyFMrwJDaAEu7ejjA6B0NQruI5jJ8+HlGuIv4FsOaIS3S3ZSST0cCuOCA0D
YX7GxMiL/0vd2apaZr1a2xRWA7rckOJMI9d+2SasoewW4ajRfPI/7pjbnZuQ
DwaInx5heaRoqeLNy3QaVgmAN/1fM0VLYshb5UHD3hUWY9ioK9R/r8QBkwOI
JX/9bzNWsXDgwHRZ/uH1BMxLqJUE3ozdX028CweZk3m5C6AmyjNCKxFQYGoe
l/K9X8WU5w5Aw2WXLXXJ4ZeuKaI0zO3aX6KQ4IF3t6Ur6eE1QLdYMzNHVO4L
p+q8br3zVB75vHqciGjUXMrjGHf96FumPch4HVQAQXhHMa7B/aYUBCaMAnnU
U4DFFYYXGDcToT9rNSdd4bFn1vvCWV2tadboeRr58X2d/aPxiAh14n3D8mPH
MVeVUdHMMqMgk40ZYdm4VltLTIsRlIenSFMr4dpQauh9D8EUd90+ca4BN8vR
5zUHdNqttMyYd8neDc8F0hf0jMHhxDAETaBHv7t0qpj7OL9ExOy1UFhOLf/4
/znpMDlfdvtPPxs3CHZoM3ZgStPCd4ZUNM6yqXoapZ+NHm2j9wQaAN6f8SA3
7wilHICkMTwrkuviim8Iwvnlh7iAjS7KCPWLF3VUXewpmn2DihmSVc8+3++m
l/Jin2JF6ssiNsJuc3UfLPoKqzeI3byiH+p6c72Pdt1Z42kky3di+ntL/oIU
OrqKgE1Ur8CJxgjdRTQoCO4NAegSt7axKDgrjOEq76yoPqDWDPz8uTyReftm
SxgLcvmYsEzBqTRkuwyJg4aF8J11AooqWFSKp5ti5BDG4AYOye0X5g0qpLxq
e1WPtxQYO7FHdPRhhHd0R8UhgpzBeRhJWY/JMPjKXL+0x2cx5mW4pqG3nUuM
uVhh2Sq8gSZSEMZBhxeLlV2NeQx+SBvU2ouLnHsgCW+ePfbj/nT+R9fJ/sCK
bp+p1zoOXpqQLWk7nWD7E2adz7PpTsZpEbAKIvW1MiFdL/ZalRNu7lYaE1f0
0YZTuXsAHSBxQDaNeiwa+NZEMPEkbqS1y04gr2NwD/SVrQOtqAA53RCsT1jA
lOw4YuY512EHnTvPPtQ4Zx3rV6JNSub3fNNlBU31Ozyb8ecBgTDcQPd1g6Hk
tgVZpGJyL8rmonHs77ZnrW2aziLOedlQVGhbQiMFOSrV8uPoZZWO2jXJoNt4
K4nB+szHPXNL91iNYMfgBlFFTkoOzRnTIr3oaz1jdfinREw8iaT4t9H6n4xR
lOHrp9kSVftvKsfT4yBGnK1kp3XaCv++zYiE9abLpgL+/xly5zkzMOgV0FQq
+zv91MpFW1OeQ55Ws5YdBTG5ZKHrWKuWs6sVqgkyy0qdDJYnnB0T+gM9L4ug
Aiv24SJFbukPIJZBzULiFW2bjMIa5wUpQr1Gdx4yRPjLfSICT0EK2HFtmsWg
/kvP73HgnFW7S1zgIuEShq3LmptpMkRbKosQr7IKQ6a7Kkk5lrtLTGE2H07u
TW0MMxiBJPRYYAdOFB/anIlJ2R2JD80ykGtGHtfcfLthb9passLyZuH3RLmx
dKwvUHcEeebrpXoK6cA5ePpO0DXBA8h/xc7KX+2w11nKsS/WwyilbNlgpLf3
bi0qvaSrOZ7ggi8BqDZMeHxYgHUxuCFvSVSjoVMTtABvOkyrrr87qGcrb90C
p+dFXDMCF0n5+WTd/sIrrar0q5MkXQuZ9OfofPV+jYvLIgV+SNMjE+marpwq
txIw1aSYzc3CnnTcD7NpO+7yEscsshNroyItW1JeSS48a5cvCm+ujs5ax8mD
cHekewX5NyPddyMyvu3YX9YRLnm9iu04B4qubx6ajevuqa6s6hFZu7f6rpLv
YZrI2eoMeWrO1aRAk5gKu+Iw+XQSD2CQ4nf3vPu7LxuCwANjRrOQpZW4h5hW
jsDHM+29lNKY/uO6nCIgO3J9MqFgbrhtNp/9gshTdhZXQ6Py7Q7Na6lJWbnJ
Wl0RLhxw+mUZrOm5WL7whkvPLJDfYUJabVBxGZoNWnOey9gcTFDKhkB1QqHo
59vWu0AZEteH+aEcEa5SyTUXK7qKM5yrTMdanCv4xNgmy9DYhwW9HjlRF3TC
hn6AzpfgZauVG7QD8XfC3DLs80Iv/oCnGMpY0TP9aNk3SMOObw9kk3cw71K7
79218UyeI+MzPJgDLTn2uwIsaNuCMKpmLQa12uuz0UkEJ1BSpv4mSCpxexe6
Rh4k4ltrSq1wRCW7kX3WkAsWSJ/U4oL3ceGxmy9Jp35Uwn4F72sOsQxl6nGa
rLLk4CwVHI9+dvHdyEhZ2UnOp+4nyHcoCwjexylLEayQD4n4vtsWBY/oK2It
Iin6beIVfvp+GrOqMzNfWr99UIj/aGhpTnKvyCXPPhYOR9RepDY+EUnc33VC
b6QVNT7C3fa9tJLY151w/J+6/4NEYoOgqlrUkv1GDU/KpwIj5s1ogFrqHlH8
ag+vtYNIpxSvoTovcnJkES9REpWgG/oMMVP0S+Uqn1T+qZb6wLniA8f/taWW
GcQuARdcNWBJApk30AKgKPye+9ZVlvhILCtc+Y2PElL1+4mhFDpYmg09cBHC
bZBwig7CYW31SwLG8/Bvj1C+Uc1oo5H/gSTxtO6bQ3axqb8Ra3easTwwQPjt
neA3P8jmusGJqQucGUMihgnMCXGon3DbZq14wxhIy1GTfn15oQxuBpSvaIzn
xExkc+MQM1Xg9RzNJSAw+UyumWxF/uPpy1h8FmDqdrmI9WMuKmpEkpANxWq5
QsPaOjqQ69Yll2hhoELLvchFgOht8wtn1ZUHvlT+xxFcij5Sd+Yr6IO6VE1o
X2ueV/CXAS+6uuur9qrArDx0cjsTjiEN2APCIQdkHEePr9H/NQ/KyP+TJjES
qA1Vp/ry35BYDLhnEECpJi0yym7cX6UefmCd+86h23uzaCpJphM6j0cMDTsz
CtK3ZzM1Hywg5wsKKPjPRaDm7t1NKVObnco900/5fPAIwDjJMS30vNx2/32k
wirx97NgVwMTD/B1E1LWgLsLNFBWgBZ4QhFqAYQki/LslfDKnciUhfvfvOiV
IpE9HI9Wp5ZgqjUstPLQX+lG9H3DyOIdwQkWOF77gaphgMj6pvldDebSnLWe
CbhN5rQCIAC9k4KQ5iKV6XfEZdX+za3FxEATAOPF9rbM58fqPb59FsveFz7W
pvnaGTHaog0l1c3prEFS2plGQTgdZ0f9zDR7oTEbnXDqeSpa4AhFcPHhQ3Yv
NvMVTZMyogne0AHAfnNdq7RgAwbXIkplZtHZmoSi5T8CqtxKH/T0K8Mz2k/D
3Fm+Sdr3fc9robRsT9WcY4y3pRIsORgmkY/uHYOaWHBMRIox//q7OqHnq8iY
AgKEP4mnMI++w88jSMkYlmsbuTo/oQ7rgRqRoT/Kyb1DOElwVCFAtk8Bsjgv
sLPvsczySV+1RvVCQvVgzOclwMyrij9j9iaZuOlCVFt+nDN8G7LqljzVKHSK
GjyNEO25nNE6xjbMbDlUdTzAfdqAYZfOudQOsApWh918wa0HEo4xvegJyljb
ZyHOmeroU9PgrxDVAfnbDkM1usYqW+laauujC8J15uIAIm68rUxsQPRCvaLK
ox7zmxXYZ756EkI3U+wmzLb9Bs6rgLZOWRnUBKZ+VX/T3ogoubxKgAxGKiOc
pqv+7SoWj1fabvl71Op31rfmBLRcZk5+g6npLQHyh3j/+hEoGe2Dew3w2+Da
GG53ftlmVqzHtAap29jKrr09U9P1HEAfst0nj1UpadEc3psDyd9HuFtmiLna
zNiVWCfeUFthbHroy+E9kXpNXSB4jsa0pzddmdvEs5cEYUWJhMM1HT2Hhtt0
kbFJS0bxQoSaMoyGTRo/I2y8OCt+A659ckO78XZcJj28ONq3GAtYqlIdLmZ+
9Bx+uikp9fIXbXHqMcMo5+Aq/zBfR6ReiQIEDUIthedxCUhGNRSC1zvd4Lbi
F94u584kXkRXja6PIiD8xnDZn7JJp8Fo2zlO8oR/jVeFnKKvwkdWpkISjYae
oMjCNGHiYVKYeRR/OzBKVdTNM3mIcEPBfdGYuT6lzAc2iWL4XHzTzyz2jM0J
BVhzRW1nFIxURRLUzEsHwkgys2014+k7/Nc8mtdj6iV9p0aPzfLsCTw57gpj
9xSLcXrykHdiCkg1/ansQ8sfyTAT3VnZfPOtCOU3uASBkA59bb1AvwmlMgkF
ijUwQ3IWBb1viV9R2NDwcMn9uBcc9HTikZQzM9K+shSGvGhDcsefxto4txPb
U5/eWJ6kPzompqPGwJGQqc2f6pYLFgsVbHQxbZ58Lhj8AH45A0DvUPkBu68l
M8eQg3pyFUiScXgM0FQrOPGC1eNWDc1wySzYPWGE04odRvu/q7aAVB58g/jn
LqoSjBa7VL+7hOI0a2fAlyeSf9WtGBLsggy+hvD6T8G9T2gfjLHR2SpjELH+
h+2ank6+mV1lhE4ZhFd3/9PdyUf3QRJ1wHlCXodins/gIEvG8qM4UJL+bdhN
lpuwgooohlBa8XCnSKPsIswsllXsePw87yr84Okevt7h6v9sz3EA0HWXgelR
yQFKbJcE8LYN9dqy7Mnxul9u11Vgp3N0MBOvbnrwy9YUhehYZWkhzWdHF/B/
0VYViKNto+pxcLBgWqL9fz0WtGDpPt4Gp5P7ZdM+0pjFuvbA4SLJxJBhcsss
IeQb2nb4zw5r7zcHNUJJUFwAXOR+iy5uE3JNj0JsOhCZspKVYgmtNVf+LZF3
859E7eIs63phKIypzJmu5FovOJkfT+DILMbVUlCy+XaI/4cj0pZuT74Dha1p
dlRTqmPf5zgVIXCO8415aFnTGPErvxC7xUMO4g64CjSO2QT7rH953t6q6seN
JGlQlekTPJFisByc3+edIC5Yw599jGUnohwby2rtXYoRq2WYg70HyFcAICN0
SoCC2D1b2Mmbifh7VydRqNa21xLjnEWadrn55ay0SIffAYx3EZsm17vXcVgM
JqlYmTEV8JzygCHoDTq34UXDz98vqTCcx7z4+A5YshgTQLSM5RD+4eJXAPh9
RVX8GVhb7Ct75VQMjuWycE4v2FZ+L+24zh9cy6WEBX0YNL833jOcLI23v61R
nL68ZrrU0+XBASJHOUCAkTAE/4okq9LfnIR2c4N1spMxHBPjHwDbQNdMJCFT
/3Y8wnvRwu9iglorLHAIaFoHtf9PjmyLBVTzRpVqmcVFmQISHr2dJOsv6blX
KzyvihG1cRySsI9T4nFK+RciVjPeY9bIklnMJnu0vvz5uSWjV59xqe74+rMY
cr+ovke5o1xrYu8Rad39fK+KCQ+fyPeIi1ZHwSaDjAMHhab/0bmOf5Ku+pC+
80NY3jC8Dav7Fevwe9/J+fKAq9E4CaeakEag2xawCSai6AMvHkLzhqWpAjYp
NKDfPgJpoxSk9fE3pSJEILD5LasvbsjY2Vzg1+bvLutu0MxLv52oABNN7L7m
aT2ko3YoQm/Hi98jTW4NzcNKMJQO27dFw21hHwa3MEkacyeTER+NAzAlkHf4
zZOPEyptcktcEknxTOmelaSSfqCD2f1263aGUOAOEXEIarwq+RA81uZcTNQC
Vsf77ffjFcqymTBf6HsBn6/RXq0aH7dLYYJVu6oFuHPS/M+6ISsl+6HOL9yf
8JVtZAGKr0Rxux78/M1a+BfBQDn3mCze97+uSKHOS5n/pN1HrdFamvgHX98p
Mj7k0euNs1qYGE2eXVxO9ONFd/5YKeP+fbpR2woi8aR5IjMXaufoJ0Bz3bx1
QfZ61qjT+7zxfCZtuP6b71Kt9UMTXyO61/saR+xPdFzBrvGNUIoCnfShAZKu
v14Zo6x9XLO9jV0ZuaFZxxazskOXqXLmV1hP+QvMTXkS0AaXKvbwxTPjZHD5
gHbtpp2YDV8E+ECCWyJHQlCu2msi+++2ViY5uGfudP/AToOVbSTrexxX4Nfq
Xb3N40hwAzZNtJnziJfyqxUxk+xwAJI6AYfP5XIUjhgeHp53zCK6eVElpXhQ
NUwyzkSeTWBw/QaiUcMSC54AcAWx4RAuOXl65MyQEXHV8ntiN1Ry7JZzaECX
jYVdfoGNGrtKchEpxSikq2JnoajAoQgjcXt7kVeiyrW1YJT6ZKZT3yIEh0lH
Rw9kfpv1WbLh7hALnGHfdw4U6SugUqvfUYtKSbAoV6la5UHPzJbfBgdKQsuE
EFW6PftKu0t2cbZl3YwO9wUZ9lHc1mpicamlreSCFLI37hM92TotenJQq/do
G7XmonQo1T9lEEWNSzntCa85dxzFONdNNse2K/aD/7k/cZfkwUyjX8CZFdvX
PMcKL68dD3fvhiG3ikEVDBJa8uDDJpYZDdWLVnboeBu3dSUAPofIorl8BxB4
ZtQQCXz9NSH0BsT4N9j/cF1jd5U6U5bxloKtya0pY2Zr5hspcSr8v+Z/GsSM
6wC4O5cmtBGjSVqigd6SxxeyUvxXPyh23RUwtgS40zT0vlw9Bte9ZRwbFrZl
+Ercbx/gLrPb4pBcXNKzHCj9M9Nhvwzwccbfz66G5dKs7aabvcrHtY1gkfU6
FaIvt6vyPkocZ0zVYYrw+ilwZk8b1IARyqqTvBJ4JGbIRr1AAqdVOYHDEBLe
2W24YkTpdlwjqn1yxlzsBa/HP9OdW3K7JpEFhvj6GR/NV+gULxgy8kh3Tw0G
IO+tdFhgnqLTHlUQY4AHqsGKxlMMHeuvW68yKIONN46fJaWNF2/iZEbcsn/4
hAUyHNYRg+3go9dZ0Zaecz3+XyEg212uSq/ylfpNKUON3C0dnKXCB3n5Feek
8GN2f0XkPqGVz+x5XvwaBh8PNwa84+h2yULAJiMhjPLkYGuSi5YMIqpE8WNW
69vvgeksCDe/GdzuRQg8atEN55q+NP6OWo9ppO+KyuHUSZ6YbhGqDRENb4xR
t6tgzei9mf8lf2RD92oxnEPMHGj3RQWmhc7LX2DFgSQxMs7QshiXBjeYO0MH
Jw3ECpmUwIibKf1wogCg056KrRA2VBlqMAUpanBQYcmQgtchfAKsAdXJ1CVl
4q0+bGQ4aCHJHrScmxl0gWlg9E9AzqTzD2RRPKpR92Lx34Z7lpE0XRgOAH5T
yeRcBojCbLmH8YuluP37S3Vn56Z7Rm3M7V1i2wmmzUDB9d1+kPY9zMGo2p0B
IZzt9iY5+F7o6OXCdHhMRoY3smHxf8qiX8ljfkWySJgxXzFGWmpeahfb+4GF
hJm+2GkIbvB0x41aw3SwtkVU/KNgFPk4X0AH78hI3I82phAOBWsldfel14dY
gqMBQTpZK7fi8fml3yC2Gy1elWZl5kPVQySnCynvYjhx5Xkh50zuKEhVEWmR
9zMKgfz8LyulzPT3cN5AjSgCkqtHRJxg3f2XfGP/RtrlHeDubWTEiGe1n9Op
dG1JkpcKs31jDBXqAR7oU65uK0fLSHudQ5wTgmRXTMab8ALmNBdpk8QaFEn3
S+hPGixDzmKUrXh9GIcteLD+tenm95lyNcP/IjDnz9++VKUlaL4bOcIKfGkS
uUDgc4VBQauTTJ/G7PeXXdfSLCo5ieP95uEGZRAyloUtGA6nOVD0Vu0j5Ut+
mXKGHdUoxKddbEwSIYlDJR6JCX9BPC0+8jgs0chDSGeRmFzA3nl5+BvXkJpa
++2/8rg1qBOkxeR/FkDHWOMrk2MB/1/wWOb5FOt7fDbh0Mnq0nCCewpaio5g
OyJeXaih7mxVEjVyZrJIbC4l+Yb5yoMnu1f5PHg08q3eAEKqy0tbFaYiptfm
SFm3VIFIKX9eUDPp6o2Qa5wPXyWfpULVyQI6QRxFNdr29WNqyfymL6n0g5qG
2M0PvgCXXVOQPL4OPPW2aRMj48gHbVXl26KCs1RZsajagpaAUpAdpe1PSFp8
ivAb0o/MWwl5SGDOn7bldyGnzkqmvxYTD9WbGvnInE5Pvhu5jvakYhauacLK
9T/XWp1iZ60SgA4ZmvsJQF+XaPoCH2R+NVNOEPKzJZbSRohKZNYRuLyHnTBC
+I4BJv9Oa7X3UPQop0Uyo2/1PUjT2OapwEQFpCAjIaECk/RMTnhfMI1z2Buk
mXGOM0id9etV17ger1lUVUYFvUABME23E/5tOLWiA76q/ob8t4yM0jOXf/ZD
5IzyX/+YRxr1BvV5g/kTECvaSpXJqIkOT/vsMUtJk/U8WSEEm2/fC8tT7ZyO
b8xnXqdySuyt/ufyoMdAm932yAk0H94LSmBmdzX3K0+AHlzh5ZxnGzEJSt7C
3A/znlZGikXeBVF9etzJ/+EKXJ4tSDg5vX3alUWlePGjLNE5POp61vvOj7fz
YeGhJgmRnD1syw16Jlm9L4kPgN4oDkTsBWo6f7ehLvdyTwl68vUGdRUq3ndL
hu3IiEKdVAjST4kwfxuODAi6x0Af0lumZkeE3sa/UBP4OQP02Ti5Qki0HaL7
S5eKFkwEU8JxYE0gdsvek2zJ7tA3HunQJ5Z2SK8rvc91/tHaQij8lODcmg3D
25fCbP1D33K54E/CgoWAqybZhgU8cUiFn8z3xEQiOApWVC23nH9+8L4B5FG/
KqAGd6K5Bd/U5binpzzRqDYzqIFcYZl9eIVlqPmi4rScwWuaa4eyTZDQ9nTG
bBx8mwc2a0a087oEN4xDeqNHsUyyNXySwOY4t+DqvisGb4kcsdEemuYn0wni
tCQR7hkIEQ6TlMqCyFthZ0LdCsLWDPhS0jXr5w+94T7EAxZiTMlK2puKDXPh
NuydK34iwvuBNdJIi3O9vaulHtX9HekuUSUUW6E2de09GNin1TuphpBWor6z
989z1rkjt/M1GNmOwnRdsnU94ohS1ATzS60G6VUVQklVU1Uy2PapWdzxsyOX
/MyTX2orc/zU7zSC6riwXLuxpNJkqjEQDgj0HUd23eu2epq1W7DWy5FA2+qA
aNwvUFc2elwaf6ZV8zsKtLb9HMRdPvYcgdXPc9r2fFXzIguOd+X+9cXbvwvH
iHJ3jZau/RzBhvEIz8T5qWMTgsCCWby6+S0LQjgzjLcg44QacJlrcmFAlt0S
wQQVH3VYlvlva5pzx08MJoaOQ4iHyqkB4Pv2xqWD7MtRK6jzyAN1bBjvMRr/
+pSE9qmgw2+Rtmx6+W3ByfAL8rGrRe/GL+tVbEdDTM8JHnahzzSvBkpewpPn
KXxAwh51bN5iYDpASy01YC9EVdR0YZD13tZfGp6YN75WyO9sdfc24eG/W8ku
7UtvSTje4KASiyHkbKQm70EgVTsID/Fq84xEcTjP7jV0ykVaeqhzxJHznmFG
hrclHqEXsRr+sdCPt6hkWhRE6QHenjOmPYX6t2lHCBVVJvsxkcRIMA6Jug1q
vqdV2jsArujjZ1Q+K/ITCgNYeKF/KSI6HcQr0kVdBY+FZQCtRHcXngi8ow7k
FQU0PQDitfEY2NKph1eyAIe+3KfnpCjYyM8ll0Hezp7PP1j/gNcLwtuZuLN4
KQZs8g/Ytp5h1FcDgT5U6FqCCYgBP5OgdOWgsFUiO9/+9F5j1P34LwqeOqfb
tGOTA18UNiuchXX0Gj8OxWZkI3TpUGpAWjAztXKkOi4iYax1hUHAR6R8sryF
zBgBmGANV8dM0cY0ufQbrPI2lImMySPFUhy+Qd3CaA0DsjH3cNRd8tj5Lcld
n8RcycgfgQvxP4Z62OWFoVgCsuSX2QNzQJ8wcltg5a/bIvvb6UodztSzAPgU
fkHMFGABZz2WBsNAheQhLF+jOFpKLKuJs74Lu2HLbkBY6edkMQOPtKyp1hnJ
UjVUz2Cl8GKfpOwfnvh0DA8PgNjvPW8jzMOVN5Cf8LiRAon72JA+uYWwHm+M
/rLXZpRKhgwqPzIff3nl81vRDedEteFp9i0SXS8rGIzuRoB3OGogQrHONHcs
c9XO+A56D4ZkOpPEXkW/MYhZEy1JPwjr/800u7r/k2xablvPIZohjKDWuxWr
a7BC41mzddYdHdPx0VuwXSiDtnCUe3DwIttwyPVXjytVJmPbfEfvcxDAItwG
bSq7tn1eDT1Ad7VcqsN7YsUwv4+kv+ofsOKCuZNvieGo7jcIUw9mwRXeE7+l
ScTmD9fATiu4HNZXcp+GUg0FHP12s7wgAy0/XuFIZ3sC8UQ78kWVzyRGhmLT
995NBCZtO7z9PrZ8+nO1ZgNg1YQQK17e9j2NGGQdQpyc7PjuHYrXd6mG+y6k
wEFx4vL40enB/aa22RI22zb7/4Dzl2eKkaVR0m1fvO7TTqsd9d8rZ8FJEZGO
0j5SlM6XQ8swRM6oTffiq7KNndJ8hbH4rgnse/FtQQnQ3k0G/brxEb5tg4OV
3vSVFKC3zgHl4F9W+NSPMzJvj9gn0Tbx1IidlzCY3KPgzf1wL/3tDn2hcxrt
n/iLjAK2gC6Gd9o/3hqwdDzAG4b1bs6FuO8J+Ul7RaUJDfXbyXWIw8aEGgT1
3oZyymu4v29yBs0KXbIWehjQa1PPjK+PIpJyfafhhltFRDYd3MLxEKSN/WkD
KEewyUGmCsb/jnmcPsnZ7r5BrpbH/JqHG+fuxEFI/QlAsS9/VxZBv2GkUo2R
nffglvW4vfV0iaeKd5GiKjbBOVG4dgrqZwCpgucYGiBoHdyy5Dtv0xabPTeP
BpQ8i7FoZYMvtdN7q/hsyblti6s7iWibfvDWIgZlXQDqe8uinRRrggGFDEDE
WfZ0xJYfvF6aBALll0B3+qEDVFlisUwCOTrUxuqC2d45vUQUMbXhRpasCSIF
XG0B1OnQ5uZ7FyliK29FEJ7IYuoTgENj82DuxCbGQU39h26DAsd3d29Vz2Y3
2WHVYCSJUwSWW5HGxz21lP0PEFu4Trm/4x/ocBoIj8uTiMfjbxInJW2dfhtM
ANB8AMQmI2I3sWiJnNqeMXolWaWU+l33rfQWeOyIWKIRR+zxhvKI5V+cYS/3
LBNueRa9etEHarMpHuaZa8Ngwu20t8jJ7AW4wnFWAc8eXfewQus2CORKsnnA
lfJtlONFx+25

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qQ9/kdbyb1LFLiv/SrAYhVILWSMXTS8auxD3TCPP9JTQWrpoHd+RxphpiiOfBJS6Z19G5Vt5ILUbZAayhX8579WPokbYUEHC6112ut+hNTszsZjNiBgUQT6zTulSqDBAfJMz7wGLQOStpFEeOHQs8n23svdxJlnenP1wtisFGF5ixHWRczk4v86MtZYp8kKLgy8Vu5vwzwEx5ScipAKazakvsLo3rXKrmPvtKn6gnAKwBNilUVHOGKV+2WYucLvePx+IXt7PCrAwVVD1XO4X7h/3wH++FFTzLBXA5VNqWiQjKbGcyWGU6pz8pSTFoiZScaePXYYRxQzf2tJ5nqanN4Wk7S0taHfGCJ02VqHORF18ALfi8H+Ryj6402EUq5OJcIkRGzeSK/WK5JFMUVCtFM884KHKI4auhp6BeFEiA8GlhY3gDWiKePvOX60UmKl+SY0xURk6g5prgwc49dE4zuUoe78YECZRq1JGt8+SmeYSuPVN+/4bsasLFbl5ai0puEak/tGTnrIS4MQP8T1yRiJSO0EpADYallu+bT4nNKu3ykir2Vm11+aSEwI+sVaVzP7zuiuoRfCjchfRqRxrLXQW1ouq5p4ryROir2TlYQ5JwzseJB5dO9ChcQXrXxaiIWFOH2IO1ZyzuTdcpvnT2S9WDHBE1hK2f6IJXWL9PCvaqasrYknKL/5KYAmhNTpRCvtpp0miwUJnqdvMwdi5B74ZfE69b3WWn2BMYiTxVHA9ozIm3/qEJOoqJdfOe8wwU/8o+bEzWuGQ0ESGqw2748N"
`endif