// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VFB+8Zbso31ztcXBFOj248npLxJGFc6z8khLj64btultfqyklS5jBo8txTK1
F0DxVECfdtbJiib6LIOQfiTiTxsXCQND5yEZwJBILWU/aXQ5EKjMk9OgylAF
RzEJ6rau3fVldljDAS6L+hDev+IDM68CeIITeExf8ruTj3utGq9D03t/7KcZ
Nk+3LFm2TSVHVbTK7zaT0fGFimMskl6JoKy0q2CHHw3n8NjM/PAncpZ8O89O
bNeGuYzIPtpe26ctgru83LOiVxGXz/tU2vvwLYrSd976BzxsnenOLu+r6oon
zxlg7ZDOYN1pH7on8KLoRc/ooPWpHRtOjUsFSlxLSg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
R68bmdWBKYfYxvX9NxM3A7AYVvPxlOSLX2Dit4NIfvJfhY0FB1ZWfnV67QPw
TDzG4X+plyZ0CcJswe375dEyTkShbtKO410rE/xHRxJWRplkKr3BhIR12hBV
vCv/80QIyvnDSyI5/3nMM1JjAOj1k1k0EJ0WbcwOisRhBOlfcYwxINRLL5xx
JulURXNSNJ6kTbnmwg7mBYoGV4xTamTYFGO6ktgW9UYhtdzcBj7ivNgop8Wo
OHMjqeTiOW+BOYig+ZFhr95z6UZZFYw4HnA57kpMYDRxldMSW0zsIBrCDMbn
kvu5QwgX4+JOo7AgiY5p+5jhyLACFqhr9tB3399Xmw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jhx8LVUPcGFCVuQTzPPxRge3bmBsQVSSHQY/LCTC3pd0KCEWvhtKB3xYHvWY
rP2hA/lug9w226jyHOIesnN35WJ0yWo9KKg62mzSX1LFL8qSMFDwtWNGwCXU
4hYP994klgmbqy6YvJsRw6iKTtHXzzU3p8jv/le7ryYgAVrc2IFbLutHGC5U
C6ut7h8wXTf1LXi4lUksAauIfEKGesspNP6J9gzgb8KedEvVxZOv9Emk7Ngv
E7088MOh8+t9WSZiabqJgiZFr7oomFx6Sh0jag4qisLnF+SO3tcTkm7CJCJ2
G+8bd4W50Y/vnz4P08lTKO/NibSTeXCCuFqDFjk+tg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oN2m7ynW2oHMxgwjSSp9rwYl7LGoU0DlKgGmw16bhBfH+H2qsAs6As50nOSl
8MacGQulC7StVGZn7uqDmzZHvq3qJqPhakr00glwvwPtZCouDQOLiSVTUZ1D
yFhtAyXc+AvJJGKnTqAUp1IuBkX7/KbsaB5wfwDz9qtbtxbU9ZKPqQD/Rq6C
5fDqD/76oyjJmcb1HR23zRfLvVifnvWeQvpTgAY+mWrahfXpHC5YoVMM3A/g
ZOriVJa7TvuxUjanPTbeeEH6LxOQ2kyWdSa9tAwGiX/ycfhHS5i/GhLQUpzG
RFrhZzwr/tItq50tNSYOb74GT7engOs/yr0MBAjJVQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jE4ox2qJI4JNOS6wmUM/vLcTr6BsLSWgRftrKh/n1QxAZNLtBt4RLba1Icc8
X0Tk0P99PiDlo6lGgS31ilikDfxpw8Gq9X9Y+l53Ueum/wQQMZJQIf+yg//m
bVZjHfGN+3GkGofn6eDO0MuyUYjt8II+02qc0fFKVuji0lrwgLw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Bz2Eu0dzBrHoHNp7Hf+6opNU811rRu6/G3gmchoZ6N/05hL3mjK3dczshsOV
RXEAum08NqMkDlo5pCsDbUHMlSUMIaKyEEm/7mBcJmC6KUVeR2VHYsqePTPH
iqYomKocQ/qLeo8Ss9MJ9ncsYLU13yeupiordIPIILWjnoXp0dfZNDFQUeUG
7R5Tw58fhs/ya4XFoA9wkakUGHJlZ7nm3IVNBPib4vrMkAR1jewTPDzponn3
NvVYIHj/ZjkKxDbKFNvmv/mOrdpTKv9mTYByr/uvBB/pXMzIgfMO/2V5EYE7
ptwgCSKuHEb/ypqioLQCkSm6X+cOU1B2FF8VM36ZsC34vypi0PI1z2VbzaaH
hMkShOzEWnqmyT0NcGuD7rCVT/GgQvqryUdjo6jQw/182hoLeaCBAKoR2AuA
I+kjtWfO2OQCqYtCrDf8XCecOWnhKhOpWG1yUL2XWUVyP/grWuCAm+n5DaHS
N/R7K4jDOdNR0PIcXWkrkK+qTPxFnhQp


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
h0YiM4oGCo5wuBH93Jcf7F5yBb0DKuhScuDkM6GUV6pDsWpRVxQZwP91uV1o
BIfmmmRNkdjciHwVA8MEPYPRvOWRac8CgT79lWhQIb0gDwsF5bui/UUf8jCh
2zB7hjVAP+cNmOcZjBGUs8psrhIDb9mf1i57t1xZMaZDBJjoqWg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
R/g7CZxXNG++56fUfOSvXgkpnKTmfH7jb/CAczVtxJLxrEAgVnFUu4edTKDE
EX9ItZt1bAm5pe2y4ee2yC9PkDGP41F6P/I6/Mvj2UyWovE5Br+hwjQBZtwz
f3yFqjD2L3et2jIOki1VYZoZ099bLmpgLe4idwU30dpBEHVVTI4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8944)
`pragma protect data_block
3kvko04XdswpUQIpL7cjYmUdhyM6njYzwKQq11hRJ9kKIX9a2nt9YH/znN11
m2qnkbxaigwwi2KssJ/W91nNkSBNHyggjFXk0mV2IUtNW37cMDUwp77mmZ+6
BwGGovrF1RiBWnJWwoxFVgbQSnNwh6kmPwJsRF9ROz200Z0QVw4AaZzIH9Q/
Vd0Fiq+5uGRFt+lJKf/l2e0KrLcqw7ennuLbTuoUOykayKvTyTHZcCqq2GNf
3tYvrQ9Ydpyo6Pjmo4IpGc3DRmPraEbxk/CdZDhvyW9sOoim9aSpr9ZFGY69
w/ntWwlc6B2fNLYlU6qK3BXdrJNBenov7ZDBXsbDrHtggDESq+9T1INXP+yu
KFsnFPQn+8AdGFwOpZV5eDCO6sgE/iH9bertFu94GF1sEwoSSDSg4b/7JjKy
523ZLzdYU7E81wVDVhIe0wPsFxZZpBj5awFTES6fUwuEkyXws3muPgljzH6G
PdX9IerjUYthZJyvDC44k125hs7TTFyQ3RINEEXBeEnBfUE6dRSD71I1X3JL
/xl8YIVkQRXIZqbf2oVcVEGLy6oSbYzxRgzDZgJPuQ88CXWq4Yeoisnh/0ao
PwiIaDkOAJTwIf3PwIDAsDcN/Ih/mJ8LDEbd9o864ExeMtU/HfQAlPc8OF5G
HTZfgHsnk0C3BAFOm5xBO2ZR+dm/NgedgO1u6Rlgo+fkScUFXqbt7gIiGypR
dKBO4ntReK31Mqzh1VmLbcq0Uby1w+QwyXyFkmUfJW7GsAOz5/13AZ/Rt7Lg
astcZfTFFQtPnTwmG+tdD4ttXfUtxaZzedCEez/XqNVlzwFCU+vGyNc3a2sX
Ub1nj+VtTSX2uH3wYZ4mEhtkZaWMDBta+Q6+t6BsM/vt/JxNy4+RLEex4wx8
W5BdVt/iA2whP7HkIj6l9VXhnOAZiK/T90dSB0HGSH11LpKignx3Ga2hT667
j8dv1OtQ8Mby2+FovUVMWeN1A50i2/OCkrybj6AMW9Xru4e6CXsd3OWFB5aR
2e3zkMpT1lIUHXFDJRYqOXbD8wjl+E6/0Fzhul7XHfw6gGGacKZbrJ/8HmAn
tDlA+lkXx1dxP8+pJH2lozEnG5Q7YiPmLWeXB5zCqiflTPRnlqntNdNfcRkH
LiLKjcePBgDDQdL7WtOs7UzGhsu9FCRbzojg+KJmDXEnGisrcPlOZN+dzEm4
WS5z0K9IFJA5iHoXrv8TSGVlqG8ZTuiD49vtqEuCHsBDeE6d/Nzybi6pEjUa
6Cx93m/tbQDiQzIryuTwiKU834N/8qhI7XrLZgIAm8vRGGe3V+Q8Ec2+YMzI
u8KwyqMINQbJ1REAKo4yw3muPwjq/6k2ovLxTKNMpzsrQHdr4Ayl7nNTLkHL
2xUKA+oc4iEvtXiYepw5evvOmE9FJyzn5uJSqGUT4lQGLnkElMKWUpmMNnP1
YsPMWLx0R0hBivHCbaFvo9yokRZtrjrZ8MjTtNRp860bd8lnOEJV5EGtXGAG
qDTg14cRIBX3H0SkquyE4l8ukDvoL+KXRhvF2WLsYG+stTPE3nUxuy83T9+c
dC5jRHJNP5j3iCKSGx5raIVV0u6tV20GPOSt4NjZiLHy67jX92+0MnGqkios
+W6Wzv6xbrRftNn5dSnJq8BXPuogQ+0EsRon4uFTRAvxi4/YnDRFxXNGwgcp
ESCqHgXSCV55XsyS4G8X6lSABhdCwEykdRWjNZU1QsAYg9Klwq2hsAQAFsaf
Y7bjvmTwXCStTxAunZeCz0psmUuCePsNJnsK2BUca8Hw5rAIoGf07hLeR1mS
IiUSPsXJF5TNv/NPQcMgHonMR3Q0QGTAaR5+jf88tSew4tSjvMsIgavHY2rE
JnM3foh+K1udpkRCNx9efh7pmsTHNEEYlp62hQpDdDqmWPQIbWXDkB6Mm+Ij
C8V2cvXOPp8Po8FwktXq7M6K01+mQcQqDY2jKoOVdNEmVxfhlQ6II3QQxH9z
4miTi5PC/8nHqk0CeJoAw6v03Y/2pYJOG2kSFg09AkG5gtdBDcx/otEaieGa
m4p2VWwG9kuf3Cj+TKvpObSwNYhuHvqkdon5k2d3vZnJa2KXespJm+ODNM8S
jYvmIKorSltxWhIDurzReUzv2hdQx2R6O12YLWLM6LeJJIoMU0tSeVugYBzR
2WIBjgXJTKIIvWJRwZ9Ddn1wl07iatOe/ch2Ib93Nlpn5piZcZoazMVXauwx
cxQVjWOquVGiY6FD0MFvxSPcPrUwWO1AVy6bB/17KMTVHXUkndEC5EpfAwZI
ZJGZxsB3/JVPjdrCU0sz74aTLFzwuo9JetSDDwYP3P3ZK1JjUNG4NPKMW9Iv
g3lFdhCULE2TmRIBLfcRwd9FePNcHFAgV4B05YLxjTVhF4zTLCHRa1b6XpvT
rugYiYESNIwSzwDzFBX4uokSfJWkhHdWQPhpG5o2AnAHIan5V9OPr0baK2VD
S6urkP7TIvHN1fZGqn0+ZN4XI+2LBguuQjYoCokszsd7rXWp4WJMgS7tcWIi
0ZERQPZu6f/2Y/bhK45cQzOE/R7UWhTqnPv+d5j5r8cG7T9FELxjMh6C9BUv
QzLBgVlrT+tCu94W3AkKGphEalDpcxEKUf/62oS09KevFchVjPdrrAlenyvi
/Llf2MKsTqCoeXV/7xl85sOVS6KlRCg7FOVT6HSNF1IWfCZ7TaWLwIqsBqEw
V/C8A07BpC7l+vzCATz6Wro/8+gO4Z3EpgGeWzrwJ9UTxbmHYvSjEq53SOcJ
iwVQJ9bFUUlkbJiNXlmm4MCZB+IDUksfABzyEqk8U0OB1pvC/avDvwg5AUdq
eZ4F6OgE/K+AOYmwZYA5csqd557qgXOoDnKTg73GeItCoFeKw0cil5ziLWoy
AuiO7VWGg5/s0kjxnA6VvjcOxZ7qV4rOa5R9xLk3onGhCsO4NzgKz8aCvx7X
pboz+tKzdmjDtDe442gLZpNHa8rzYRI+GJbW8v7pkVIY79k5YGVy8aRU2bh4
8AEiRbNotB0h+n1mT2yJI9JB3s/vbT2PwW0o7MYrkJ8fV1C/70rXBmeejHXR
gaRY9Ti7mtGuXFW8FhY16sKNpEsGR0pjioweTD0QdoCTfNc5fQsq7EY94Bsj
MXA6uablgmDuN67rX7nusK0ruxAplFLJ0RuJQzz7Up62UJvhI3xgG3riflkB
NBVAzbWGOY/1j3tKVLcZtm/MymqpNxkDvrcCKA15WeILc299uoFIssBU/SnB
LeHTZdnN/pHd1DWXzFdtV+KDhLpDwvklx08uJ7ZjJffHqO3j9J2iZvSjdj+e
mfHcAF/itxXvHKwIk+wcxP059BldETDLFGBXshKF8d78dEsHXHVmuEF+Gyko
op8PUTTu71eKTXNxZnBXpU/Oexk4tWM5IRZSVW3A6OUiJWVeQdXmt05tXM0s
Kz6Ae54rtzSc+LeRhL5+3SwcFiPEXZNuwHkcjGABBt7rdnOjkMVBZnYMtkaQ
RLCmCT+xrSDOg0flSNeL2MaEUaHmDtN3LaXhevhIzTIsmX14OpGbEKW1HIcP
/0vsgPrWA9hQOkucNrINV3p6uaR7eqqU+WpBZRUNU5Gybnt6n3tP/0A3R9fL
yRSLLdLoSOYS7+qNZC4cBOZD4flxDvSFKrz1fUicXzzSodRde1dEmMqlNW8R
85saJKo/fy20f73XxTv2VHwsgrjd6nWi/kGoPm+UmO68gCtRzpIYG37ZTigr
S9IQAuQQXnbY6/C8WjVamzq2HymlVMDb6bwxxJiQmegtucRcscrZT0p1LzMY
zRhphP6GII2guV3gUJPY891OeB4tv0wGIB85hWFEIMLlS+ylgB/PIbfciLzL
OkCvAV3a0wJzJPEUW+/rlAl/JlSdwRIMHG5Mwf18rbk7pWp1xrEaDZKTMxYe
OAicjZ0OCS3Ps5WsBEFStsSoXlhUZpdy2X5o0B9e0/SyuA6XSz7ReTJUynlU
EkKzM//wgpYIkUdLayvW91O9vMLzlLhDlF7EtJQdeb6W6+Rw1j/o+5fEJ51o
PXE6sBEvs7l8BrCyMtl/KMY1LDfn/pmo5PnuOoaaaD1A05c8V2TfiaXIM8T7
F48Tk+Omoh6Pqs3QGk208M0uy9zrcflYSqRlHmGlMIgEA132EXxfjG8klg7y
vVkadJopXn3jrWVjzu7052rbKcsiBAj8AYkz/o5vlSBvdGa/cGP7b3Ft62yJ
h3lKKlME01A6RW4gN853eApBRQlQAAOhEDfG8zF2I/73ElxpTqeonll1Ol7q
x0CdtpejXasd9M8z/47cgDrczR1vVmCQYa6tmNEhqeekA9oukB7EzR9UCyqK
F/kiKRJBXeXenjLDLqc2TQ8rb+2forn5aZebHMWiXYLML8lvTZzDVzw0bo0I
4t4zGzxD3tBH/s7VwSDlQLUoYv6omz9W+ppqJoj61PRXSPcZn8ZvUZ/T3hrX
mPt6H3Ftsd7sGrfhaGNXL0/749S2/V6SzfFZEQHsbOcnSJswsUkx/CSKmvU/
hKAKWn+CIMJFMHNBVO9HEXhcZw2QcUl8MuPe14J0ETNQWG5M6sjCFvuu0NH2
OxXwcG15Ft110sNGsVaphn02scB2VxxVtbAFe73tyjstb7VcmZWQHAnijAj2
jPsYIKbfFKW+8V+lYq5WTM1HWRurmjJAa7b3AenIsjr7RQ/Osr544/qQow8f
6pSiQ4ymjig/fop01d7GM1MxyJDs6/F7m3WyolJQadzboht1Z1qzDmNTfI+y
e+Ms2MZnYJyXEeOpN7P8lhCPMZQcP7d8iWiS/t4KxRbmD91HEJjULrsoIwOn
e4UWGcvpcUhKnI42cZ0IxXHfbI+KIEw6EYHAyAV+vinPQv/K06+04ghEzA6M
8JPMDfgtZr1VwAG2Hb4985YARK18aGtiFs+et6yDvFr5gkNWFDhduZWR6bP5
grmUCxRKF3L02wwhPvJKqSA6ZXVh0EJZ/sP6u+qEO6Komg0c0mjwghwDWq7r
SuQyh9ynSBodVTAO8Uf3s29wn22KNvmI6AC7YjvQd9sK7YaIjH/4DQSVEKOA
oQTBd0XIdf6UvJHC4b9khe6K6eP7RWAkPKgbUayvSRK3DMCkvhnzqydtB7Yz
vHbLcecVFkvGwQ0Kqv65qOtjjLRghWCBK/TUYlbxw7F4Y32we6+AUizhn3hZ
RXOQeo5bL9tpG4CQs9OW3A8krjfrTC4t2lmjllhE1JC2RNwcARdi0RpeP8xm
I3QHpHJLQ1xsbwSIdMx/QZaChx2sYTctIoC06ysdZG/YtJ61p291wzLfNPEp
6tkTYa1nebQLmHj6hiVJJWeppFRZU0k4h2pHm4U74XlqcNhrzLdJCEtws5qv
6zI0cfzT9XpDg+a4/H8rI60yCEn0Islr674u+4jCoZaUaJ5UeFIh+6z1prEd
eQAqYgVSdDhtVlD4iqxnq29LdRpxJRly/3w2NXdNDj4r9GZLKwzSkPk0R6OM
uv9pIheK8P47sXsiF6jInseeVES8LT0yoDCo/Mhwr0JbWnj7bGKzQIloIiy4
Hzsg16z+e7tL7TU98H435gsFxgniJrY1idx2D5i3Y2TqelVBtrGVB4aPS2Ga
Ii9sJo933vPWqcM69eB+yv79gZ15OQXTfBErqW7eaibPvWV12E/t7dC4ONFr
6qhWUqZdieY0uAg360+DI43+gu+G5CoWiyQKFzCCMzcPIJ5kH/rfRLt74+Aq
CKHGAwOVHNyzqddR9deVXolhkUI8xwWew/BXujcEdcfwWR5+rX8Z3J3hak1L
J3Yu4wHf0kiSAKPNn9yu0FYizMzcqoIw2x2LFXlEs7Hw5+iq1m75/j89/FeG
6jGWogljR5lK+2cGhMFvyAlxXxr4tCKOsVt1Wtz06PjqruCsLvwYc9nzwDM5
9IWekmbbXl9gd9vkiqncnI4/wl8ObehEHtg6Wbl653ydvANWpxv4dFkGYYYt
4+sl7XN9xygr4kTdoknvQ9V5SUgqVnaev68sjwC+PwvakWuBwVM+xF2v6sxK
TRCJMtHK2jRR41RUcWdKzVWF7E5dsh8fYGUwT1Qrg0/u59+bW4uFXyauzgWd
y/ypXYKIUc4aSY80AIXZzW2pYeUTszEkkj5MzA+ydo6/J1mqOtokhSbhoRrA
8wB4v/IGxem/kU8ashVlQ0XeC+/JXSSljrrg/4N9U7A/fh/AAPf8vFtN94fz
oDTVTDYlx4MJ9RCXq+ErCHwe5cJa2yRhLPyyf9vzU6Nv0U1KV0K0P6kiIOh8
1nVQBzN62fUNs7cZLM1ZMwbElSdaw7FHrMo6V4T8Bxx8gIV4hF8Ngpgt+7IE
59iNyTex3uUwAQCsfcXrc9cUhGk6cwyqv8LJsHtL8STmn3in1Trm3SUTy/uP
Y+uNz2S6ggWMtQMwkjTwRMtJxUkgCR+Bx+Gdqi7aWq+nxpNXtLFMmsqMfwF+
xs8twyiobzezMMUvls/WaRQcBZJNxJf06RJEa8Rek+FHPQJqdSQjevYEOYCi
2QYoqWBC9bOKzTNwHY8E1pZ0DXjOkcHAs/r9jFsn8zV5R/mpCJzqKVyPnbqK
q08EqjEW67QVIQtMjaSwKLneSOsQ7XXHSk52dHFqySPNpVr+elwVOFY5HpSe
LkQosIT3noAwlv+zZz7Mkj5OC1byDu+3ilq2OfYdciHU1iK/JxOU5K7Z+2qb
iRl2F5LZ7s6LFoxaVehzucs0KuL43Lhis4c2CJkKQyswZ4pTiGhSHJTVAOTS
6EJjtGhWQbZ/U9GfquM3TLmeWV6RCE3ubd/uTiEhD5bHzTaLBmuf7fIJkpr2
fstakyeah5EqqlBLqIFPk6vqqmlJ+SRKMvK/1PaltidD6CZgexV3EKGzxv+k
6h/uklfhv1ebWrDwEl/w9G6CP+2aHbSldADROyUJymxSo1GOMuWuzTxH+nNl
y4w1E60E/lEDQQwYIFGRBXQaZZ3UNaZsXzVhBZMFatiofv23RGwuydXLAmrl
DzfvdmUXVYHOPzyiBPiZ6UBvv/T0kv6BlpX/yx9Z2/Xwz/QNJ3L7hG3JsQQE
ll/feK6RqRUa8J/jv0vR17JXUbpKw02PB9RxW0ZDRD3eJOSXM8jcYYFAZrUr
Eh2SgkLRV67yK2UjOdmc+cWy7jQ+cmzmxxwoPYsJABLu8qLftTDl6R6Iv241
be7trXN1IOhsDYGWq53fwyBZXyuTDsUAzTYbH4L3bj0OCpZ8/Ztt0iCQVTN+
LAnh9yx9QPO+d1+bwdFNT3dMz29iA056HBAO4gjRG6j62SwRIF06bi8yJxuD
MX2OGKCPZcl+GRoNcjAE9INJwE+Uqj/5ymFz0V6lbaAYQ+pxCqBtXCQNYL9I
VNvWZAlK5k+Z+vFNw4cBFFJNaXGVCyUyTaQsvbVFcMTLteBYYxMzbH8NnSlR
KfgSBcW33NSevKR2Sru589ghv2ObGYsVLY8S8PVdoL3HaUCYcwjJfrIEKTMi
EnXI7T76q3FHvFHXcDZ3C3fEhV/oE7SegK+zD4HM8wW2SQZgjI6Nj6w9bqoC
ZLJbp5fHlqtT+GTzNMxyrIfvDCu00hUsOpzzIKGMbqavjvQxV0Dhyxag/Jm5
Sb6wZzNcZ7+hd5Gmb/FORVHtEFkLZRFx2yaPF8DdpR0Qcx64znBENlJwChab
xg6AuRrrgd0Dq+C298grv7aNdtC5to/14cwhlKc3SJOQIAOKc45O/DsNXSez
WTH+XiFcWsqvIgltEUJ0rm/AtrlbaPtAHtVW628ITNWb1y8J/G4EO3cTC9qe
KYoMXr+bebPbCyDym8SbDuMgCsBpMXr9Eyi16BySH4gX2SIqaWjYq7GgXWcM
FtKnic7EqdLGbmHB7secygrxRf3nL90cnEmmBF3IoCHx+3hxRYOGT+3PvQeq
vpTZjJldy10L4HMZSPTPFUQHZi+GmKc7Te0qm6itFUbzInBFL3UevO8AdNCm
f04JxljlVwyXL2OWa71lWPccqjirFyFIW7E5/lis37EIY+Oa1TsSTs0SrIE3
EP8mMK6GVFyvY+g2qqmurrCW3ONzOVmuylnfgwyJ+ZBBUL4+9noacVBG2svF
6pXyayzrangV4Fv9rKPM79hjJPMlz5brY9jZFZb+l3L0ShFRzg9lvok6/jbN
jsWpB214nIGOU9iGMDNk8jhMmDJsffeTmsz/r26Ezpv0Ruj6dbwMkcd2At0M
g9TlTecjhoHqcZvOmEXa+lSSZXvgu00drluyIn6PlqQW/2d1DPUpt8DKrkhy
ctBRSgSOiEq+pAC1wN0CPCUf3eVlPBQ0nREJ4za7fusCY1qYFzP1p5bjEJRA
SDtv+k1Eo2jQGzoLgNZs3AE/4NoxoFd23v3kCCZ+q7mJhBee8A1k3lNBoKfZ
QoijFQ9CCcpUfb8KhTdzAI0eH4t34uz8Y/WsJcpCs8GhFJ9f7kHvDzJlbHxt
wMY3C4i7EXmwB8rmGgPDVwkTw1eKjj/CZuW1s8ezHyOt3NQiUN1gXeVVlHKM
Ninn9nMLawEomhL6eE85hwlMBUSr9YkdsFdHCUYPslQQ5+Z5UxEf7EhpsL/2
dZAPFmuWotV1tr3clvwJYeq5ZsEb+aY/C3s6QvpHzceBV93fEUq0PRhQf1zZ
7Q2/bXRHR/ryobK4d9BvS2LIRy5+UeiwZTRyePybBx1RQFYwh2o26ktqoHEz
pC6DwXkmr1iGS4mYxOhaPxSZ+Bei4WL7Qdt+L5vjWc9E3OED4KJdfiku8392
tQ/ZcBL4lNkomnW7SdZDLxrsf84YI5Ws+s7qU6jTMIlCl/kBIXejJORzRwhK
8kfM/ExGeFLBTztWC5AjGF/fxR+r86mgqjTe0lTGSfoTuxmMwOKj12/5PVeB
Ih1mUP1EJueLcj9ZoK0bRWgxbwfu82h9KacJEYOyX7ja+48V5QZmEcNjRjo/
dH5lYYF/PSsMzYPvZu7gvNozYKcOr625LngVteZJBsLntRdje4ZwFKQWf38F
6z13qkT/ytLfBatY6x/jbqEinqiFC2MkPg9426a4MXEsUhTL+JtJhC+0N5Rs
OW0mPeBlO85PWmPsTiQy9ENIPspakqgHr7TONBbxPOuNjFBgS53jKKsgh/ou
rJj9NP+LsVR67cmpXjt2B+opYKC7eu91cv1waFAh/c65bpAgFTLWYeBP3rRK
EZM0s4tF5Fsd7rojaHy0/ht3SY2+nrzdIvQxQBvHagV9FkwtE4ISOWHPCh3H
7CFfFnXmvVZcFX2aGNMcpliWPXm9CLhVWJuL2wCH+G5lIx78TprDfTGgAeB/
hrADzm327IHmcG+biw6rk51GQ1Q73pYW2qiifHJKRm0F375k9uHggIribHt+
I5S9EfNbuuIADLJGKHgo7E4IReeheKG3gzeQWz/VAxT5DyrD1c1PIYLpsWPb
OgOEuI874XfsQIh1kg+ziyg/C66bHq+6FQ+V6vXe/vZ+xP7Z+ZbnkoPYcq6f
H+tq9SLYovcKWC/yjmgcHjEgdzMcS31a7KtpZmAstk41v9JKSHJM67wVabkG
SL08TZMkjNnjsaVcQ+nwMpPqjVPBeltFRncr236vs7NADquQ8bQOhZTbmyPv
zl+4txU6ZAe0ZORq8MPiLiZqNRqDYzUiKYCgsUomku9trKukt2Mxk7epm3AS
TaBnYujXoJc41QiB0B/6RAWuiUJknM/d9+2oSBekv6wTSFrb4l+qiiJm8o9y
yWi0GPg5Z3OZgI5Bl71siNFdwmVJKKMSiBqgoKF2tiZmBUVqhMTKIOSPcdz/
5k6z8P6VyA2+t1brDc/QRiVS75XB2/ecm36a6Jelmc1zkdIkCSbW7hatXzG8
AUCOf79LryPFCR97cuCBV1SrFMguNw5jE//oXYOW8aQoEuNO2ja6vPfzoxoj
zSjGLh7n2BPryd9ZOQ76bjkNo4TnBHuOhaAcy44oobfV9R4uMwGW/9PcW8+H
1tIEsBOSBv23BhO6B+qchshY7Mi8h4fyMq/k5WOi1pLmhIXuG9QMWYicPszx
CJqUAHd6T7mNLjpHLUcxx7VqNvktbOOsZ2Th9I5soUC1fEry+H7Mnltl9/QR
YCvfHPBAJ983zOAquBANPlVSlzlDvM5JPRmImFCtuquF63xc7lPWLN3QkfZ+
X8l5WhgNopYYXJT+tSvVeZhftElYpy8US96GMl/LUEhM0kTyn6WpYEmA4tqg
+0diTfEgghxNBKpIp9TXTpeJDlqzq4csNXDyBtvXBco+6pKIbh46nrJrieBt
wD7NmNTWjBnvPsI8rr/7ZXtai29vS3pyhvmdHiUrEA2Snv3hAzm9IgCrVREp
zyu2mH10byy0Gy09gaYEsx5x27+/YjLlVIoCYWcUXFd77CJcoBa8w5NjafNx
fXRPP3xlyOyOi39BaKYiPwr8MwqUfB0nNCNtZ7mGkacvhtMhteVqbkaIwmCN
KWdMn1Kcncxt0Bz21jLYbzuJcx71LsV/zU+aQVTzsv3Vg6DC4s72whBJbDaq
L1Im+DGYvwLWmn2DlayOwCO/sjObPEN/O1GSxrAdwFWmqFGExJt1pak6QoHN
AvzEYNLwZJIGB6DQT3j35BOTcEeyoNnbqn88PLtfQQaNHQ4H41X/OzbfCM34
Cri7cTCnBhqXeymyptrUDTW8c6uyLy75jIa8sdvrYU4PY3j1K8xW9t5jLj6P
sXfI4N8N8/yzkqQrBQKm9Cd60tpGF5u4eHiM1tfbqzHIcCSLCt19mJe3kTHy
F0pi4SYXG81LCLarpG0a3pgoRYAZTJT551K3aVjzqnSW05uZl4Papv9gSMND
pPgMdM3ruO1PCqtVnoFOZzJzdZmKGf1W0hS0rSOpn5e3cyUePFkjtViL6rfU
zWbrc9Y0H3hG9BGMcnvpfijg/WTp06V06ypaU8EtZPhkZS3l48IjC0KZgwW/
I9UqRIIUO4GtpZy2SvOuqgUoOSBD1ZfyNv9DwjWRZt42vxCgkURkySGFRUiI
yLL2BFNvmh1QM6Pu+BAU/hpoA5RxqhEHXJ8IguOQ4PIexPFoUFyl6cswH6fs
a+cL/CoYJai6d6/9s7jChSF8wqKr/rpTXECg7QN2UeadhJXs7Zs2oejJ+f4z
VBokxdrMHz+/DDw3UDwmfTq1PwqSNvotiScPq+7fUVnvJcgzcP3a71Kiy1U7
pymgatFE0KMUjePH4nPXC5JrXNizqoaxZknxbrTYDeYJNXnBP5ZFYfnLE/V0
DZCdkN+kwMt+646cj/f7N4lL+VWLR0FGhcV14FxndM5aShiUZgrjc10JdPCD
60g5YFYxTCodmRfuDe49w5P/3OgO7p+ayAJLPFiJ6gAXVHSrEyijpxiIXYBZ
/NX4A+lJLtlgh1cqpTYQPAjdIgv7rT5YQ2HHW/O2vVX4E72ko12nG0R+2Trl
cfIEa8EnNr2io+s+7p9OSQ8JoWEiuUsjbHwG2SCWwBqPVaMa/vt6eKvwTiTD
1QU1fqfdqc9nVl2PVv4xhP8CJm+p8eZavgq0jlTf7UO79YuEWuUkpnW/ItAM
mF4YKf9B21nEuxB528swcxQmfb3WiqS4+rNEBw/eImS3xbRwksjvxyn5lZUL
XmfP0kyPa8ZoqkHJznt3BAlM15LGPVJGVpAH0JtTr094jdYIZv8iSnZZnIDb
S+Uccka8+N4GXaql+2bXu2TB4JffWRboOjeesKcjK/zZW1uRQGP+AWBKRV+z
bu+ZS7tgKcLuWHFJxTVibcoTf81tfgkE19BP0VdlwcpRLAtq9tcZyowj+66M
kjZWiwZIqURcF9rxxT/BYcLGNF9aupr+kr15waTvpLdBT4C57fO0OwbFgMA5
k1UnDlTd96jqEHwWijOVf2NZkT9Ls//WXM8iL5tj+xbRc6s+PHgV+FwiGKmQ
ETnKzxhlhFViJFWSfB11hByXhK6E6/MvzgcNIjjOZw3axNPs+aefJuktKIQ3
SNgTK1oMdkCs8YGZ7Xq1QRJGcyd8iCxg/H3u9KWD2qyK3w==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "hmRb1hCms2kg5lxwgzvVC1ojkYPyZtVhUZroYIGDp3nv41l/XQfn8gMXcNw31HDDWBFvru7tQ/av+VlNCOY8CAEc3dS4tSN1iCLWoSLzjcf1An3u0nZDKunxPUWY57wMTkfTn6dFEXYBYGQG/cgNqAwhgy/sA9kmZ+yrzAG/xfCgRlDUR3RpN+hQPPycj5HNM2pIgRPAeD/5T2qj/frBFu5c2+SfDL19Hg79cXZFl7XTSKRAv84QoXAhg15CQS1cLdprDIiWjfSb64Bov4NiyBhMLbbHvh21BApIeMUwK4y6vAl19INlv8HZF6OCYFkaB/JHGFwooxyvzrlaPtJ/4s0EbHI7jWBeeQ9qR4g9+mie1DWbyHkC/cXjz7YH0auMBx2Y+dEMIAjKrUH/MAYUTJst3gg5P65fGi666i8zAgU5a6YXPqiqcvxb1glVL8sgBIb6cSbTadC0+xRSdvgYekcreeqoxGh+8SPcnzCfr92EMyjpohTTw+JG1GjPhIiIv3CJ5jsIdEeSySJCEkqF+AZVtjuFr3X1e1bDdKbDNL94ZSkTiGkYZsYKPjLTOW5WYcBx4HhZZgyZTiQ8Rr6h9EW3S4wsa0S98AANdeQSoE3uIp4HLTMD1+KXjT2dy7eD3VsmuIJB8AuzjVwatWXmIXQKFOCIMZH64V/Pv4UqEF+Wr1togsyhKAyVQhZdBgtvvKgDJm+OW09UAmP9/lGbHn2QvFcZGaC8WCP6qV7wEblNjfUV7WJgm1biyEErb7hxPsfP9bxVO8LA9PTeZ8gTVjSSHbqyMumIArUE0Spgd3MpBFfbtkv7FI23fedSMCNJCM1ECSr6EX2FHGTO2ymVbjJagoHYllQe3JvL6PXWYJmNm0vZrv6rEVDSwnrD+MXLokTakUP0b+cgUOMQTfsPZVbbeToDo6d+9AeTi9TK7H/rczT1o5dqY/OpJeQw3jG/DcwUK2wbk7afxDw6IXiAZ0UMypSUfffb51pgW2ht+zFsyYBup5mbCckhT4xLC0rd"
`endif