// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PSt05oeHDn8CF1I3OEsNydBV5DxQ++bpKbMR6OHzEdFVwDdiq2JVuit1xgDp
VZ8OD9Lq+L+26hAzPVAzyHsmB497McmygvJ0uFIPlb3TGg6bMWueoS56CYUf
mc1hoB9uN8i2l6pRNimp7mB1QgJeK2D/+VFpvaosCKhvxoMArzHmcXPhR/Vx
70wWpqDnHmDuz/ilgy5wiCOzW8q1GvX/zFBjvZWsAIowGHQicj9xQk1DFgpa
bylGmELMrmTuE4rOn9bpZ8aC6VwZPg0A3YjTFRovmk/yVccW3Q+StKgBxtYg
O8K3mVdoGBbL+ziwW8KrqLmube1/jQr7Upi9Zj96Zg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CJKFpMlMDYEcOIF11O+Ef3yBV7xEEKYLsswLFpJBevXx29Flnjomnyq2a8Ro
SWnH+fdQgPhfXPBT23kPSw95B0ZFQdOmeKZkyFyl3kAJaWTO2S4r+T4TKvKs
S0+w/C1mPoeNmdPzxDt3ZJowbjGsc308EU39lz+nTg+GtVfTp78frBjIBg2e
Jr6B/oScVKNH9A2tAgnhlT55JycX9/0Ok5ofw0OLzGOZBvg2yok6HBrAfg1b
Fc0RIpmLueuem0qZzQkilxDpHl7JgXelJqG+vMqgHSsx1alB/EILZrF9/Xml
pAW8agu3EgwcxLtZjq5dK8pxdFsaa1jFNLNciQ9RNw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JshaNchaKOUB9YN1beNW8dKvgPQdGlp2dlAe6g5+1/8tIy4b4jI2hRutZPfP
af9pW2Z0xxVi1vzPN3L5BjQllb42i0yBBHIMNiH8hhlzNAcl7+c0I/NwgDqA
KkcrfONcFLEvW5l/6tytbRzTfK7+8KnRd42yoSkkrFTLOBLIKJNUZyv/THew
vGeAVrHUPI4jc89qsCCr1nSmRuR79QwkzgfF+RkUZfntBdBiGitMLACVurcr
SlHjMIVL5D+wrJIKBXfVLWFk2z5QpQPPRwcjXRVROipgdYmq5el0M2lBGnrS
8cojIgm/PHYy8ntqrpYsehamK2oiovIQr/NvGOmbiQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Qs/6h06JOgluKQ6cN+wksL9mBPj1AhXQ2+Jw7oSCI2BMGy5PzBURw16jTcBw
FhdGAah8HMC18OWW2i1XUl7v16qA6r8K/SkMMkhK3yqZb1sdszPissC2EK0d
1IgpBqlWTRJOlutT5cxlkMPhmXQP9N+yWLIXyzZ+MoLGhcIS4DKVU3VGfzaF
JPz5mayO/XG10ZjOJ2egQTGG8oD+354wbGWZHYNoad/3uNVMF42HN/FPvEyT
X8fAbQrYEqr3g4IpSt9YHuCguOiTUnSaj7oe05vvIosK0b1KidYmAip0N8e8
XrUtPP98/H05tnFK7bnREeHlU78UUToX2Ygjrbo+yA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YvS1Cw4h4Ny2Jjkmgj0ChXbpKWzBCZfRGRoN7kJTfCEkEp+txCLauRMNH1oh
38E8K2syIGn5wloqnXWPdUn/vwKmdCrSB8kl1D6aChS9AoafU7nfL3imDzrp
oFzxwDSfV0lT9eqJH/e+KTpkqsnAicaR70HIvpW7GjwrSUHvJc8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
f41GE6NTfzBpSDyAiSY3sOtyXtiXuOGeyBEsdbFgyjw84H2hxWLYQMij5cVj
THeYZbpVuS/g91Tou6jxEwEHlNE0h33OWop8o0z/150p/sjOKjysMynowpVB
Pu3hnKOWfd7OvihqHc+Fl3cg1fomhqVDuRQ6o0eJ92BHv8pk+BtLSIVfKOtx
c0/Xnb8OU4T8ray/KLFNiVmcQqUPC3zNxq1tr5IHOSqVKsp60a99TZ0ueBZt
1H1/w/yNRMjTpS6Kg6C+wAPXo/BBNOGH+DBr2oICELlLNzcc3md29MalmPZo
IPQe0LPv0MQNFHgfY1llcRkLCrHdyVXU6dMhVlSP10izFAQvO70iuBuwKmSv
Tn9s58URP4SwEjxivjGXTYtCeY8yo3IkNjVF/tvvelndZrwwvKUYlOFaSOq1
XBk2Nz9vYWe1TBFHns6pxfxQP24CTYn3UM0ZgBeQtGmYcE5uhUgA/nPNqYAO
52jgpiHXpaNjDuEJd2CaJnc4AfwsHfLK


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YQ8+BnQhtFfLg9772PXXQ3/sXkW82rqYQ7hL/SKQ2qLNytRhXri8fhQ3mc7Y
QQfYPartxttW15tw9WftChtik8kN6nkIGGCSrL8a8+uCgRbYS2X2OAJr39VW
ATZ7ewUCAk8CzeCPzyT0qAxClxAaBoeQ+bNcfxMEm4fUKrwbVqQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
C0L61W+Hy8MiHi5Uv1BQ8JAfNa3tzHbFp99MQPFyLG+zZlgJiZhGL4GeFXOO
2aR6tztvBddmgU5nCrGh1Ca2dRzcM3zK/9NYX4hjcZ9EgZjqU5Dr6xSreByC
hMdtoit37NgrAoOPihDBwXgwJsczgQ7ttIysbcRObg9jTZ2zq90=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 44864)
`pragma protect data_block
pHJrGmmWcEOEy1V10pJVzLXEsHQBOqz7cmHK/+xLl577ilf0vGcfQMmgosh4
6GqrWwMGLJZaEZ/yyIWdtp10zs9ZBSDmmGxac8ezruFTiSi9eQbDb/ZhNxpP
qnQazYptCOMagBpCzfoe4UmI8a3/f+eHOQtyKj4XVwsvsfvxa7xh/UcjnRJf
LdOhbUxONmoodpkqNvgcYmbQvw0USmyuB+UcjJCnwFiZKbFrrIQGpUc/FGfX
UwwwqFmjNkAlbCKCW57sH6WgxRlogSxN2+qzWuFLGur6TsYmvz5h5TbRHq1o
3xVussZBoX7XyVvpo+y5VOEOevEV9u/duKlzCi+Si4Rj4PJkD2AhkGICJeyT
oZQMsryo6UEGJAEZKm9HKHDSGiWti1Sj9ZJ+INv894hpZ3vjmZPOTjvsl/Dt
T3UvbwtDqobABi3jfuDjY4fRGA8ReZPoilGLGXU5rmS8IRJ/0oLVKSsjYzPs
LtWdiyjfEhWUSztZnf71odU+3QWJdxKsyk3rU0/ucifJ2wPtqiTXf0Kechbg
9bdGEzCM1SRQ3TjWnaDWpBj7WWWzTvwgXBaJJcmsMYuiu1mLwlKbqiHddpbg
Sz100bJA3Txq5Ug+MoHah5rZVK0fwRc6sVvYt76HYCJckBKshmsS9wgIImWM
SPwx2Xjc64xA/Kx86CgbP06Zv01Y2luX5nepJDwyXuZXlvUopFQdw0Sw2tqB
Hr7AjhYylebO+8K75QAniwiZvp9g8mT1BtNUqQ5uoGdseyWE/JbmuzeiyWhZ
eM3oHUzZO6OY8zDeUavfnDmsU/iX5+FBMOf+0+B7qoibRLGvpukSEVTL8C/Y
qId2QhDrSWKENJwUY48sOjxwpZWCMpPkd97qRdtyWwGhNcaesOKRJOOqFBlC
MKiS4SfpjTQseF2BnvmIeDsC+40nGEOx9aX7nNebyOQC+KjcgD5rCeCoQd2w
+rFBCksNX0sCXTvkMcz9ukC+ml7seGdbvFwqOJ1AoVMtHTTBIGVc3dCcRoXP
e8ybrDxz65m6OrF5Z1wLcnZZY5We/9nSaFKCHXrw2EKMCuQR6Mz3/Mx51CuS
FhMK4xltvI+rVYo60aLdGCmNkmtwI0m9eaCnMpKf53Nzbvw1VqGUIWm150bG
MW6y7T40ohbn1EVtoEpV0DYHBCZVJwNsY2uvAY4/wtwDftgHuTc89bblFtpp
Um+mrPptUuVfle+tXxsECeC0rcQLWslsoLHPe6k48x6sPendp1xfMvzhvW8o
PIv2EgwcssBHlu/ErBa+1HY8UsQJWwejO+GAQ/YYaHEFzhID1s+3CHuYLKRU
tPf2aecGyHtO0BX360QbqFHZU4KwEIPnviir++mqw+LaeYILLN8PGMAP6UCB
hE34oyt6VmF4+Hn6GFQ6Lv4Wl2cGeoOlCiD5ZlMkDCRavcYOfI5ipc4fzgJ4
pigNNiZivNuhhXTpTDeOeZ9hkHN0hkSZ3mOaeZCYBbYvlRkDUefH2t9tAvBs
mrbn/XSit63Xa4wsn7X8lvsrfAH2hklPnqsxgUnnen9xlgEe7jLHEVqzG1pZ
LGvCLG7Ogc85JCrfr2EfDuLb76sXb81InIu0rvFeF5I0GMLnMC9qYn1m8ilY
w5N/GzO9NaDRpNICK4RSOjGd9q91+dRI0xmzfOi9+jjJ5M70vJ77f/v0QEKz
s2K2wMgYVvS15E65fTPJjjXe/UtYHl3KcU5lazYQ8gITUV9HlYS9hVFwEJJo
Xx39xtV88b5aHc0U/cY+o1DihV/aEdxKORA79V2wvB+CCGDtj+iM35CDzU53
t3uBIDuKAKtSHo82+rgeSCimVDKqAH3YLRh/sBXoAcVHlurBNNd3Sf2gHLgm
6nez2Nk8U8Su+6wH8zICIzY1j9HJJNiqbv5OKWkKZzwfCRL9SvMkXVQDbG8Z
QNO3Ks75PNd6xL/e6nOt5LAz3EFQyOaZcCoibJcc4wqjUJMdRW8/oYdZ6tkX
t/iwwsqT5nzZDdeW3rRgDswrJymCMp9Zlq7rJh8quTLBjCda6yD0Z8DMd2J6
q5W4zqMr+9UxRr89RIxAVUELhE5NOINZhx5Yzg1zDteeHtrNNKi0iqxCs9hz
cSW2phAc54FlUYFnl82X7bIKDJVaeRzStuqNKpXsFaQvS4TDx7cvtHhrGrb8
W/GJZKVlqQX7oFK8F8efkZqxbbrl2WbQyMqjCfI6nN6tlrhccV6ku4luWaag
5w3N2dKYjTdezslecxI2bQ28K0gLx3vypOzn2HQH1IfkGeuntxMCpwdRSySb
2AGochHKieLITLt146hFIQZrLbn9PV26XCvz485mSjYi3hC665PVsRdvURiL
JAxaULWWJN/30SPciKQKsuGxbmrsJy9H5XOKvhhdzZBrI0T4AxpLK7kd1C8t
SRElmviV8Le5bEaVWjCfqoMp+QoN/4q+ZfQopCjYLhRqsCVJE3SPCV/Tv3YP
mk82XWus0lyZIVhx1LutqMf9xs10FvR0VJ0XJ1NlEruJ5X3S7Xvsh8de51WA
9zv9bNGHLphCXxs/wIdSwPvz+wvUMDItkHCfS/b/SH7oY9gJr3Gj6pbDSQTY
JCz8ARe8ehoqHk4VH3Zo9dOJfbznyreO2GwTCJNpa7EelAAHeT6iDfDFt3yY
zr4QaBy8rrmgL3/Z37M3fWldk6T7EIroNuL7StH+NXHyhkrdve9xu8f2UF3G
7EvkFei+ftJm8FGYTfiVNXrU/NpjgR07ejuvgSXVU6jBkgJE60RN8lXv0A/I
ee9pWnRIkRArKUPfYutwLwDiBlXb446WlCY/aWi/QmrdWeNojZrhTFMFagCG
rIcawky0zJhLUqAZDJEHSHS/jEsbvmU+jqcvIlAxoxotJ/7zEO/eT0Kk1N9S
JYdzDkFSCTav3RUlLMh0Ka//0Ca5NWGfc5FxKWZqWQZGFtC1WvGMi0Hw73Bl
k/YxlKxI1PVfrUfm2+rdXtn40cqrNplhPAeGe5sAfEgqqUbN5ov1kj9Xyr3q
/V7wRDXA5saQFW/JZum8YOQbWybxd3zO7JVg1BXvMFSFeDCiwwS7AwRq0b52
y9aUzf1x2LwT9nzWz+i1GKo7CGgyd5oDBB779OXan3OORSjpkH80smK3ycH2
wR+ANAurcg9xOEk1d9WNNRI7g/Nwrcz7BLLAXU77NPMeljTCSNAjkbqagl+q
PIxsjP8TA8ALOZyJtO0PUbLH+UpgzgITwwhm4hTxENrCd8uBSjQM2EUbuH3W
0Yqv82rGf/Cjnf4NNNAJaiXxTrYpSbzcWhx0lXrvUW7MtpM0x8d1BHED55/X
CI7Ru1c+xYZB9DejXh6aneuFyLgjL1X+eITCzJ9KqT8Fehi7HKB/zResSPX2
TTthCkK9pcFau/FPnw+9a+53ItuNUN7QEG83bo0EGOycOY8ScZ/2XbvCbjhN
2bHTKFPDH2buSZWZCBSJLkiKysFXCFozlZ28wHEWpNKdaFOOjddLgHuLs9N6
s7cHY1C/51w+dcUqWxlf1sSemcSM5P6nJNJIT9vD1Em+9KwnyQYScs4L2r8/
vamPolIlb6FhJMKJ77OebSNyc7r5/WzKAA/OjaAsUp0+hnrkuA6+yEQA8BHf
tdzaHG3gLI7tIbHi+zqb1FXToNdUanblGTh2CJ+SFCXt5qsaLrkVbgeyFS2m
bgH2keiN/naNVEslHMTWs1wRhEqLhMd39WP06PofelmW8erDB0Hy3bqkhdOW
PTCHyhGcvE8ozBf6QzOnLBxorJLxpDSrm4E5hDNznnug9LOV3B8wZjrXzRzL
cvBkBJfIuWvVfNN0OMgxc4BjeX/7moCCem8qLbpJSVLGcPn9tNUnTyjueKEU
vVECCQrn/vAmt8+/w+onrV61apbjHMtxQAvDoO26WhGA9yu+BW2TKakIlbY1
s/7NW3608ueJ6639DexmmNhpz0yFvK4v1kuO18eh/XcUnDaQBNykDgF4pyBf
f5UKsnaQcsqfj54cyCTHkg75C5mAcr6M216IxMPdfcQefM9oXjeBCBHWuZCY
MEFaG/X4lNGIA/rKOvGDN2pBgM/t18tmUPgTynhNcOlucs80Nl+qxqQWBUQl
LShqsZowb7TGP5gZFI6OG3CiGho1IUQl6v2+rSn0Tjbq/Qj5jPFUg0U9RpsJ
NB3TAHae/wCWElmXlFo1eqULoHedRzktAgQcKp3n4LLx5lNhutBof495kTl1
B+wcXemsvbwPbB+X3FH6sh7Wmi7Kgeol5a/tK9jQQykbhlqJysArKrr5PtwC
sYQlv5Z6CvRsgdnkLIVFBMa5VYO8+Qqsg+p3QFp69P12wqP/2ZnDc+FcVBdF
7JEN6bnpJ2CZO4Q+2zchp7EplJP/lntpUYAQpU41JW+a7L4yjRHDWCSEd+ar
VGUNXvM0qx12jWrI8NKQBiTXqjjtOenpOl8mRfiYV7RCfuX8JQFnYcti6hsv
yJC4FjXfkx/nS2fOIjIk8jm2LBa1h7/eHiNJtjQSxb+XUJag9wnnAPrAAAme
/a2VUSvsTcU5jOLTqLMALHPH2gILmQToKS5NRqK0hf87mgUdkW7hkeLkUMxr
mlrLzGMEZcvMAkvsUwgBeTW7EoY2JtYwU8PuCzOQb1BKiaJ6yKNOFNmgX7cO
4S881Nr200PzXUensanj7VVXj1d3AdjuTQXViB70SUyccuE+X987JYI7HSra
f1rmhQg3qlm23TgijxcuJmg3nJ8xB///DCwKOJ3qPz6e/YNx8koeOx7EN8XJ
jhJsMq72o0NUVyMVZKQ3dyajCzPnQ1QFaNdnkdZRV866LYY5szAuKcJxmPxk
G/DxkCZywSBhDtaVD6xk1UnYavnT5BcWaNhbXVgu5uQg4GzMYXflmHMuIJ9I
iu5KUhLRAuOuEAfloIScvgfjVIL+VY4V1pvmWlVbdN0tglfTnJBhgEtYT573
gg5C61BffgOPK8Q/W6K7enLk9H/zjtDV5rtGwXVoDO+Ie9PX23NR+Vp/Flvd
enHXeTaAC6fljiDsM2Z/eIxv02jXkDfZYSHFIEtJiFh6+J6SM+0jlguXu4V8
k7cNcS9ThZv8X5kSWAo3kWOL3mpjA2XzFoDCTJbn5FDO+TTjRXHGTW86NIyy
cvuCueY0g9L/I6BJnA+6gYImEQy5D2RLqTm8FIBQM2Ropcwy39/jcFucNij6
7VWzbPgB/YD3xr74sNL2rhDZDRYW1iExm2+SBtw9j57Pl1Go6VyccujIMfD6
oLHcC6NXbkkAnTWRXhAQQQIGbjiY25lN4imTcBvmaq8x3l/b/q/t32P3BWap
XrfFLBRN1E3PwRSJnBYhvmL8HNXTVm16LcLTVb4T8jv8x8GPkg4YJKJvh7NN
JeOEOKazTsvUpI9UnczlT+pQwxGbe0Z+XIEPKOP4gydA93FDb4+BShYFIb61
41jebvS/s7ag8qLpwKx4ziEHG6uhtfwNMNK40VgcSvUfcYcpymqIRUgAAlJr
76D9Iqcdo7i67sJLR0Ds9SRo+zvnSL8MMkCQI+amb3nVtfPRUUsY3rpCJYVF
X4HoOFQZBKnNdxDDut/dk97cPnx7y0gF+l5MnD1rm/RRSg19/nn6HkrrPMUr
KIoUzFOuI7uIpixVorwIf9OjPgj2MJv2j0ZlrxDigIpGUhOAC3EQI5k2691S
EGjJpPVy4OwkvJ+M63LhtUqCBb9a3JVOID1QoFCGORXr+VHV4hwbtppVlMbT
JexGASSmhFsglGD4Dp6K3y+j1mhpkVLcat83retCAvURSqWA17OzCrV+zCI6
+3lYjK+2sW6TN5zCuh0NgK5/rH+bfFopAFQc8b+PEKTQcLpE5incPbG7fCFH
1/5nSkmP9DAAUtUFqxz8/atcAsk55uwkDifZj07ztWU7Lh6f9voTyWIt/Twk
3oEPdvKGEwxFzTL8Fh1yvKOb0DoRBKGXbyIOwxnatvhPRjb5csjMpds9MXqi
KrxPZlG893K4JRLwvrtZ9g4QpAnVmhY0gkrm0M0OCkJQAHYNf19sgAVCfj7R
GAjxTqneoXLQbfRHNwn0FDFawtBO9SaMV3EyTO7hqFamuSG3DTGyo1Rr+/rW
hh/IZc0ofr1VVd0oj7ab4SPAG1Z/cmTK91ugidvg9xG7j6XImVSFN/TLS+zu
ySBHPKBBzu4VQqvGbmgQxwBvtkBrtW8UUaNfZurwCTjGMaccSsDbO5fW1VYG
CIDr4EpGeTPp8x62iJsR9Klm4mdg50f04GTnGM4QfBpmbRPjRKNeSi5WJ+dD
+YvS37TmmlbW20W01lpw2mNg0jI0tHyfnRvQV2n3H7PqnZfEOXHaLBhXN1WC
DeOFW08KhD8Ii1pUAVllgHi+lAr39Q/q8hu4XReczzPeBSNXVH39M6A9UPFw
aoAc8bZ8DUQSpEBFcE6GD/dcl+jKaP5fmZNR59JE9N5vgveDfdqXVE+th9b1
I+kxLrdw/cuAsmLs9BZk9Kw3DKvGBYazPsuo5wJ71kh7WgJD/THO6lEZRaZA
K748REsYXwxsubVihSgLizoyT4fqlVvsmIc3pXKqAQ4pxCz5g2jhEOM1fXF2
GHNjpBDiJoAkXTmfvYkgJtzsxvLhomAK1FNtakJ5MD8aforzi+Cj70g/5L75
emUwJLn/kOo+iPI2cY4cpJ1mPPIgCWNuCYct2tx3cJpMKXq/hqEpUDQ+odbk
PGnYQl/k6Il+SRx+bsT1JZJtJIrNHeC7UNIihZH8yDotKsAadLy2SdR7eR+Z
og680x1lXgx056YBW1TZomFMnSgRTJt/+V4L6VsJPqeLPMgJKYDUQEoDJ+Cz
K9XlGAFhNZhWdF4hMNnG54QAXRW2xQxOs3VqCPwspapmUkTxDFzJoha8QqLx
3JcItUeskRmVcr3ALwLg6gGIEA6Qqn1FvvaXY6mJ7HExcVxC4+iNDtw7Gmjn
Kh9E4haakCDmWuSjivTM07cr3Y5HtcjaWGS9fun3cfyAtA7GZagfabmw+1Sg
ABDTvfhomk5QPB9j2fxoC9FLBVNvq749I8P32M8mLb9gz0r9FIK8wsBgP3Gr
ef6AI95pST8XEvWnPQunVxl+bJMPBb9nhTcWaeCBLD3vNe47jsm5jhBSxgJT
cEaAR8cWDEsVS9KtEQofakIfOlXqTdk4nMMH7W+7oD/vWVTwVBTfH7DvVO7i
/URKu/6oH8FCIH0fgdynaCOZQcFqlbteH39KGsBkwvwRGiSMYNlTWBRIOD5X
T9uwzArykM6rYACnEz/tfqbn+m1maZo2egBEgOHX4/UXMuMNfpPiFccJqsGJ
599QTimksxHBDxyQG8lrqKHOR3UegfpmbEm/9H+dOph2h5CwlCWNu+nc249w
ZuMqzAbOYgjaFk14PdyulVv8R6P3wHS4jf8n2S3JFfNAPO3eGO7WaOzfWwS0
4nWrGCV4NGOaGvT3YafNXxLWZhz7xGP36j1dOqBEo87wsVIK2/1CUdclNOCe
lvkef3e9vOHcjuAlh0g7jL78V3pCQNedI5IcNS4EyYrEM4ZtGYidzTZML0cu
QRshxWPA/Zeg5Uc+3J+qFJb4xUFxY5JrW7nZPPifIhC6jT5zF5kswHBQPWmt
p9ijUuNaVIKw1gIh0NDiP3VGJklJ8SO2jn1mREJ1izE+HAupcaTIPLadfomP
kjLc4mlGCRP8dBDn/+DHAVNxkCbdskM3qXsrIKN3LBQAS7Q2jI/tML+ptGIO
/BPYvVCGdXgPs6ltmBdt3MZvxsABs+xkUdtI0pFhsmRsc1eIsph2lXYnXGzL
hk3yK4tPWWBI1JICo125tlI6ZMBGMWbeSyrPOg6nB+B9iUVSZxFEMcjcZGRC
pG9grD3pZeybu0nnrPCOirTgMp6dCNbswZWhe+ea3KpaJduBA95pjrODKyuO
m6pGECBD7cLA6w+M6ujK6Qw0Ecq0et3Vi3H4HbzRX0PLy8iPINVpQCaecKEt
pTsrgEd6lhC/8vgckNH1I+myzVM94zPaSIi5/d2G55AmwzBf0r/THpBtPNfF
0swSxR5LKryGsVQlL15jxEu2YZZ+c6+gDSG7WBcox71rFMsMAh21HxcUrixU
Xjdpf5HVS6uAjKvjJh16z4/K8M8Q/o+n58XFlpP6JT/FNC70lqCOjfEWvI/6
UDzOXaDWB71a/jwCAfYcX7GwllUaOUQrPE3I50VuwyTSo9xe2xXno1QrQvfc
9DbVEEPwHvD5uRk4KA5MOFyoESAPFo6JmKqP1hN7WsZJlqc0HDmml/Kp1/KJ
ezaCs11I5J8Qc7mh3KCICnULr3M6BllSUyhFBo2UtLFnEqv4Egl+HgYHNy5G
80Wx6R+a60Lln3L85CF5JNAtj2gnJN8wV5LGk8ufWkwejROT6QkEDSYuR8qj
7iYIVhMLupmnKwVPvD6qpKYd49KsqQaRgZZbkpu+GwDcitCWROF/FF27pBqZ
iTorxPYxq5WeUXHMA4sECSNRzcMKV9PVbb7Oephi7zoxZSmV6ce5fkXgLK5W
iop+6eLR+dqUhdo8bZPpJ9VRGq4BWfM5pV7IQXGDk/ormG3nL28MbBIhX5jt
bXwNNUr7rRa7RSUw2IufzmZDzdOBO+L/U6ImsN+6Iqe/zKA4ZSYFKvHWul4N
VnKQXiUAwOHpJLSNAzRfKAaW8dOd5GOiBcZmXtmA0114Zus5NBxD559GD/NG
6hjTMcySU9vJLgnp1228R8/3e6aZDIDHmg8YCzHY/+u0D3Ad9zv58A6vZwGI
yxKKtVkpr+qa/Ctg9NlcRLGvMVOWNqkm+DPqeGJs42+SxquTQ61mQQl/q/Oo
1xi2n+fSY8jTJOuZgz/wLgwrpyzvbP/Gy9e83RHTmy1raC2iSQj95KHbE66N
x727qUzBVNCzOrH7oEjognUJ9SmxXN69J9xqMJO39Fk2r3JHPsj1mW2i9Soz
0yaPU1T9G6iV2jGlfpspckxfBAEchJxKAHBCSVVkHKNgIW0Zi+B5R+MU8ek8
EFy4jlQJik0fZGlGvqNspjqmj2NvZKxC5G8jKzXd91NAM6JJlGky7HjCtQQN
iL9CToB5nVKIY0ZKk3lxEe6Tk3Zbdfv9o5tofQFe0CVOTlOGDFbYVJyiW9C0
FY7p73aPhw1P4Jj6gVbRY5c6Ig+kq58XOKz72cPj81u/RTItNQR0rFNZaE3u
9OWZS5TB7ceGU33DmRfJRVFmAbY1GIumKdJk5K+/TD8AaWLX/oaIvrwZI2/p
mDj59PCWMILq53JyqnxMspkhVUWS6uaKIMEV2pTmreEvm/+PXmKDfPoGpLoF
I39/Nc5jP2DF+aValW0UH/xmuqSRo8OdgXi4NcBQ7qN/dbZk660S0pHJ6ocN
945Z84lZhOh3VDuhOilxF6m17SttZL9GQoMQM4gRHWpfEQencZ1Ub15XGz94
eu/YXxxesoJTWppDiQIMzdf6Pk6piLwe+BgWsnZyJi8N66sd65z7p74fRyIe
Z9JxwYTHjLRjdgdPa3O97+6KLbWc96vt4EBLRaaPSNX07vBLC5vTSgmqDp8g
RadB6ap2s7J1gXf0hONFtm9TWzgxfQ2UA5xYE3Gvv9/iFO72N9dq/rzuZOUf
fP0eJg0tDCKI306QSNcWjxKBgneE+qCtB0bu2Lodch6aYxHrlumChNvwq7Qz
EC7OTKu7BWi3UJYuucCI8fdNTM5V13bJVN/x3OTvxzuLY7sslm0pL8060VmR
MRf1TORSKfyRX8xWs2eMz0htMfkNOFkAtzjpbWmA9+8JNxn6UYfT6QwKgUm0
36t3AHG5fmeaEq7LNm0EoC/F950eCuwYAvUsQrCwFcqiv2e/X/UYKQ4nFIJc
M0M1gzAEToKkKPwzTUkFx2xwSAyXb+WEJ9Ss9V+QU9ERmFO1oWMBBw5mHQEA
x7C2UYzK6fq1JEfRtsH5+WKxYbvhUcmlh6ITzfZ5/ghQCvJLLoi6vor4aKi/
Dc6eaDacIga5hZcH+OVnVb0/TnuISwC5DOISaSzZA+cr+1kGKcsOsE5wBz2D
PwFdg5xSMFpqTm97vzF2a1gGH14xOCMOag+T2I/NuIGiSpo93LsZyXRxmLrI
ryxcFCHPj2xSeE1hOygpSFIKe3T1N4G0QiRnZKFXVzmh20o48hq48laqLM6O
GN3E84dvaTSt4oZKokRIr5eBeU1FzF5oLh2s8VnrqcQ4MOHRHYfIEuCQbrYp
fr8+iq1QuRgMsLByod6fdZobtKB3IaqcilC4qWxDzynK3Q2itF5mOuDJoMNU
Xf5ZVaPWlq1VJwIIL1bpmSPFwC3BCW2wgiwYnOY6Awlg+SONwih1egtwjzHC
LM1rr+bdUEikEPdGcKX8cLIp4zl7Xh88/trV9w37WiBnIIVbztNjlUgisenc
aWlK2HtEfKD5q7yVcSkB/eq6SsrhkjKyH6R8sqEhVVViwFyPGcUO2ACBWx3w
6MWeLx52vfGQ2dKDKkWuFZEtCxehAnEN5GRzZ/mRWdPtOtfBFYsa9EMulPdP
kCUmz2CARQY8agGEyV1ZfFxWMRYyv+ke8r6MQded1UJXAVkzo1k/uIFxjFxL
lx0Qt2z/ESHNUVd8fYduSiqbz/joHZRnoSFzSNNzffgGUuENwVEcqjKKq5Hq
l4i3Nd18ftr+eiH5GzTTnL7B/djz1uK8tkRaqo6ceiWuPdxqPIE98ZfqPz6n
A31f4vmTdeSEN1vvLb7QSUQY+tbT64pMhZKSlK7fCbO45ymR/PMSHtHRtlIU
iuakb3iHP9EdzFbm6Z91Xe6gXTz9MUbEWS+zE3I/QzJaW1CM8gXBiPeEwptz
xit0RSKBNeLT97FWkavwduQVmHmn+otq2g2EQCDH4vuf7tHED+Ft2HP40lzS
S6T2JAgmhBGLl4kMI2TYPgzMk/2jeoDTEPxx61JkU6VWdFqM85d5QMpsRprn
30pC9uH3SJRwHK6ezohlIvXx2yJs30LjSrhRgOl2hHyZyeZWZjnfZ0nF7hb2
59KJnqAtVr04U6OexVxNb0bgwGrvBLgxHT+o2xWvtz/XaPxhQT+prk953gSJ
vonQhHYDJufxkbw6JuWIPjjWPUM9XDw+gGRN0BqYsSi/3jW3KB+FTyTC2uiA
CMDcS3dda2AFnSY8ss+0IG+nAtl7YquMT6dCIBcy/7sUH8ROA7lY3MGm6Sic
0as7+U7qhX9yOuwQUliCsGytastNDsk4QFW5M4VmY2Z/Vc61C/a7xzI7fKLD
Tt+i71CSAkPgCNb39N/TuDY0KlDsTv+w0Kw4gSvB8tI4fPDKCcbe0v3dCP+R
8op4KVkDOl+gsierRMlHiLzGfQ2cE8haR3AvW2Qe3DCz2dFARVc5wzoNdkr/
6Ee8EJs4hmNskqdNdYjuDEJB2MQ21Cz7uJN60FAy1Xhs0nrXeQ/kyaFA5X7n
55m/atnvl0VzC7KhhaAbgvQ6N19AToJHNTnJtiC9D2WYFjgGZB4nJvAibL56
CqJC5QFRGyAXEthAA3FGq6LZDMd3KK6b3+iy6ufwa3gVlZfGQMvb7YWaKEfM
QCKQYeEIxMVeBqNwvFPEYAQKixPXsMsCJvIIDGj7+XWFuZjCBcqIPfRMe3Lq
sbxb/GDaAeq562zrmAn5bPxooIZRUa8THFATLcjzPxxP7Rpy60QViLCZEfMD
3sJUVL1qnk14PmEPynyqMghBxoigUaMNen5EKpW1jPt0Rq2oSVQYsTf5vtDt
d4NKhOhHERbp/yYfNeoGtg822G4E01XYZydpaE5kMfZw6/N2MJw3rKHJw1tp
OyZRc1VaVWZaTtvMECN2RzSS/QA/ce4/ExhKHld7hCS39DIGqUM0gugcRWFm
U5o11cQwVlxmKf7GEcdaPwJNspwbYKBSyJy+Hzsz7Htvfi2sXnjSQVJ2B+Ku
VF6xo3p5PGE0SZHX/aeJ4Y+C8Jykklcu8P3oJ3PqMMk+PB5dKU2rzUMspqqP
fn+lRjKkl+mdu1nIvDv4xfk4BELzztq8eYmno99Dqke1+/2TmJkQ5ErkT1Fd
Xr+cN5caXJx25TRHNoc49OiaSDKSmYdtWsnvcnpFKEipIacW7Q0JRollzyKA
nylypMIBX61sSce4xpbwZ45L4OsHkuRMpRzbxm4b6omADdaEYzoPrZZRDq4L
812D4YKRll5g0VIcLn5vznBF1mmvTqwwiz5hD3XbcAVI8Om5Hhu/yV9VxI+e
ra1DD6U4QEF9Ppc1h85dP2OMYUs7yyguW0VPfvWhN5vSW1KfGsL1vVF1kqFi
Iy0ouAJiiW+hAAudZmf8nolv/V9Kv4whuEAMFmfalIMhSGvmLwr18dS8tLoc
gVGPoPLAlk3lj0OHoSep+LHdgmqSgb2HnNtRxqNNzikaibh0NcgsXYHFE0M5
bjgnlzuvplXhQJcAVpvw+KqQDTZrbvVyoNRcVLDD1h6nRJx///lJNABDBmnP
sJLu5TvN9rhKzBn5avWs80fw+20fjHrbKWi2wKBrC792HJAYzIm29ESVJzkd
DG+JbvNU5f3XJZhV5X8ypR9R9eUMFcsdZDGDHDE2GGfx1kcip4ZxXdPPW9Ix
HsaOAlPwzYH5ByLnhmcmGCm+wMeEN40LTvli8rQI34AZg2mTcR96zq5+Zdmb
mfw4CQ9Yx0o7MmmrxmNP+67jVoFpIK2iKY6nPu+fktOWQOQdFedcPr5VnEZ+
dcCldmdzPUY792GgAinSFe3hBW8erq1mIuZmpj2dmFuZJgm0dqWKSNG5pSjR
Y3G9sd51n9RnPj2qPt+FIcgP4ADqs2JDgruCkeDbvrLYJf24RwjoGgDH+bXH
vK8FcgRa7RLT3kfJW6EosaLqtFQqoCsd0phLzHC2Tp+yb8OQkTx2E5qERYYB
Z6F2ACChlHWHejjpALM0vXoNuZhvXJ10xjuSPY+iPjHG+/Sok1T2RDeFY082
a0Nvp65i+4kxbqd64SXzCm3St2Y3mD0kr0nM7o9cxRvKYOnEa8fIjxLGOCkm
0KKD9cuJlZFjhMcljabMOU1ArMK/nnMAm6lV1RiaJ7QnvmpkJAN+3vF+oRFq
BGmbk90E/NvxR5DPMzQnUCD2N2ifOnudWtNgrv+ti/I/yNatBh7PJbrM2vDI
m8I1/1nOHgRSItjTnYCeZFLLwbxWijm+qAnfnoKDwmk+ipf/Sc3NuTSMwTX+
Y3uyAV+xlwpfR7gO9s/Hz42Z/1lPn8PXMbWh8AwJOnAXW8oG2As5d85Du5ZF
0KvOtuvOw/QGhlAZj5bQOCaaEU+VWcmr8xKOBrgW+Eb78tdwJ5/WnOESe75M
GyD92yPG9LWcYXwAhDos3Oem3BzNIlJb9pwBJ6oAMJZzAaeOGRdNviT3+xC4
altNedB8Xw8zPZ8nz9ZQ9fmDIpUZTy6gzBGGr6P1XUw2tR2K6cJft1IndC4n
7WzGVEEUuOzrC0z6NjBn3UHf5pjh7mp9a2JWAM5Y8YZv3RHuFgY7HRkZNAuK
fB2sX32LdDx0DGcoHyOGVDdQAKKWlpILSAKwVVJVCAPjcE5wAHj80EOMy78f
ereUY8B5yEBcBWNy/tN0zcizt5VbNhcK5J9LBqV2S1Wdqmuhm9eb10hTyjTy
hY79YJ0CobLpEkSjlo3mcpKvDpInLh4sHgFZNxxVIv9KfL3Kp+gCeWwIukYO
mGzprPxW95vncN+4tvPa4Gbr6N2mVIOxHeU1YvEWUyUfGukF86uSAIpIKlw7
WVNFOY5LZvgJcn9+ApDGVCmdVezmTA4+Q53090kU/zj6HrYJNpedwiax4nz3
wd/anrSRsdPb/bilhqAvsNc6z+tRyNAeStJou4ZJjZm2MQuxYdfzmO+5GSAA
HH3CPXeqSetkCVjBTMbAcz4wOeIaSNHIlw2NmJf4iYh1QQfkrEa3hJbNOHMe
MhgJ+bgfDt1F4yktkyyCw+Ye7fGb+WKVoY92XMhv4ecSzzXeFM4bP8bHU3hU
/8hG5Hm51qOWyUWrHQ/JZI2vA8P2LdCe2B6pouiXG9GbFrG4584XAYJMV7qP
5I2OoMBouLr2jkuBsZCvkmUGnK5E6hQpv4tw+Ghpgci05SZCBYOK8ofGmx4J
3vQlMq/biyCMqkGWjU7CT7X0IlH5xYGH2kxGsVTe7+4ThMptRwxMQb2g4sVf
v9ABvk8a/a3VFBAITCrgtiPzveOIAAuGUfxJf8Ih0Onai4/f9fiCBiMTA4Jc
+YPAy/qgovCvk5DhzfGyTDFEDdSVGdnHsdYTVCi+m5CfxCHsOmtVhEP03GOk
L3PWb9PCkSGg2IrSDrXeUYS4sBHRWzhoyhsB6Z8StSv5zqi9WmRzlWQqsbxg
1Y7+YtALqiUh0SyYZctFBWT1GXTbZFz1zmnlpnY5jqrNRdG2MwfDEXWT1Aef
/Ots1CFKkUorcgh4nXiKxSe3wD7yDuyG6ZbeGf8X3uzM9JVFd2AIKam6dPCX
lZejor0lx99xXOS2efEHSVnvRZDy/2jmeu4mgKUEU8rmkqGGZXLyfdjTQv5l
0bJ2lHFdpKoltyXLWCtdg3APGdR8m526LB88HLL4zYMQLUro2UzwbWi8ELKi
Ll8f+OGdSxDi3hHTzZdwWvCvcfQvOqll029zl4LloFZT8LAc/utLJUyV2X+O
aqBOxJEvn3qdC7VpNuCMBJFq+MlzzkZat18MqKugJQn2p/WZJRpGvhnMi8DS
ZD4pgmC+voIWwzLlDMxThqFKqnKFufuxDZj9C1qLfBzYGsf3S5Brje1fjxoz
d7F96+Jtqg32jrxIts4nhn1/pU3zX8AG4S0zb6d5Bpr9DdcdTp534Ducd1it
mm2QG1qcSPI8YQdCD1uOgYccUlrPthbJF8KxhVRd+w1IE9k2wv5rsp+KjkA/
LGtaa7TZIoSVBDM7IvUMgVt6T+ssQP+AUKzE3c+T3/9Nu6e6k0kV6VTpQD0V
3qJ2j0SWElgNJIntcebcqK93JUrUhcr8TQKq1ufxjqoDSxLK610YF8LjxKPr
CHbnqOeD94HQ1V1F4AT9JRlSg3B8WksKURTc2M9th5lSsHo47EBHVFPViIQZ
c6HuP/1EfkCqo/wexdXOcOhHSSjZt2ArMyohmb4N3OxMLYeA4aPgr7hUceet
2I7qsGyFjQ3iBTphejch/50i+HhEpkyLggAa1JmmlMMe6Z3ZTkOUqwt+3o4A
Jtei1SxzlgFZGyg3qSajGER4kI/i/kvxuokGdDZc4U9y1jM7qyLZDdIaH5CP
g24KHZQjtP9n0Wvf+HVG4aA3Qb4ANoq1/vpS6H4f6uePDeQBdUCfSk0ovzc+
VVQPleUodQaBlmDTG0cmh2ix1WiYawDoIQeFlsZff43jP/ZN4konvbFLdqZ/
QgSyv9xCpJ9KwSda/YQybXjvk64A5CQt6HRvoiC177xclZ4UQhS4/OfrRy8i
XTUVs/wd4pl8ZHUgLXXyH78ttqk6NYdagSQ/i+SI8DsdDJolsJMljpq470dD
5Hn9LzIB0Fii0SJIHeuoQSxUQHnSiMfFlZ7irTTmFH72Sgjv2seS0fRnejwU
Bk4J6WE06lvkF+xqea8VlGYVUclqRrpKYrK6gx2/6+HuCdx+BB+VdnmnLxMK
GHxdYA2+k91vWrt15wR6d1CEnP4GXYyIekFjvSJeqidLmymXxsE5AgEDuMkW
v2908xV8PqNuZN3m8/oyBrksSeNVJ4oJ1afUcp+Ln2nUeEHe7dJZdGpL39zK
zwWgTT4QMRUnqUX4qseQNzxbsJKhG7amnEcIwQEB9oZselhG6J7Q68z4+8bd
PnaY8NR/DHVg8eXbMe+DYcfvmRxt1IchxGv+5406zovxDNwyJPvPQS6N22p5
XXdtESET+FoFYg/1MK1bu/f7Tco2Mjd99ps/RM7bW0HJSOQxNamyKShnQW7/
ELNA2WdzwqRpBs+7FE99H/S4QgJZ31jY8V6fu0xt/wPnQKribmXI9lvfR+UE
lpTtZwlihonwxUeF9tRur2OGTxb80lvnd8/ZrxOSQRDITdGC7wGqnTq259R9
4Cv1SMtKBj55q+wXT/YBp7G1KPNm+fCDqJEbj9amyVdA7p8dWYi2Pg2q9/vj
VKo8YeDrXA8MfiY05GTb6p91fP/mbDkuiSSp7GJlQH+/wOPNaxjGh5Eo1vRo
iOaHJCPsyRbVKpZhSti5l6OqDLQA82g3PiNaLv5FNvSqQRr5PxlgAzLXnEEL
yHNhdsNbss4rp7ql78BjxmFWdor+As5egT9I9QLN9giq0Sx2sh+Sa/31kSnw
3RB77HDPHULkQWFTG5CgWMKxM2XatgIxu9+16KcrGl1uW1vZmjvQb1/6/HIX
cmSSueYbB2XSNA1k6XIoPf2raDlqhSkhrzJpRBxHKINHWDWyO1vR+iNM5ShG
KkqKiXgBfwiGIao6qdkLzLWn1hYGQizbwEZO3mVjhma3NC8svxXdoj4Ihpf7
ZlDXVNxpg9NkVFgREkgtCzi6f3//diR2KFgFxiP3i0Z2uv4RIUkiY4p6l33A
WqofErjONcux4fvvxeaUVRo88oUksPo0K3uYaIwKo8hW+jcm5bRM+y0lFNE1
1cJPcpqUpJlUykzp78oHoyTQEXqpIxBAGv77D0jpWktRfPoUh5DqNg1idL4l
6TKCc7eQMmfKMt5ukUf2Hqth4/pTt7Zhc0b8njxMtQkAjAP9NeCyTXpT4Mz9
r0p58kVDvqkZbGCNm2eMo6gJ4gexQ0GuhtzB8Ob4hu9oNAYj+NRAXDuAeD0Z
mYoQxNnEplNfBfUQGE7cDqdJ9JnE3VArFpsjyDzmn6lqkdKrVmWYMrUrgw59
97NF4ebffiKrzq2xso4ZlgfBjQMhcskg4Sg2o/6PuuPxxHg6SjtHfvz94v/l
kwTYjp9T8qzunFUvuv+0c8gmxv4PXnVkubKNYElan+Ctb8PMWdIK/5qQvJmM
CpkDnYv65LLKcnHX7e+S8DsguKSsAX8odzJ8cmr5DSZ3Q/OQ3a54y9PC7MAx
3kqnmNe/F+FcMAIcAMOrsArtXEX2Yb8xELphIN/YALpUcBDgJiuZWMsuhfIx
joNGFcmKKiWUZ6uT2OdREOkc7YbELAcmGinsQSRWlB/emL/NuaVTaYOFGcHm
sxRynJD7s7rhWdE61TJwWOrPTXFs/6f6r1SXdpRwnBWoOkD26wTiwCiNRcnM
DKKxAOpPxsWMTsTjRwTM1YUKCegLo7J8VW5dvtrNn2F5LJ3EStTqcKhw1EV5
rXdLvI2hgSixbma4XoySR7hzq36vFlXaWiv7bmym5LxAoW3F/4RESE4diob8
cy0lP1s5Cg8+xQVZhQ3t3QgrJLUsDJnfyJiEHR3mAKfq/UCdwwMMHZlZNnJ3
DIQTXtncJPqDX/eFRcdYgHQ/LokdR97PqaIHSqpk/GHGBFkpCvZlI58nIfC5
qd3YZBAXzH7INfvf2e/h1HlSK63teX8BQ1jEU2NlOeFwOVvkIoq68DDZIXP8
qYELoAjlT8w55I0g+NgJCDg+8l5x4cyqEHUwGqcgCEfJzINHfDKkzPhAN0kW
6g8fcZMPx7Aq0Q/7mtXz9/Yg4M8hzY1E8kXlY08jbJnuTMeiilzb0/YvPaRC
dwxJCKi5wZ3PkzhTFydsmlQhRTY56a2h5GOnu5fGe9vhDhD29KDtcel1HmYs
95mh85m3Cn6eTCtWMK4FwUn1FCYFV+7ZOSCh4I6WsyO/PONJaFd2MRD0HOs4
svsDnoTIfor5fTgm2mClMFcgtSWnUGXkO7ao+tQ9m6ZQu7AH/4pbMnzhAHWe
tHJnCGa65qbsWkBsYil86m3xL4ev2SqmtruqCH4DIFAgWSKy75vlg08XEYjc
NIrR5l/w0zbWP0WQSGEU8HZ2wJaRfORWdDg5GyewuHbghApfR/degrPXEchJ
bBL2vwkHFf5ZCn4EeHz7clz57FHHzJHmdS3DL3RYLjzS25hJaIYRKBzDe9Gc
W72ikCV8yWM1KEKSr/uEAM6h0TUKiRV9NhCB+MbUVbBFUFFwbRwZwrhiTFuZ
gE88lBJKe+5Me0p8cZ54f6hNwkAV+VRQzuOIpj2CY12J3EKeZAFVe+zLKy8B
+56dow9AqUTYjBTyHV8LZKEqRvBad5gcctNcXBM+Ygh3jd7nH7fGcjUuIGKi
BFje4eHbHpLXOShnKfDbqutsNz2WMOBs9sgszdXrASWxOOUs8m1V04cYiD+m
/M7MyBZb4tW0Yl6hAbsSQiWqb/E9IYXw1pNRddBNDnFW6zQr9LI34fLEwjrh
0XnmSM5/Aw+9Xx/AXOEE+GeDw46+4mnysQOfW9aj+/uHJUKmEWLTtMi+rMxj
z0FM7f8JpRgmMkKFm9XxNe0WJ8FqonSNx2OAdLGL66IfKZ7NdKSyxdDjt9jK
mXZwzGbMEess3n2XB/EGgUroIA72HI6aIYPKmsfPwGsU8NKbchivrlS9I3Yq
FF/Y1f6xBies+rzOZANxxkAl8eZquxWiENtbBaR6HD4sKAxEfzKZfnnU2SHT
A2hr6FwlV+9VqsrBxdO6Dch3MBF705guIYY266ghIvk2iyQigFMV8UFqqTdi
jwA6GGu0DSixwXYuixFlnW/78LDQoKvc4p8a3e/3xIhTasB9yM0YJoprQzwt
22PPQMIWgbGF4QCacSpIPeojVDOOxYki1Ixmo5WTOBy3J7NilXoUr6nHsW3e
eDxigiZZW7Ats5bI7zgDiczlqgU0GtmLLc71eeihUpcQsp3emkoEpND91Nm0
RigYbGKB71O1SONZE17+11wWsIBPQMG753kbi81bxSEH9uQ6TAtr98mGAAV4
isynheX57ctBctZFw22i9p6cNT4443fVB+iZfkEaTGOpBljcE/M7qMejeTBG
WPEJpoWta1EdeUYUzh1fMBvgTJl4Ag5WKjWZ197V13R0cp/mHe5qvry1uwl8
dp+WMyXtjkLWTiVKHB1wX4HVrjVvjn4xhy6PxPqEzKnf24DLAf0XLHyQHD5S
40oH7k31xrFuQIFt9eEWuAbPda4GUULvCDB1VNcM78Du4Db91wMY+KUt/xC+
oxGHDTAKOUnnVpzNvWcaB+pO8M7OUqbtzdE2yF1yfSKHibe/2eDCcNotMxbt
bSLCvlqd+lUmnY+D0ZMzE97O/Ytyf8QmCmZN06UTk61SWzBJG+oVkXVG0nia
JasCof/DjWDyXe7tO1u7yk8xHtc3s/o3yXn/yk0aKYJrggJ8WMJ8Gp7dbVS/
BNFKVceGG7RoDC9dFRO5HTHvPhE4qrRGiDSIln7Xb5z1f29O/sO5etvFayLo
SQgLmyuEJt1OiXsFv5MkYNmFl3xk0Q5Yp4ndCQXdCJytTHgWn2wMxeVZHN0r
Ww5o78wpzkSbDMtXgNES1AZ53paKsCWWJ2GrViNfQ6tqWAI0qPcENYGe27sw
dn6X2Ykdq7SOqInxTPwjkwnqz4Qygbn8++gm/UWYTVqSWx25w2JceGk4Tup6
IEZTWlqIZentG6Dc8ePp8vOdUPZHECV9bNgNSZ5d4yATcgKs2aBoGZFJRD7E
Nd1qBkBde5sGUfYxve8EA9hYTnPSRpggrg2BKqC3aMMUk21ykhkbnr0SnE+A
5n5kXaQhRr65TUj5XRB25pW71SXQlu/5T6FlUk9uH2eoF0twrGMp3psGoGFV
D+opJMG9ed7LNzQDl6YYqC4IikA1Gr10dofmDewOJcvGyb+XzzRsMC6ltnIt
ysdLPMdfNU9BXVDOpMEYmzY6FDnFm7CttIkkH+3A5fBRFBGx/UIZ6rXYak16
jq61NueaRBJ8R9FQ9ITaOUzhe8rvvXOhQ+9xG7rfdMhtqB7xL6hLV8IN+T7w
7cAmLIHhmPsUazpQ/yWHw1VccAf5DdJMfNu1cGSK3oxwFXBrcf85HstNqHWV
LpgCfiwcWjfrOQYX/8mvwsO5yQFtMC5Ha5tfU2hRjrzekNvY8BJnajEqhqnK
ZBi6TNpKbzM0ezTQ7dlDdjE9rlu4iyHUxXKoHIPSFg/uI9cN/lgIfS44Jon8
2f+u/AeZVn+Wz/LCReOJbGiDSHwc84JxYsXjIoEPLunySg7nMPXofhaMQGsV
jY6wSRqbpW1hhF6Egb4HVTW4+mj3HXd38oKiAez+IZhxz+uNpZqdpfBCHHdB
ArOoBxqWqMLg6zgo781wRMQvXVO0YVXkdqd1shivByd+ghpER2qP94vMsrWk
NbWecN52C5eNXp9rSwauhaVO08Xep1BCCz6dN1meYV5uyaHV1FYWdlo0sVsM
nrkO2w27qL56x2A/uxBnU12QuUytODlOk8duOLHslDuTQcWVLh0d/hP4WWgX
J1LbtOC88ItPSFhb3lgwSn/c7MF61V2MqQ8wjhMS+8VXvRPvw7XJbKnfBncm
DgRZKTH2yG0MTIpouQU1COZ06P29GBkSTG+gYaipiuv2A4Kt82a2xahincqx
+ful2C7wIsnFEAF37l8bVQF16zZYaBYOxOzLieDbWh+4PEj8yLxe7yAiD5SD
SXDg/XOuYDd+VMSOXjfgrzz6HcRcDC3esVHZqCfNDlEgaOTKBfFpiQeptMxk
4YliK7IJ1si9bBydtFdn5cf+bqTral3TSfoLXnXo+o98/SJPqaV/rHni2meC
4oEc4LmKZ5+AknwTVFTvMleeG8iYRRHm7KwpKoVQAmaVvjBbEcYoEMwZHHq7
Cy3H9Smgulbr22GDJGs7KiIfzt/v/hdS5UnTkDVc0j1JCp5hoP5Kg+soXrC7
E4wh2elD9GBorTrXZWuFMiEkAt+1T7vGvH8byE/3/naSIoptqqM4IGwq9PCI
simzggnW0BDrCpr1hdOsybyyUbb1F/uiPefu7ysrSNtkDKdOcbQZ/a8yjjz/
8Gd8+63jOM8vAcgdnzzLWj0B7T31W59jpWCGarnGK+XOEA06c3LuD+rZx/SV
VJLmbFTtxe4+l0fYTtcE8BVmr9f6uDCqEMqHLXGdNjFvO2hPRf9nkIREP4SV
bMPSre/+nVkDBX5Vp1X0VjkQkxELuoGQDax82Bc4Gp9sa++KJZ57+q3X7DxS
9MkawPA6N6C89+erN3PDcyBusvK/K/duFLjzlc8QLE+qDTr8gujJZ3Dqe1pm
QQseM/wdrLsVpV3iWzMiz3mzJl8o6XhjfUhCkIvrTPTEiZZDZNGYf8toXXNt
JhXTU1mQVriL/pId3RARvUYfhweMMgEKa3rElDglpDMQmwunfSU4zAVq0Jlz
3rYKo3CGKP4BH/3/GIz/nPlRUwAyBKKa/jGGNOucIyayvej3waL+v3lmyPtJ
bpcuTSvOfqFpplVOjeJZZpicf5+kLKfxCDf+oJWz6FHIJn9LUQLLonJykCjg
LuLxgraB0mvxL3QEr6tOBAjTq4pgF9cnJZyPBjYMho4XWL732N1LJjmlRIAk
1Z6sHXcRwFofv0AZa5BJhTt6EVE91rMhoi6BJ99af70N6oyc4ALHYxcJGpxZ
TL2iayPDP17l9xDlV4epE6G19mtEnGuEmcuysFkA2VRo/SmHIgzJuC8pJmkd
bwp6Pummm69vf5D+JvGqXM1LIWHEwk+BC4FNNNNv8S+146yegc8B09DHmO+E
DJYSVXFwwwrkhysTwW8yDNzCdoc0125wZrEf8zymnpNb+lT3RA7vqZGPP2er
ieH8PRMFyBELg/QyuZtuRIfQh5K0fkY2Qln3Bq3NEZ+hXYM4E+VpPOnGMIzX
0aU4sZDyRAksU49pYTkKD+OmBNArJexlLcY40UvdlUjHGwgvYm5wPICjlSTX
iORTDXatBAcKLkv1DOEnuI2Rke01V0CoRzTMUnTJRNZz3MzHujb1hyDyod51
vMSMWwymPr/27Sal35tcWhX7qsFe1cYnP4ZT5wFj7hWUTLQoX+cCvXBB06mi
+/dg14G5BgL0RrRPBt45hr3rf2NAjpuIH6tocwoFqNl5/gJKQ1BMa3f1Urx2
x90ccLJ7bdwf9u7WTYpJSdTFmdlSalOSJQDx4gB1Q2Le/szQq9aClMpuvjar
tPsNhbcEOXLBfpjxI73ouf1h6Hc72FTEhZvMvBltI+oJAg+Iu+Rz1XQHO7uN
/fipaQ1lNbs1GGrrKE3/jTBZ9vDzJdejMTM5A3PU01U1R/fCB531eIXhPc0g
7xCfTecmmGuM0AUgq0qhCtz8qWSB6halV856U7r5o7ik8h+nG0Da89MoX7BH
7OUVIPu700wyRMoPal3lCpX/3g/PvAcH4lgUoH7zcS6Q2OtAYZ4AtiWX+fm6
lZ+jZtBdNveNPJZQ35LdGf4v8uARG6EzGtCgtULXe8SlTp/ezZrXSZF72j7t
B509/d2qqjlGrqjMxOkVL5IqWYsEYlrVnsh5SQEWbtRaNBYJB+eafXiVNEKU
u5rjcQKPbO/FyVEPdSToGVDjlgrs/9k9nIPoc37NDtY7eCFqfc1+JKZtz6Lw
wwflATUYgCbWvr5k3RKr1a1ksthjTMeIGHEGe1miYruTft7gDmssGFUg40oc
92+lykxFwBLikW02KGGcAh4YKWBcQQ8tHG9MJqIIEPcDDJyCUyilM29pvlvV
3uRx+2f7LkRvJN0m3LcBPxttzHYHhz4YGASnh1k1OndyLH5S6ey5UhRzA3SH
WraqcDeJuMuMD/gLcsfis04vb1TU0ogl4GZcocGbS0Tr9gq9YPA/ZHZGppp2
9rertLWrJ/sJ6AdzgGWOz29aubeI12ymTnSfT8rk6OCEjzxUafFt6rJt82FN
UQjP5Om5zq2pFKaTA7qoOwFdM19yRrY08BiFiLJLgRylCZ3yY07mFoluGKlT
Uz59PpldX5m2R6PIV86vsnWtUmEbPg7x/ZlsrB3/xj/bt+3aJ19UPmGIL6Y3
xeep4ecLrTQMEjSPAvCTCORkMhiPk8Zy0zAWSVC8yIMkRtqXcUxqEJB4+5fj
xw3NDhbWSOjQIMqPzdlAAtnGt69ZgJhft+2LAIyruxPsv1CkhNBOIz6VyXTq
Lsm0AaVwfxKmprPORQhyXMXAm1sQdi5lKVM/siAtE8+dN2B/KTJDFdQVs018
Vq89KXAK9RstOw9rYp6X7pmuUsG+sZTY02ubCo/PWI7DxZGghYIm0HaMmOUQ
aZcbhHcAr1VBF941FY2U1KAUo5m5Fky8q5Nt8B4Jz+qkknjM/soks/NZWE6/
eMt9Jrl298RBGiBAqpvKhcZVA7x232MHRlNvkh089vg+EMDxmU4gW1sQr6QW
uECTEGWLJ/ar/NKNPKu0mhOydbmLTLCK0j4yE/5eJ67UYwokCV2tnlDfxKer
LQyGP6ZnwzB+oRQKhCxtd0jE1gbGsp7KRR0KLWEsGsDuzedh7nS1FxP0L5Ln
pJ2laHG1lbSTevBYHbNHasjgl7gbQfXaiolhVKYKLARj6z4UEQ30XtJvi7x6
mZOS1Gbeca/rqt7XpNhUBD/0yLvOrCSU123TcCbpnjegeRfeh5Dw8swtc0lX
WBXBP5q6Hq6ZDGbJbrVzGPktheVn0+8JGoSheoYzxUB6Dz4Jh/SDCYENMHU1
tibEYbCntT360awTrYE6SI/GT/1kIuB2NRFiw0BFelIKsVPtmNxDNU3KPdnE
dPYQHNhP79vQF0CNytr+CRFOg1aiTL4jKYnvViymOELs+e3ccZKIjfh/ujZv
0LTgvC8f20asrbuG2ARliZg5y5hubd5dbmuOLn4ruPV895JeVFjDA04m0bDG
efdGybn70X/f33WxnXVQpuTlfriL60beyFXjgc2PzCstjan4SPCQq9XgYlR4
qH89jXroNWWtUi+b+uE5aAWY5Wx/wvenvSijy8WYrR54dvXMd+U7x7/fOotg
+VY2qciaR4JH2MbGYvNza4vDOXvSEbXOOolx2GPvXF/WlGfz8n9Cou7ZK//Q
IxvPMYS86+eAQR4n+ws9Q9M4F8wNa3ftXyChgD+oLXo3vI/g7ASU45FKJZib
KpbuVKyedE38C9oWigwXHCCnCMbWtMT7pr0w66BHfzmuStWlbbO/QegdNY5s
OOGBISEvvn97riB25HRk95TaEZhbukTvJoFJYhO0N2oKOIWcV2UxraOQjbbt
eH4OKyHxifgD8v5P2AHnsrw8tXZ8A0pxBwRRCSRpAGv9nFJzIJHt8Tqd99L2
ZOL7CGEpXGIMCaYDi5ss1avBVEyHNEJ5+ki0qUdOwGZqxR/nRIm71wJ+w8il
pTNt04S1w43cN8+QH+Qz506072Iwua3FzE7w1LTXWLI4q5jmM99edRlyOl+x
noDZvhb87PKpfGgiEGnHEOrS5a0I8OdiHyHQQDg4BuwJPF5SifDM35TvmSVk
/D/6S4WAj9HcN6C12JwyqinXDcUGRbpk2NBiQQ+k58lsbxxFegs/SwaR4xvC
seakNbz7DEJAQQHDfqTDndgRyvJh54yImDQ7m6Mlq2k6MnqdjnEGfq1k+H94
nCl6l2GZh+WoVHTvCbPxWzHxIlfP/8Crdgbao3zC4cvBMTrPF3xjDQ66EBKN
Vmw/fgAOH1NCY1ZJBXklI99+4YbqiB6R0+r/xOk1aOBs6D7YSlDgtmTChWOW
tO8BfKZCpjLKAIOHQ2mp6lFwhsWRm5SqZrKeELuqwighLmcuQXfybOv45QV2
/FTkCXJcoAiAnqVhZR8ujdk/IzHC1wArBvMud7GYkr9zmjPLy3QL8GWRLWqL
z3BEyh4WVtFmhLggWCYTwRXdk1daNrcKvlv2zngxCqaj1P4EOLsCW2hQKzWi
7tpgpACUW3eOU3jExqQNhUO7GSyUoiIXOE1s8qGMSgTSQJXDx2bk61m8ej4x
XktMU+zOOevzHxo4yxi2DqSzBPrIRDl+P3WTKwkhGw1kaaPqfJKHxyKj7LR4
cX4kxrnbIveRxiF+71v10Yp8AfEVdArrEf0mMCUDsDfp6d5xIuO0oJ9qDyaR
Y7jSnV6EbmI6rKoSRhFmewxIbGERJ6PXAXGE02bDSzizHIcfzrGBF8Eu8bz4
NmNXxHeB9sCzng5Oh8AhA+W7AFZh/pawF+12AYBIJqFEq3jNbfz/jC/yweEI
ByyzXxG6PRQ50AfRHpecnjkjkonzqX6f5tOR2iIiAjQMmopxZi2m2iC9wbZ3
PFOOxiLpy01eu4tLah/jdPt1celoRZvWwfdBzOxy9A+LI4HdGqq6EhUHyTHJ
icJpzSJwuKGJtbmv+Oic3wyVE4zms04kYTUcwjxkol/hQWaUNgjjdwR3Um5b
gjt/etbSiBjAktGH+gQ7pLjT3DfQlp02L5aYGvhSRi8Ejyo4TX9F9dEhY/n2
oNKNNQw9hkcMNI5Nnt6q7bUGkEn+RKbgxEjNRLFsV9WNDaLf+jXMSyBBJqIN
ppC+Z5t5eX3+QaamdmgHOIeeaQG0nIwY1WLVoNsut8KMK5WmTgBuOOcZzGXk
1+y0qchLni6/JfV57+NhqgqjmNFbYjQJtZJr8AyZbUiyHHOSSsTDaXB64cP3
X1A2PfrmkTuKw3xOXb4cgKAE4sZvCk4FixHMlP7+a4UBARjbz8yoBAjskr0u
1xWiThUPHnm2nQe69E505WoqPvBVIS9L2ZJQH/mZSBuigQgI9Yfbbi5MUIEh
fTstGa5DkOwIcyMA379bintx2uZdkEICXJG0zghecL1XQjwXzG9Amjga52DS
CpC4Th5n7pvhG5kSAD4X63y2FqY/5YYcmnIFyRwMFtJoiz9GhQOvA9+NCp7R
nxyhbUDfkE60qOAt2UcDmR5+bdV3g+bGF0KeEVcBB/fqHox9gHCiSwUSs5hp
6kX2SC2fiWz6zYWuStWniKq08C0+wDUG0lQciqIXpP1F4MUQhuc0gXZ2yeYX
k7ARJxiJsY+QlM6EtUOOgSleiTsy+T28bty8qpTlQrNKbSseKCeWPc9+Uxp7
mz3o1FEAhN68wf9bDC8Ejt/NjyCUFALmiWTr4Jx4eAxwwsmCBsu2ca16Bwtj
miRR50l4BRRxGhdt7Y2y1/oe75nTcHshqz+qBqHJOy5D43jAPJVsJObr75ge
OLi4uquOpOxEx2m3XvZ4W25oa2EZ8QkNbL/fSqs86tjrD2rCD0DlyCfTaIS7
AZCD2zAp8+3lhPDICCXJ6nztElrm/QwtUvnhBdTNFIO38Ax1MLkHrTE/osTU
UYyFs7LWIlAqmw5Kvq0QtN9zOuc2aFywsElM2sg4tm65RE3HHO04xFsT0icK
ux+xu4i4ajXIiMxPvKRzsyGvQ62cGeXjvi0RmeBSa1qYNitAVzHPzOWIRy6q
FN75HNAWbFi3w4U2nOhTZ9rj40tAYsD3M4WUnnS+n1c5kYPsAJtSOkvhUCu8
naiOFucuD5CdCkVb55eEPg0RqPxRuVEaIiK7cPh+ijuf8WtByxcINVgTZkbO
TaTucdN2kJKtRQim6qcc7J/lRywgZ2u/49icjjfCkViuFPhExvYHIaKlQzM8
cScEnCE7zZ3x2/FL4cxeMfwUAOZtjhKNYSn5e4UMGD9JXUbhgiHHc6H5COJM
/ZBeqvpfEGRsWaeJjJdukesy0nqIkWOk2NvDiWiVtOpxmAg1xQOMbRK4dSmx
0qNycO/bpHX7Ty3EP6kOLm1kV2x+API8GTiR2JVtNVGbiroGXJi325sXRtcm
5YilH097OCBlpvmnFkb6a3Bo+Fu6ZDsrEyTdDP71H9kAuDxNXqZ/6utZ2iXQ
JnGubyFM1aUwSqYCHENZYzYo0YO1H/ZJ4uDifMMrjyGSmGRcqENqxrwc1UZX
hWrcDRrpy7rybyeUQN1OGfy9Ea+GVgxsK+9plKm1VnM2Ex9MslWHymh3DJEz
HQGWHWFnTfYEdxULqIE3E4yMqhdFq2eHavNnQUSzj7eV6QoxntqjTBOr0gyF
d4tQZYLPOr3hEdrjBibAOeo6MsuEbFgWela1eisrxvb+ihsnVuFPrjfKTh31
o+r+/go9JgKyYjBV/3W/fp4eTZ/OK3odqd64WdKCkMpRPvkUafFDN0RHGXmJ
THYhak3J8yLHP1K+Eg8cJIZr/oAmsLg6CFdHt3njSF+672mKyBajKxiVjx2q
RlttecaxscAaa2wRT0NRNcFqsfz6qoHngPUURIV4HSSkW36dVRW8tLutMxbH
KnkkRGLHdgXM7whVTvvO31dobYSPq+mtGNB18Unp1k9U3pru5roG2nuH3W+t
HFNER6RgqzByJIOHML2wFSRBXLI8riZjR//0v7O4xkZuUIPtfDtox+EY737w
S4WjWVPu9VEY/lfqtc0iXRtbD14ep96a9sPNZCI3T73uodlMkjL2lnCvs9KQ
vZUhybftvBzd7HS9WQpoYsWaGa3fUwMwU1i3IjZx5heZ0WYm6qFARUJuYxXN
IGW1IHaw75OishspkPVbBZkAs7kOCQXtu9AmiKNzjxzBL44NOX9jb5O3Qiwp
1UtMad/01wZoRSKnOxLsiZNWzeIjN2u7gof5QgvNYSsLZERF04J+y1Rqujxs
i3fd0mREbwkpVyOFc9l5UeygKoDmoJOBnnHCQYf3gP/UbdmWz4qnTFQMoSXv
uWQCiZVXpfAdh0zrPBwAYd11XUh86EuWEpmhs2h9BnyYCtq8DxnYkWsR21gi
WNB/usFrtEBHPt2ibHICfHMCqR7uYWoQYM/xxZ2VMDCgIJnmVelnLU7t7iUM
8ulqvFnbt+4DRvSguPAHvKZYwcydy6ADKj3afVzH0lkOZb1cd9Hb8/AT59Zt
uzjj49rbyPDuCVgfD98HplBZ8NBU4Z594udydbps1T0FD2pX6eLadOaxCXPs
W7rQJHHF37Op12NbsqnSPVYIU/f6AypjcHQT9b808uIhpegi3X3RcwzB/h73
4XR0B1je3Jd9ivRelcmrsbhVYpOFIO1bBT+3gJz5AI4iWDjvKanlDKeFa95P
uF7ZqNKFCtz1017yQNYRkpRZTyVXC4tSnCEJv7bafgk8fjHxTKTk2k5E/IFH
L/WBhJOZereHnign1f6KQIJ/WH+eqcXMm6br4FxL5FU3BnojBpNurELx8EhW
QZ6d9dGFZ0uf5iNouq0PPM3lxGwRB2E5d8bAzn62UPNmTkwfd7v/SiUlKEyH
sqGs6BvP91unehpOvk9j5as8YX2GLtR2M1Iv+tLLVWalpmvOAMmw7PJ0Ui9v
MnlRRW+WAsjYC9BXlsarz4m+6wJb/MQWhkRaBhnuyfrdz+eWY7jsG+IVHR9L
7VI1jCtFo3YX4YQUv3jYlvgiTGmB+sbBKEMmzvGm5bH+5R9SukrCv3fq54ee
ol2EKjfC7AJcuSh6X5fZT4cNwyJZUeNgJPrTVzwXZprVZL9Cuh0fEymU6qT3
Hn3qZOok/kspAwThlC5Eym2o9wxZsnhqExynbH4VC6SUKotS8xWNvN/lCwzY
hs9WeSXYULBqwncRMNBBYAo9noMvZFv2so4fwFfPFob3nkmd4uyYQyv16SUV
WmdnPzvecUlC4xjwqh8t2g+lDA2Zx32f2KBij5QPyEVuBZP/q4QYtCdB5fhR
9JSbzLxhRW2yxP8hN97ifmnzpxgRbomA66aieoUasIY/tFL8wfCuzazbh5Fw
p67aqL1aAswEH/sWYS2WN3/7MYjP7gRCFgc/2cEcXWBYGn9vSOoRofWXHUEx
bzpzjTcDb4auGB5o68VqCskcTcnYwUFytcvIQraiQqnTgcbexwycuQifhMKZ
XDQUtDyKSHqRbCx5il3krSEwxGiZ1c8QP5B1tz0egES6aiKBPOk80rUHsqaZ
cm6Ahlk06oF9Ip/OZwvqk/bGGFc2fj518yjTWlzUqC09LuuTqsAFcFINZ0nt
jWc9IurDSPSYP650ytu4Duwz8d5unUnkAFcTCpx4bYWekGhuaVRN80+E2oh5
PyCw4Q6zmTQrDVzFYDzP9kdOdXHqD/SzDU4xCf+DfJd1fP6gQ/cKjP/bup9S
42/zr68PfCBichTHMQ6n2scWYQ7Y8sOGXcUK9pPZo7R+aQCd/4AcNTNaFqeC
A4/TUfbRLy3yxqceZ8ml+nfiQO0UuY8gDz+DmqNsFf/ZWY+1UwPlJp1mluv7
KGLkFrdQLK7UOqgwXMIB8cYMKmNba5SsNNMNBle7C+W9j2rxYBQfAmjHckpO
AGASHUKH3IOTP0Ko3HuICLdNYtyMNB3wp0VBQ4G0+xkcVvgZ1q/kAYv1uxBq
qeuITCMdyVNo+pHK8RyGlQTS0fGEyMj6lkl+T5j5/6bqB5PbEesS+s0CTKER
emQ7XdOWRu5iHHZkpqav+MWlLJ+1fbd1hSOfXDWst3m0h9X5fAvhPn2nOtBg
3J/f5/oCkkCgFvnyBXsPWlmzStZHj4lOl/N+uYXeDkbzJt5fqh7iMTCojqF5
djiZJlxhqez/vGgKQphWHq+2lDATsNfvLoAsTgOINTlOyMmhp/L7skZg9MSM
PlL0vVCOJ0ZwL2PN9q6SHIbClXJDv2tYK+jxyzsQx0gvhJ18jQY4tTE9s0dC
gqzu+O3yYVimykrxIpBExCz570Vt4jXYEXuLjfD/PH1Ip6h0yjdsRbIeChBU
r5agDAZrNvwe1b6JkEkB2Q3ySzyPdzp/bVClTed80tc9qsMniEJP4c4m77uA
T8YSYgXopy4fK/jeuPJESymWJmrAVy/c9yIvShwFg0YYiTJPjSIGfF6XpVzz
1HRsUxRk7UaB3hdb/mvBP1GzvqX/T4m00Q3c1gKhejUZxhAYHU1zReb5dz4H
dBVv2wHidGvWO5CoM4jpvbOgCre1yDBWH2CdgfQ/hbgV2M+h1xjK2YhUXr06
UZTHEZokx3z/JaikoZpd8naBMhbvGvp7Z5056T9xswxzvKDXZsCCsUt1NbNI
3PEf8QYZG6iHquewpR4PuMgeFw6uJpyNe44miFxSP3hOrMcMY+YBt9RwmRrA
U0WBYxgpndXs0TP+wo3YJ+/Ho9lk6pphju52VMcxh/CFx2UuilIrOMihkh94
dBUNsHpaag3UMjslv4JiM1CaFqH5BMY8omKiw1txPL108pk1l3Hvor/hQcIB
tM2gsWINEvlK8TpNV4s4BGxwqaJ8Idbdk4A6T0L26waqJMpkKesj8vMP8myj
R74jqGQTuq1BIi2ALitKqqY8OVf73iQ1eMQPr6PJ20c5oOiuLtSkami0mdFj
z/Tei00uyOiQy6Bbu9x/KzvyubO22LEYKt9WH9u9+PeW/AFqWnrH31nhCkQ7
TWJmfVPimFr1PfDA/ww5BH3GED3ncyL99vETxpD4N5KvjQeNFY8WMT1RZHn9
SSNkvk1bmOngb4ZRSbVoE8Y+w9fe0SwiZOdSwwUR2vYCQ1Rz9PTbr2KuYjSg
j8tCjGS25+fdFEj4/ix49rAzL5aYXYtfJU4caLV5ZRT8yDF/44CMu20r5d5B
44z0BbAzqIUzSrP4ex7xnrQD6NxXwB2mpJnwOuvZVhfkwaxzy62C27UHzy+n
hT8g64PPx1bBteReuP1i4qp6a+u+hKV1KABfITIGIxAReCp6rJYTrm6QYiBt
TurnzUKt9nBbVKX6lmkbDgEAb+tQjPeHGLeQrKpyatUKJJz3WUAStSQeryl2
q61m4T9g5QxRUu7w736VixpS3KAMwue0gaKb4t7TKYpMEc5bcUvKnoNvMq9c
Vnvwqi43lbKSn2xduLdAuowPI6PaDhJlTd1HAJzOGnPV76/Hv9c2qL6bzCxi
jF4Hfldpjoj9XTkkmYkY3D2ljE5qM/6Njs1GwjyTvfEkP+OnbdZQpQJaECOo
LLx7RUhEpyX5eBLmcdZnb3u1LFMm1ZdaeZvxhlFvNIejiFQUcIiEJRcXbkCt
qS6u5VySfV48Ds8jxtREoP8a27/UK9/dCDFDZuV2vZu09irY1mqI1FEVroVs
TBbs2sR4rU9VGAY/wKZXsnMRO8qlC0oxkq/HRvLx1m9/mFBf1KcKXFtuaAqO
IFtz36C3Zncnl3Rb/zTmO1uf0Bc9QF1dszFqZVSaBmqrnLGfm0zzHYlyxPCK
QEiJR6sLWV9u+WtNANT3xDj76PKGKXGMesTi/K6qM3JfbGc/l2sPNPgexfrs
L55kDVDpfDw4lou/Y3aTFg1JInUt/hKnXmXeGpmLlHEyInS8Ig3vm3kpy/0w
TO3kiFjGS2+n+Cqp6QKmr9OwwR752DOFCJI5NVkhbGPr6WeIjLM/4AI2nCoo
esdgmRzQSOlNNGI7EsYH5t/z3uNz6Wuya7hOLVwfXjnKu3VLRVh7t0RjKjIr
ul8eupprbsz1/feDjQT2qUJSek7UT56qTIJSDSntoDW8Eszv6gWAe5LQY8eN
GPfAolXEFu/wcIqrfqbhOqzvpDU1+7x/VO+GH/2tBzehJI5iUV38XQHpE2Yt
GMbmmlslsyOjilMuB76i1jTlf8zywU93n+i4ixR/XhGt4HrFEj0DXuKkRaWZ
yseQoZFra8atbNV/AII8xSvhk/8P78aPN/HV/wKRVmQxIUdSn8+xU0ttqbcx
uCIRLCjHY5D3I+1GKVoBKRBevToooyvqwSGEQr+t/+tvVOSXyq3V9pv6A5vq
HwI3j3WG39jwRiDQuXZmWDUOXOtSnHJVFNoh1H1WLzzNmYNnzJjMLhSxAAPC
l34g7Fxu2eHPjhR6FEynfzCypsSoJ57kkji7tqwfl9PdRYxP41w25NzQ1gvr
1LmcQkjwlPf3FZA/6vnyz2Kv+63cvxOF30stJVVzwvp0t206yIoPaY4HDIak
YKM7kqtxcw6QfILwMKwSwOK96iXUP56levKBKpLkvLVgQfkhX8hG6bLOc7Uf
fa3xX5oz7C/yjRJzsFV8cDVbvZ6jwhnkbYO8ruHbtGIkAzwCIxRO8x2m8fGc
f0Y5BRxO9aRRMHkchmzR15mJdoibOlVVHCLXgXqs8Kh5oUwWmRuz625M3MJm
DlE+p1AvAPjZzdCGnXE7juA5F8vft8EtRxbVzE/zQpzESWzGmZOZjoK+2JG3
EW8AUKS+IeANANL9mZREF2UJT4A4IVrsuEp4ZPXLEC7MYAPLr1MQFqOfJuEV
aco2ZWiqkFtob5hzS8mGacnYjak9w8LX72TYLF+jiHCyppg6G1COWKvMU5b4
g5RsO4VZ1RQ2Y58KhO93VexV7WvbG3kvJqYjHse2yDyrJnb1mLlUQ3fkbICs
e8SSjjzbj/M+WzqtC+mdpzDUUZgjs5CxrUVe/0wIzVhSoy0389yqrWb6bc3s
0g2NXe/wkk1M1ylFuU4ZXHbx7Y4kJdDkYf2pFdmaonc96+yeg6o8zqwVMDSF
j+q/XyjbhNRZkkbAfI40hnPdSkwXzWCpZiW7rDkaXrwT4UBVZxN9d2S7bkzi
Yd+uT3zeZA++lxv6lCnvGir6BpHETSe0dbOsZedrdp0iMVdc/v4NXQ0pXTuA
ENsJNinoPFjZot3yjgDoy/HgbUKyxMZv3MO4vjj7M/eg6G+0HHjq39QwMPAj
y3RH7F+Jj2CrWAQKhBxvp1NU6AIvAX468jLs4T3kO3KE/EQsJiienZ/MAKzx
yyG/mkzKmwFzwXt/+jYtOzY9OFl9u9jxvJEKIgBSYK0DAOvsHi3JyNAyUJbv
0umE9WX4klyJiK06ZP2Be556YzTivWDwHsJkBNeC2s4yk7VsVFMwgAOrW4dT
tIWoYgg3sFt16BYEfAiUhx728+54XevCfsqtx8nr5tcnplH9ndoHohlbRKCu
sgaGguyPy+apegpnGSi4HJ/Qet5Vx3buqtwwhRMiP4gnkDRop+Vc7ms8j/b0
YvobhN0I0lpIt72C5ZYmlqUpTkd5RuikSecswcJXwOk6QQusHWr0jcMviQVk
ONm2nvYOSKRNdxb9eaE/n1obU6gmhCeV25lTWkza/yzQalw751iko8AyIZye
dqukbjCuQmxfsj4iymbPaYV3tVGarZ01F3uhcEevlzhspik9YowMXjWfS7AA
8hjkyucK6nY3j30opoCG/Yl4Wuk6EQDdWFh9+jwUpuWFkdygAl2al7+pgQXs
zZEs70KHQ3RejzvBbAPwsmImqWY2h6bEcYjC4Pp++WiNVn/6bwuXTtVFAhhh
w+gB+rXYE4QEiptC9Nlg1bVfKIpvLJJ43/5YBuzmp5YJx+Ulzm/bNeQWVGLl
zPOPGlmwzplan9eDw3CkIcdyvojBwWFX/sXO5lsOgcSFY1+Z9BYG953sTGsj
Tur9+l6C0YHySKQbzwy/9rYTO2o7TXLCEFbaOFmgHH/LJU7lzSW4ozLD2tPe
814JP9+5pxVAt5o45HysncFBlK0RsXU+PKsXwkJErAKcL3cmMBKRvFkEeZkh
As+A9VbNlzjgO8QiJYvPvGwD2InhOqGuUf/vjFSlbSy3CiQ4kBGF3StXfnjE
XHKLFkpQNy/wbOI3IO9Te8k59FAjIMmneTAt2uOKaRRKVFKqFn6+Ko7PYysn
GSTsqpMaWcdJQYsG/k0Gfiy5rOqRT9MTsh5cK7ERCTxyl2d4GbszPMriOyHM
G4kORHTvxjpx7xQNwv8L+zq3iL83REFfonb0ZM+Svp5oedMwGm5IOPUHzZ94
nn1Z9fJvTf0nng1eZ1co63UAjmsKb4yC1C94y3SsRzCKq/L0MVu05m8KkU04
mpsZYa34pjfi2dj7GNTVpbY2cDz3eGi6NH0y2Ms/UkU7Xgjiur3fHCHTXnx1
c8dwGSGXxn4NXMsYlFMqlhUYAeJm14fmTlvz2G2rOuUXQe88P+kxP/KagGQp
Jn5cqg/fnl8OApF6XQtBjYAROj8yHiQzUDvixjXkshDWZaTmYHBpbKg657Gi
Cb6eMvN5O16QJSo+vMkOeWKoZHeHc2tFOdvfas6e6Rz+ljV3NqJc3fsNqfAF
8lkyDtLi0OMpIMYKG1kxhEA+1bTjwVeSA+tE6dNvVNw1x83bxUEQil+3hB2x
/zW7BIYi791VL+r+b39wmq+6BBc9qXHQQ7MYvEfus+LXAJ4H354V0oFSJvn3
+9gyLd98H/kJW2tKT8AfERiU7Jw9uMUkvjx06xHcuvCg4mRhlWFrNskoHobw
e5a05HMsxsGAV+PaFoVPFfZavVU53iKdwlRXtXSAeDvNRX3NkTKEYNXJAZad
rb6KUP6sVFBMYrTYWpRHHNpHSQIIHVeWfBgYG8ZkBnxiYLwDl4/4PbGQjDU+
c3tkTBQgxFcln+PilCW/gzDJou1ls+o0Y09Z6zsd/Lt3rCeZNGiKwZ++Qytm
bG0kdUHSrckhW+cjMN7Xqk1tHZxvHREvvxsXtxNusxFjZg6W4wMfzStuh4wO
QUXaGKy781KmyhpeqFZVJa1cw9DQo0X4QNMuekF1b3SJDGpQInzQJO4DY48D
yszXqZDlMqMNrxT5SHDrQwzA8Th8HbUOPjsygB+S23vDvxWn0A8HU3g5N1St
sjs2aWF1Hz77r8My72A8OUFbHqnO005w2GTz9Sb/w4TrHonp9YBcsvhXYOVS
KW0YXeTrUkvyZRzCXqIYRKUmZrapH1oCcrJq0iqiRPAZS/WeuggqzBKCUP8D
NBfjsQiDCFzN0A4g9h+Sxp2nZu9d/pDDPMILp9OIs0kLdwKOqmyDhMcKrSOV
FGgAyUzwCgkRV+us/WYbpYi3hLKScEiKNeKS3KPJNGT8i7bJvzqlpICk8T98
lZ7GPW/iooHCyVPszCTmYBLLvd+Vi8MlblX9I2QxC+PHkpC1xuAKTFNV4dov
B9ZE4PdjNWyqX2RKYf99fcPvHN1Z7AyFXKm3fAGkn2/68xjedT71Ew6E1aC0
8b5B5k+dUQLYoWRh2PeDqYLEStIsY/z8ZAgbm+uEUR1ttTzt5Kb3jvAgWk+G
ff71kaqmZTM7ChmgP13B3Du+DAnILNcyZd4ZawMboyRw0SFml01gXSpkQO9t
E0cIYDtl4nw2IdQQqyMtiIngDBWzSKOlSJNSwO2CptCxcpbhWO5XlpJ5N8gi
M1UNnzW3+I9Lhnow+NbqmVHRiyK6MP+oMBbiTQ+1trlBbyl9IqWnLb/LKUqt
Cjzo1o2cxL6hAxdQs0+nM2Lz2h3r/y/ac2cMBEiaYRLwhA/hMnEpxM5XdwUy
oce5B04cy6BAf8WoUbsvo16u/4y2u33iQb0fI5+pv7j8zz25qlLltwOopMIX
3sbkMlgv+GP1zA0n8cMwt0kk2ohiSXxRKWTp350/rpwP/iuRf63wZ8z3WySZ
CqJigdVYdLqZ70fjJUiD60UGg6v5zK8jU4xWF7WLQ9bGku5t3lBW6vylKNDk
rVCxXaD44S4ILk1gbWdMNqvAnjddev2C1qWANSdSYSJFdW43e7x1bQvki6Uk
TUCgLxxd76dv/dx46MI5dDl47GQaUazsFwuP+b3wyHc/f82vOshY8esV65Go
xOovqnVOoCpyaohLDk3+tU6bX+p0YbtM1wnhWCyHDYCopGu546u8JTaxEPsz
iP8juG5jsSDELMof9p6cWodd8MRNiaHvu0BhIvXlgbR3NN5g6QnoWX0DFchm
JO1q0N8RobuPi0m1jZmWDvlKJL18+N8I4oVfqqHHaviXmW5VeBCkSIfDqlWO
DfVlYjB0hB/SDQoMwWF2FgzhAwJL6/+xhlEXITwXYxLF19jZ3uNZmo9MhgEp
T6NAH6chvZf1m5/yuZ5NenzW+DTC/7NYgIcBuCrdYSvWoGeZT631ybdzy1zF
Hv4I/lA5G+u1f/tQzSQdGhfef/s23XnFNJ1zaW1Dkpdx/v9Bu89QTvPx4eHq
7t4X71NmT0qs/xhPEMRVPaZ/oULFDjWD9o+ZpXvQHEGGWD/yCkW6ux9tGO6Z
ktktCwGn8NlSXOUTLcim/Ov9cfdpO3BPPSgfiN1fe5iudbQWyGNBJ0aLjF8A
EaaBZxJhLjlb4RHX8uQPk2WnXJ5rNFUOQ3O3GA4w/oJbcwVwBddRhxT5XulW
BnX0AOrI+XmpqSsfcnTkBKLPsk9SEb6o4Xy9U2420AY1/MfPLTgRz3K9221t
IWQpYSDTu1UzvuD8kbN7EEGVTId0D60n+naUA06HhqiKKvnWAk+ZnVz4RlXI
rmnrQkb2UPXSFQLz37wOBLdlcfgRy/joa4WmEZYJ3CugWKC7WhkjI2UGYRSV
s7WKa7UT+m3VMzk3tWUwK/azcybUON2Eqn++Yy0CRyOMvb3CF4wYW3SBjEfI
RLCrEpnFSWr4qaqi5HAbOfQvmsIIm/3LvR2dg7LzpuEgOtAQ7lh1tz2sEQRM
ZV+m1vLX/IHTdbUz684CQ02WRSyCh5uqq62FZIsstJgOEBXPcF4Ju5HSvLmN
JySyN31eoqyJzl2iUdSxAsRN/BDr+XpppjmbYNBiP/mjhsivV/xv3H99srMO
roI/RzifVa4GJqFWuKWxg/AJUme5J8wgrKDJWmLQtxE1vMNGlNJk1DCFAewr
Ix3DNhI5N8Ak6eoNjKpttWnZ3BbqEELT1U3mqgb7L6q0pwqe6Za7f6i1i4nN
wb8vQLN9BpjRxwE/POWqZpewDFivvjP1eTV3hjcyko5yaM4yByL11l5+txa+
Llswihtxc/Q+Seu0xFTaO0wFZBdoknOWUR9b8qj/GKmCQZKO45uJ93zur8xu
BiKAORouLA4YqKnempB5sKOWJ8QmI5hylEO29CHFL0jiECoI4z0+/CQSCMdP
fSoKkJM0k8t/L0Ozt7uvb4v+zMTELxCRjVZOdP5wHs3Q6alHXK24zRnllVfc
gIwR6LDARVDUQirYHe0/b+k69L8RRMu87krYjpN4Uv1AkDXB3Z9JGEvlujJq
eec48YWkrjL0KDO4N69thuuImZ2Z3L0VJetXmsbZ5YRoE7C9KVdytoIZ6BMW
UVQl+fcOTP6/skXlFWgBMjmWGzqQKIngbNC2Tv8sjJPL9K8jecL8Kj6sCzgI
s1/5nK2/uF07xHVC6tFaubDi6z9vCJTUiIDPsXAr/Oejxe8DnHUuPPGdNfVf
4Z7GTvtwOYDMPeI+mxI323VcEfBeJGL8qvL4UkeJufEwTTlLMjk7n/WrH4oL
eZrsIFGeyeE9tLRulDkUl9K58L91gbsg62xHj3THLeu5FQ8w3wokOZQZxy3L
H/CAPBCIdGe8i3/xtRziHMZO8HK+5seAoX2/qOlYDGOz2X7ueZX53oIW1+LP
G/lYuw1ve18mdAfp8i8nTDeO6+mnFuTc3ZveX5t+GSSkKD3UNF0RYNwPfgjE
Bu8D+gKw4m4enlm7LfHU3eZaem18SJwjGzpqDKTlr8FVNJAbwmrj1fcL7wwD
hZAeP5EqLWWKwghvTtthBQg9KYZyoCOP+8tSBSuHJhr1vd/hC4OVFpvLCGY3
+j2fKg4ybk7Xfx6yR/LVdSbN6UmUif0ZM+mMzU0wMCj9dRhUW2AtCLXNc9H9
6tnbfn0O4de46+sQLNO6Hus29EEqWyu+uMyOwe2Ys5lOVzOy1oGaUU3y+wiu
MaqH1Vk/Z69PoirlL/PyibIxX8s5S5ptWTAw3ouuoDzsjxsEC49GU2Tqks+q
o93YyKFQDq2lanjgbEFV/zvHV6qAbwy7d0/Sbd9+4gQzHwajDD8qfnTW9g2g
t9WJdKemf/osiJcSwuPkc5BdLHzWehmnGzsQwwEWEW6vIRiNN6eWPQDwCsPi
W4PkGDFYmI9Zzaot/QQ+xdtDhl2qF1YbTxuW7SdSQB6pXjxnmx/z/QuyNZp4
SLiRvYbl6j2duG1bYo5xoBDY3mxVC5bGL+gLe10AV76/S4qhRpHGoRj9dOl5
N+p15X0Navf2NvDS9wtpuNxqc2sQbwS6Zi28DKqNV+0VPEoFSiwjS1l3D227
iwtbPQX7wrmGD8ab3DhDpHS7rsQBMM6Hc7d72eZsAWMCod7mQWoJkUinM3SL
Bu4E+1CW3SofhiSTtFqBOCJBpt+Y98IeZMW5N0SI8lG7fS7DHbI/yuqv6PiB
F2OvHMTMmrjm0MkSIvGaFtORunVEzuiRsw6ZBIMpkNbk1LRDFoTp5+AWDyxJ
FA6mcdRv7N4KZK3Y8lyi02PEmFYhZkebV7ZC05mGWkjrCRh3XD4HyXc6K/fz
ymHJ6HoH0tNCnHWUmZiBzh6qrF8JPFmCDO0MlStqMy1BEeEcryYllujwt54t
g2rtxUWzA7Een75+tf8Aj5De6PxM3HLANILek1xkJmXr5qRCu7FleKA96QLf
BnQjoF+2tYaTFgKyo5YUPaZonYcHUpmbjhRcmchDTM99sUEQwvujcdw5eHb0
5P0Vc/Odyty6696sNhKx6sjfXi06gOO9p8pYGrReiUrpZt+54I4/DIX4k5Fz
dlyfI+Q4INXfkCaYHNAgWa9W1k+2XMNXsFg+5Hnaiy5OO2ypInd27R5/6kzv
lF5f6Y/1QlAE79tRf9cMqyypxC+zhjAPWZwx4tI2q9RIjC58j3fDnBD1czE3
I0/JwJTbQQZ8zG8U1Ce4rkYC2jINHXEp8BctT+nTVbhlyWlsh9UBujnCrgSz
3oeJDNREPCvI/F4O3ZFNcA2JpdePj4ZlXztG9RJUMik8P0iQc+uosza0JJuP
6fDXwgsNfbo/m3tg26sLXcVhnCZdLhqXIVSkvtULKqJx2bogKsXYrrS4wzlP
ZTD8o+ZYjeVSkCMmzvM5xCxquWDpY/DpVpYHVp7RoI7M9zTiGjoxcnQr03W+
tzCMlNgefF1dRc2wM9YVTaLlDiu6QA0BMGzozj1XqrLqee5nVcZuhCuTSv/o
xFspYbmtoLo6gfmOU0b88km11Q9xVuuZvys8XW4E/jAlwtPEmtV0Is1WDM/2
UPq9Ah3n4MVsD2dsmgA99LQjNEHxEfYjYhdaAYV8vZHzfURNdVaBj+r4ouZe
nPA1v+Hug+OQMZMkfJSOKvuRts/Do8pBr50CwRJQ532fwCNjd2VFy0RVArJI
2dUDf9XSHUJFCCwpDhX6JnXOvxTTK65sVcmMlnBsQwS9ZnfKj0Z51O7J48h7
hu+z6JlyblKB9/+n3ZBKKs+6+Wky82aFb2KBdGaCwwyIJ69nCNe+wVH7p0Ke
RLHgF6j4dt/aEzmgIfhcRPsrQBgVAcQq+oyW3kA26R7DPJfRAmTBnKJo3KTA
ey1LeJyRL1MwxrWaFv3ogjW31triYMzG9QMw2m5ztYUFXbiutfqwg6LAXi16
imfKyDfvGYPhnBtAfu9EpxI5IkWq32s+x+qru72di4et5bI35QBHT8yk0fkE
L+HM4nSh2TB+erY/U/eCzWT+huFsGGb1GPIC1c3PXGZZtz2WxECWWTQdBqcL
TEiuHGpEnhKiIz6604+WBAtgR/DOdUrXth6f/og+QX3npwtmxk1bK1+X5hJn
JgDZl+X4NtZ7eGMbMMJ7qO3cUOC1YuX0jzgL3oHkeM1n+spcSjeOcuieGHSV
NVl2GkgP90+wjMCEc3m+GBA7exKNQxUrCMRIRlNX64XF4iWy+lWdS8qBka9S
69s3AOwnKeIWXVasTTGgIPouC3isbKbdssnb0SN2rXduQ3vvECDKMEqA9zLC
6D1SDj0mAnlQidYHmNxaJwdx88wFwEbRaSNAHiF6xMc+gbfq+q/e8Fn7jLZG
nydohpH8PySzwtvEyQRcKprEAXVlGxTioxNnlRt5I9wsVwy6V8Xlh575gGlK
WdADwUHK4eOfCpYtvH2u9QpoWqzikl/Asl2aveOrARuV3uULjfDztLpf1P1G
y3Tygv8PcsEQCWUmkvztegkrfGS6f2tabh0lYZMeURnW08L4RLqdtkhaiW2X
Yi/RjjODtoAJ+euAjEglTnwgNOdl0YrxlCCs7YztNhWnoamZLNpeOBsLPvjm
/rtORcIAWvMNYx46cGZn2XyYwEvOEm544Npz1qt/K0F9MDOL774qG+73O8x4
q5+pLHlkU+0kxNiMMUNxk/BPLTL+QbZQhtZWc1SoRFN3xR0LhmQmdvWUqutd
A6oh7f0G1sbPwcpU4tFAmiMtktUhmNRV3Mi2W42TCflzW2/SmKnpKYDRElrO
x1+TLlSBKH/Din5j+G44vb+YCjZ+mCC8XCE3ARZyQrzOFP9p+4tu/kxCoIu4
LSvNpjELxrfNxw4jXycxzhj0SmnN2h6JbUDVZZbf/4yW5DrQbfekypdVfp/y
0qQ4PJ4e3HY301rZFgc80jvy6JqJfD67uf05Hr9ISOJd+o/LXiXeHVGA26/j
n5mFDSYTwHjUGLvzoC1+Sgosf87mrAMZ5glkEzP8queoOGBbgzL6zPHQPyOB
3ttpUonjfShD6EpIywVuWnJ8bz5iRrkVCxRxlKlLsNbgn+gsfq3Dx5QStM77
wY1U6R6EwBt+nfCSTpv3jNTM/71NszPndIDLkol8YA43I+kNq+/J/XB2iYvX
TIR/V/Dzwp5EKvyjIACTs+hzXWWMQYHilJDhp5XZ/bskGPmIz5NJlLnQeu7C
Ms27yUpUHBbhgmZw5xVhASoW4Cw+8lnJGirD9l+pKB1Rci/5ozjtbi6yUUtT
C0ubMHCMEgOPnxYUmvyEJ8wl/lOJ2CeSPeN2oh6y2/vH0hshnhnP1TQa0eX8
6H0bjArhZEW0VgSF95lLCOV5FuzKCMnNDtlC/M1/FkSFVqMXw7LOcvKr1cOA
VrSsMVc54Hmpbl5Rb0eX3KnGavzkC3mXaLnUNFER7J2RIle5HXP+INOEHN+m
U1mEzcSDqY3kU6Y3uwpwN6/2tmxRNoH3F/4w26+zEB2SsBIIl2eR/oosTYNr
jAJpbmZ76UeRrq9+sE7gWxMIMMg/pT+ddiZDIYDS+gVf//GikpgNEuzmN6Td
3MavO82NHGqi7Vt/uUi0o5DRpz2NEsunV/ATj+dqZFTmVrwgpULMSurRq0PX
ymrdl5ZLFW4mlWpJEATpdR4RKJfigIvP26OxrGqoReS8HtyF8XF0LG0MICNA
AiKzlxL2XHVNU9P0PScveW1IVhJhB19PtmBGVX40ZOE2pYJOQfG8yrEdGARR
B/RiTmLeZ1zPSZgkGoRG6C8gxFjF+JVneXBRoJj3d/SsDMJfzbqLBS9m1fbU
yNKdyulevW0T0a7m3rsljabcqk8ZuaLvE/vKa5jvfIOVmC+3tBW0rsKmhfQn
opTmxRz6OdzmNahFnDNdGXtElvlvUzHsFld5+y4Z4XYhHfLuFg+KOi2MWI49
fmdMZJOER3WGjcKXpGEEZb6G/9/iNPNYubhLkw/CjZ5rfk9IHr5ZogNPf45p
ZXAF9WIgYozMImBGZQ3U2Cp9c5QtbIRI+1+lwvA1IVrIsj/DUY9c/jhuiiDP
jom8OlfoNMTimE3Ee3hRICX8GNHCXM6h9ol50vPcPy5Q8A/hlbFfAotJQC+N
YmOyOhBKbFue8XADn7RM8sBcdoxXfBt1xq2q07lo+VklGNZMRjypDTAn+P4D
OQvPwm4xX6SULIMY9aEBLsXu3/vS/28tlITmXrP5u6eB8VbhuAypW5Uek2J1
q0zUHGUwvDTyeBWagKWm5vQjbDdnxTv/b28nCE5Z6ngq18uM6eJUcZ+zmDa7
TCRoVc6yiwUkUR0feYalZYYega09uo576IVWaSchNKG40qvr/gBP367j9myB
Uc62oAtmgkitu/pXLmeF4lKcfa9F6sQIE6bpy3Yu1YkYJ97wY/ifH0PdU0lH
OMFe/bSvyhN3y/NZ9q/hFeMuMfhQ+qZ/F+M9amcLIQSn/isJgZhUO5tES8lg
9QI7dwqng7nwXJPa/STjk2DZX6ThE7FGi/2jvgHHdhkPDNagik31diqBH/Kn
Ekl0HaAdoj28cwTQ/Z66NuVnCaH0YaKbW8p6W0N9md1UcNwEd1BLPpKi0gFk
TZnHgrrp+q9jqVVyjeu0ZNfu4rrpRunhweGVvF7+ZUr4xj+5xM9qbi34z+V2
G+rpRnM2eqPS3LnyWeyFVZq2Xv9rWC+ietKEXnMtYFX9G1Cxkf+rMZRUWeHs
Rnlyg6K2dwlaI4yfWU0JwRTMeY3ayoA31HU/dU3tmTfpMkRSlLfP4yAau9WQ
+aXvUrSm266A5Zc0X4RVSwoCY5J2q5zlwz+RzjJq67NHcdevT1rLDuJEB/pT
qdnEQM0Edut9aL4jwSKpaH5aLhgs0xz1Y4vCL+KptG7DNmIaPvtf2skbDsoE
9yYr+LzUZwkn6DRQ0jChvgnvPuqcohWeDf8jTTwdI15y5RrFR8d5Bq7M6V3A
xIYFHD79jX0DXUsoC09b/jeU91dhTNaVR+uKPdQsMhTAn1LmVybo6ZznDM2m
9dp65tSZxp6Ga3LovrlUIhV6cdU1/PkrR1X1k/V8WO0uEm95cn+1Ojui46za
JAQI9tg9BrxzOP422ujzG6kg9C5O5GzohI6WMYLE5o2x2LvFfBj65oRlEiwM
w+7vnLXZW0aWY9YAqHBlLbVhn6QqsTUSfBTctCg27BQubZpgipFOFizGqb0i
m2Z6z8YbFl3td1LLVINwSVaOzE/Ds/nbJoR1gnu2KjmyJFcCIGaB+w9g+ZHY
SxhRB+VMsT4I/0s6wAL8v7j60ghv/bWO9EWdJFYgrIITJAcy/A1QvPHFfv8i
RQheGDL82I8+GSmeC7TLge/27iXmC+kq2erWd7OHkxNR/Tq/NAPKaGt2svHe
3PSlIl67x0pOrzKBvhwcJQvfY8FXa/IoRpkyLukq44yqZfo8l25v08WBf+Lz
5quNgaSxqXvxrwzBAXFiKW6k9W9+NAIlqgauz14t9WKLDNT0mbDeWDaBS5wT
lzoywlwXQYYMTTeeCiSHWl79yC9YwGF08tWdmJy0QxdL1tloBS+PBTHoQpeo
T5hfLAVrfWay2EsQyOT2JfZT+MA3bEqNHQUyX3qbRvT+Slqh/apgz/Q5h45p
CKvFaPWp693mdew6q+ABY7uZVVpIXkMw4KtIloMd6r/Cg3meRn1lbWWY1yZ0
A4+/q3Z4apVZa36EOjB7XCQZdvyEwAn59erYOF0Y6+VqbWiifU6cw8tSZPwo
LYZDbO8DuFsB8lqPyrLFiB1hz5RTVqZ40j37nH76BopCwzC0Gw2NmqIgT4DK
fAcWDxZvETwZkdK7RSStz34Zu8oK/o2AOZC/XKqg82UBBkeg8ummOIHLsYgT
r0+HzUhyy/WMJHEHlpGcYlvU0yNyOX8AMqoBmlZMAZkfP614CAaY4HxbN8AW
ORF8Fzh+q08yMFVpx8DMXvggxlxur//UvAzr6wosMkJSj5/GBAzNcaI8XCqj
7qnlcjpzlkEQ/ra6fgGcPtbsoLectgr3TgVg4YY1xEH9HS2qrT34j5mcB/i5
lK26OftzUPTDt4YdtP9Bdk/v+VUUHxNLOHAAEj4vAc67JF/1ac1golBI6DsB
poPYT9PDu8ZhJt/kNUxlwaU7EWNyQJW8agS/8LYuiiK0yMJUtxcPo1unK9Ib
CRgZaZsLW8g02DDEMPXYxk3idak1dZUkd400muhJ4wBR7d2cZim5xR/NiMyN
nmILsHz+kBGZlQRANGGCcpFREniEuRbWcqB5pJJimxcN5NbsNGgRMrqBSOp1
gooqoWhbp/1vcLPyvMtGpKKD++4vFErTDIz3lKJ+dElQ3lEQOZCYxk4V0KOG
K6njf936CeHhkGklvUaIsz3jcmP7QCxCXY2wHAFJMS6RWkbMxIbeR4wU3OcA
VVde2CWskJnv2QtEyrGUaLJ1URwW7hYGUojHMKE3+kTGIXM5ZEvVBnX1bom8
EoRXIhuAXdrO2atTUA6HW54blrmX0QPmLHdB3N/g4IFuZfSuqU5tYUP9pley
a341cq1qXgTFpiYRLt0nXWUo/MMmgwIhcfQ/9OATbThp6yRbSDBOHAhbux6v
sTlIr3qUS121jKNRcXAoqfL3aZmjh4yVyv6klgU126v654Qmv0HQ3s3Ygs1h
a42SCUYxv3eoiB/M4Anug0TObovjBdlFelkLInq/iKWoBhj4SyNEG4igOtLw
ohmC7y2H/wJJjAHCfK6faBe2bZMsdUailp8Lb0QlI9V1AtUJabWr8J00JHo3
7/vad1sBv+5waDcbcxkpxa+Zejbx7H9zeDo1sdmlrJJqisPRiR60vieOEUC1
FKsjFHuZPSlD5kQRlN3fTFnuEZUy3jaeZc5b5nqzSrN0hVYSaUMzIG3XBpLG
xud7dVFxhyPTXyzNmfE0TJyOZvJdRPfzbevBD/x8BBTYIt6/mBIItWL4RTSu
xdj0+zZJ8QKpy9IfdpNrCjfiSd+cmN9pQOLxk/MKwQadpv67UBa0NbeFmnrc
gm0igz+W+p2NqH/8u7jlEqjPfpNLHtmO980avD9EcoEDGTtuDgHrPqqtOgB7
TZPRstqSBf708qsgXh5E3z0Zry7fyodTnz3ZX4PjyroB3RY9/RXClPHlxcjl
m0YNtXgQ7yO0dg5ZCIxZgoZFpQHgBhuSMuBcNKEesn6INg1uGY7gB97LV77D
cD9n89D45Q6Dh25ipgZ+uTo+qIQSfQYBnecsaDDf9c6YW6G35ntk9hd9qzBj
ItBq/OAt9L3voqzGP/AkP1lmGwyGDfUJ+Hv/B+OF1FdB4IYckfAn31TJ2OTE
4ENfYUSuyW1pRMlRrf6kcR+0F2MTXl8gU5AVvhSU2WQZgERKakD4QNEzL8zz
nuI0SwsD1FkbQdDoTfYAr1TOYwz45jK4LS/B5oVKVPGYWLALy3eqfjAuXdR8
L2XjaRYJajrfWpx5wNK9GeUd2TRR1+ypfn4UeWFU7mHjHR1otIspz2NagtW9
LMK46YNOBZZfGHst6oK/DhUo5lyzkjR2L0mZemo9H3OBkUOXxx4Fdnwx49HE
MVbfzAy97/PO7b+8jhytrt9YMJ26xP3LG5Yd5AmPsHTCyKf6OeDnf0FOmOSe
HdaZVQZW+mBjYarasPDLdHOoZ1joy6LfUp83jfDKiZWhhtMonUtPODsQ0f8/
3zwqkP8JKfCa88lXNI5oXjy5E3M/3AZ+UiSTO7y72m3cLbvA/30UfmocIYfJ
qFFnHM5gcFbQ+64QEkXPlVJej5Y05h2TkinGdSWSpNs1/KiQOFuApN7Q3HYp
OtP66mFt6QTGmrCg0h20RvH/ZWoJaa1z/hJjjrkZFnRpFzCAW5/LE+b1EOm7
y/ZQ28PIgiHuvc8wQMujk0c9JDREEsE30IgPXi73a+vbMEj5u8iRU7eNJJ2I
FNysSSULKynO1tCRpuVRABHjnz7Hzii0YDZ85i8bHa+1fJr+a30GI4zs6jz3
WPO15ovBOdtYZ/cnNkW2ItMcJKQIstSG9X6+8YA2hjURBxrfH5oOGdcmI/ef
O0s24X2EgS/OZDuBw+jyAabeznllc0JGRsaivxLChxiEaxkbxYDhkOV7FigC
TrMMjDPi9bjVdIwJtDAJLZeLRIzv9GhvP8IfXOjxD2trJ4/rr4bxpmnAyojn
mZxKN3R+JWW4vgCVWPEj31baIiTI+LDfBYLq84gyHt8hLyyfIVDwVYRY0k/L
KqAXduKTOnh7HmXTaa8Zqp8x7oXpFbR2hbMD0ajmOSf5pdaUYsBqOo91B8ev
m3MaAgwTsBT0b+9h7814QYvVagFD/PV9j+G85y2t0/QH44Es1jb96xqcFowX
A0JPptIuWUtOT3acS+tX27G/9JGQd2cqVCS4RqkP7awJqvApJ1CBRETQYXUw
O33Rh9iIsZQ323rt4P3udeGQfS469hf2t82LG1+M0bvumDJbbJp/oKN73lUz
iAC5GpycrLtvPdYaibKb+UllAOuDG4wKNkJ1eBZZKOlLyKcvzKrSHLjYDqvY
sUpNLl1QSes5u4UsWU0bXqLu8FStTT+Q875XPGKVaPS3cv+ivrRJVHmBQETR
JvU6JkBJGu16M3GVUnSjUGoiLrX/ZpNJcDXqpeHM80EfOXx5lw5Txpxt8NsU
nITaRFzhUSUA7/xsLBV/+C6oDnDeHJeRaTG58okgAjGwt5L9ET2ALcJolmlf
xOdo+bW7oYwmJDJTnigqo9Zo2AsgofJCIX8KiJMi810TvZtGcDrCIFW/ZyZi
6vWSyl4whOdIWaZvHgcR0J7Spi46QBU96W++X0//lASb01l9R5Poem5nDb6d
syvG5vQWS6sc48aF2Y8UiRN0DM4Z3IfMZCaKx7VbokXrkM9BnDhgr0eupz60
0Ybnt0ZRefggR3HhHtd8GZNSDQ4HW8qO+cxTWdyxThvTpyi1SDsqIWJdrPjO
0If0m8TVHIwdPc/wNyNRJEYu3ziyVJsJgoVoztSHNsmf3O6DUACLfQ4fVVu7
GuOxokEGi08PQFXZJZKtTW1SFQTEDCLOlrVwziaqh/c+LpBsZjX9CXE9c3EE
r7+8CXplnP+o5ghB8GhPal7dYgNJqIWyDNpBSjJG8nxduc9RRga3UcfR/PZ+
m87ixgNgdQKDpB3916qwaZVdWfGckWgnGNaZNMd8N6rLjrYKCrOFops2XWJ5
Ri0nFxIk34Orke/sHE1I2U/EmmO5HJY7s8B2sMZXjIpNVTKjRE1QY3MhO/jD
b6xX52KLV+hTaMbl3mWmjHD/ZrMCcNXj8WCoToFZ+WBg2qD6M/0gxc5byGQq
sMZs+tKMH1jUkonEeEi7PMVQh1kkb9UYdbaZ54hHTQoBpO/jtTemeqM10pyd
+cscPTtGHEuevCSaWqHWnN0YlXYaLUnaDgcKxIM9IPYIHYseDVDG9iKp62Zx
8d18980kUD4YykJi50wnjZ/SFdYLGi7xV+NUXKn4WskT/VxaUmDBHG0w17wJ
D29l+GRI+fHybKFf6E2oVYatNSQmQ2X3MPGrjNntaTudRccKNdtt/UeEjN5V
l7PzJqNcPEvEfouNjiQhXWY7V5vNLA0HT5WGmO8NNPDKk0xXDM7ztP6lLfaB
n5CGE1p8iJpX+hpZkaxFZSzA6RUniM9kOPtHEvcaXvwqc7mJrv/FRaRnQc19
C/wtqVuXcpnNlCApmPZQMDHJpcO87pNXCIUQTnzAUQgUDdeA5GI8gx4AyPv0
TSv3kpWCHKTLSw1E5N1jiMxxXq5Lz9bah5kDaQ32ghjAP0TeUJzWtCy0lHHK
Cpv1xMfBFN5u3UUgQ0J1t+UD4lZhfyhYdWIHhKEAu9w/J8wdFA1MtopL5F1S
gmGCB9ivYC2YBfpIHQPjMV90KiuoZJXIXtzIH6WYt70jHQsCK2kD9JkW9AQe
EQVtFP7D2BCjKHmywUL5Kg7YkqWfE0rRC5G1VfSG2DV7EfEI0KSYp1viQ+lM
wgMaQ3OvLv7tlwFAWnJGh1BOTJ+iE1+x/daxkqssgdzPe0kz9Dc/KgKM3yHH
atK5eOXEwhKgIhlpkE5jXlnBVVo+5IjfHm9u0SQV+S36a1sy047lBDUbcQvY
Ic66E7C8Ams/LgFwAuWI5POnRgHNPrY/wnnyFul2jActZ/kCvaTUagCzk+iP
qghApjAh2fW5US0SdXe79qfSfd7zDvRmUkQNsTWX4n4CYEqndAtiBgQ4g2c+
L1K0MKlHy0ecTykICIoJmaXTADA+SbkZ50mvH171llovvMuORc0fkqYS0enz
BA9jxakOWrsLIOSd2Ds/0JXRtE+U5USIDpx2xwQaxx0GGSp39baaBELTgsP8
L2ncdk+GJktmEApCxEphuOH6CpbqZ1rFDMF8gi83kZ2GnueQZAIwZoblIaYP
qQtZTr796qneoCqQKwStRiMYiwS2q+ZDDpADDzulbw6r25yPNyQfmdk2Pr7E
NthWZgnPnnYfINFn9H4ZU8Yn4G96kHGfQyEbk1VuYa+ok7xbWaU4OVuwtbjV
wgc/c2OglwuPvsFkqDgAGZRs17dLDQwfzxdATY880T4U7TW36TP1LC2RFu3d
G/ep9n9hKonaCK2pUnt7dYgTQhOB2heEYjmFNX0DY7QtUNXRbF9Cc+u1nNyS
OVeDqQeEuvSc1jqVWgtbm003mVSGoHQd3MF1zAW26toFpXLmYWw599Ggo8ev
C1SWiTl2FpdBVBjrup+TsazPP3IDcm96/PhlWH0ARSZZ9mvez4fAlVo2AjGX
1lizkutSB8iIhoCeFPRO2Yxnulyde/fNLenJamOGjxPv/tM4yFSSR7WujL9S
FMgTSX2flB97O6H4QUwctTpY7Rj3B9OIS1IVmrOO3crNNWTtnNk5Evjx3hxh
IWUR9TzH0f2O1sF4of/PEcr73MiZlO6QslKuEJqJpqlFo2ZQSdbu+CCB2+tE
LIxn0tV/hXDlVhs6kTcG/Svrkw2lDwjMb/f/E3FgUOy/fQbYuot/W1IgGaVk
TLB/7UmfYgkE84vIvL53JQ5Xbb2f3wbSh3Fr1X+uwN075cogMltjGdR0yK9s
JHQPHbHC30io0iFnQ80SoxPZkfPXuRT/BTbuHcb/P8oNLggAcraNt5EP7wsV
pwNLWDkeDzBYPaBP5DwGl4ZalcK6zzsTjZ2eq+MeCU/yU2N5agobudRhXWW2
wk4/fLe74GaMg6i/NMOpabSUnSmbDg50v9mZ+FCaCi1eBcOKFyI6TcvspzPV
w7t5Q7hhmi+jUO31pYFRt4ZTbox5rr1kCEg/E8muntNdmxfzKKApSwOhrDrU
0ffZElfKbC2cgndb2+94CJRvuv5zBWFITvGRDHJ8RLjtx2uEV7DLr7oU8hyj
587C5URckZJrNmqVZqYNXzO21wFAl323ZeendyV96c+0phfJz1V2vLP5OWn9
/QbOLcqyQDmfVsbN1NdXPZNFQALwwfHLRNNGbZZ9KbOJWpv7d8GpU2V5wIE5
HJvEqRacrlMqWkYjJG+BzEdBe8VJz2M6ZV4tnzvq75sknYeLudobOh89DJhS
2a/6D7Wr/ulOxk2eyQMWsVQWoT+dczTwu10E3fXtyAUExTBMF3EK+K3BW+Sy
4KwKAE0EG5aFJROkU/5LkwnczlC94XG3bjoloh+EKTL1HTLqr6O2ghLXZu/o
ZciMf1xUAnejcdYyPzlZcIclIWDWZQ5kVMaJrfk6igsuxzWrNpOfoj+eIY0X
yRKUagNKeFs6XEGh5bUHVWAdnEiXP7yvbdQQ3unpXwrCc/tWF6h8tTL9B3Ns
Hlpm9afszrrrZYNUbvyXPzXX+UiGCyRNRIG0Kl/5ex32QY4cb9n3iI6HiZQ7
xn8qpqpx/hx4X0QlA8UyjjMpm7rvPuqi0j/zQz7GlVNn9lgv4jqedqrjy3VQ
l4L6+kQqj5el7EjdgJ2D5PqiW/zWt6bRcbxMLY/ls8eSkefbXiSffvysAbSD
DLAUICMOESpvSHMeMWM5m1AF3gJYM9RY+NRUi1O3lolv85j43a5H2SD8i2bC
YhpBUx3jDmhbkJYciMsGTo/7BV/8Dge5xUF8bWJc7weL8MfFQtYA0kt+Oxa1
hCQ6WClQfD5lALuyBzmz6E30Ial/TD4+FXpfgA5qQfyYyf4qjBXGzdxzNZ3Q
G29A7wYfcZSbQrrMKWhGwS0UI8Lj6Ze2IeDbi9wVtBzN+gnT5o8iLuaE5aVT
COSnfATK8riu6IGBmcy5oG9/aIFQeWInvikSy+GNZIwvPj94qTN0oHs8Y2VX
ORVdDF8fUG0jkQvdeQHI7aOi5szU0TC5obfnTe4w3Z0PijahEW6sk7Qgeqxk
3iXZv8MJpuBzGpg6yI71NP4XldrYA4hIvHL+riJrdxF8V02rTLq1udYSiiG+
MCUd4P+N+fAZbPh58+5GnLik+QKOOcXQEJXub94+QDDpDndm31hMD8hjIvz/
8ekx9s7lMZbs911eryulgL0Q9r5NtmZzcuhgmrPc91XA9b9nER9OzL0cAh54
Plr5EOnQ93ZIp8m/7KQ4aiya/hyfYGnkP08DMgylvTHkf6Auc86zqXfq8gXq
vCsN+Rd8NMZh3w+EKAHQj0A0MnuHxCnvTuiwyWJMCt8XzGMVgHpfj9ijboWs
AZgeh4vh/mVTsL57QoYbxdXbkUnI2/bgQObHAdiFp8knKg776sMH5mQGbvYC
C4RXKtHAOOrGSDBfp/V4iRNkxZ3MBGHI17gTH2mxwryDA4dKHAzVONAFSMrl
BMuXA2y0cLJOUuOnKCevcJM0RgxWIYEuuSBuH8VyhSYgGVO7sIey6RBYpG4t
txEGEqMO1FEaS+Qsx1jVXKGUJEKfrfxFb7c3SRWpUXCo4dA4mSNT7a1zVqap
7xr4F2FzoJ3PLOZF62fUgbXFb2fX/Pk6EMUHS0nzlYfaisYmIADGM3NAPg8u
uSPWib6q1RjLy6cHL+imiBRdl6KZJ/SrvDQ+r2ajI6MBfJccKIh04NOOecT7
RoX8Iu8OYGfV2LSoMlH9ta/I3H5pb3IDLAnK8ZKocl6xoVASbif6nqfRMSHB
rl+K2HiP4dYjMKtZdg/vn2Cg8vi8AR3NvWoJh2SmyFj4Q3x+zoY+OmGm9LMF
B/QIJbo0jw66X6FIJKJ5Eqvxmzj9rr+9ETL9okywhn+k1SYHfTaioMTORIdE
cT5iE5a2YI8TjVyStrHYzYzBX/I+PQFaMHjJlt+CV4ITJGae49VHVYdVpIsH
rB5YLlbrVfjlibZVdK3Snw12LSM5ybyt8B9+ZFFB870B9BXbpZczcWIlDezN
YxwwOxyibzMEFwwAk0LcorAOjBTC/L0vpnfiW6rgOHhxzAwZ1VXWXy5z2BUy
Tby+f5m/18/SrDyY7i2fnDNVF/ApivpM0aqxihlYQFazLazFgKOH3J61BCsp
iIIzjWNZs/+Lkyy9aCS7riELpSqMQyZ3OU7wWzJErlIurXFUF2OaUd+U/dx8
6skQgnZBkoCOysq1UN9eIleEOF/hm0gJBg8orX/ny/nu4DYBpa8DmIYxYsfF
9dE9yIjSO9YWzk+6MnRm2CwrYXqClT+X/4bRBirakjmKNQ4BRmLq0y9ZqIOa
r2zb551Wmif5XlDj4Q9nFynIyUXii/wHwVH2JunEhY2beT9GLUpg7dF10xwJ
LjlwUiSeiSWwFdhJEuBm3UK5VZrn3L6QqMD7e/pynUqvLJ4mTuZqnZYq0xjt
rONqOcW7nOP0ToE25bDk5zHyaBFU+4Pa+vKI1OktU0NvglJKG9zwmTeyKsEp
ynl3/be1cYtnbhzkKN9TIFt9XMRXmjMW/WzZFjNJCD6kueR8T1Bswor2n+E5
azg/QslAB9/ucXavlMCa7jf76zUOLh3SmdClatV5FRcunG4Ob0jh3AUbWDuZ
cD7yJ90fSatpSU3pjhaDUsSdgjxE7GgkwYL4KUlXODwpwTCLCnX/N4bAezMw
6FSiyYCMf8ClGQakNMmVJyaPRxf2Y/SLXxDAGOvMcewyOGvuV2u+Sr5hUr1w
vOtrEImezakAVIf1JpDCjLQgNxDDASoIFzfS5/GKpm3/tIJZIGZab+ZYBgRq
AMzfYY5kC1xKrJp/aLEu/6wDcUNiCjrElHtVKMLUJ3cJAyHC3daVAP4eCgFH
+tRpK1DS2Ntz3UzmtXyhtNn6kpFppX4sEzRpEy72Z54sgdnLdT4C85xmGLVm
hXpODmUgz1GdcnIovHVYpq7tK/eCYslLhHPpXIxjO5VsOJxBwxTdMIQAj+xJ
MHF1eC1IEH52n5mPFZeHRjHcKi1HYQc+3urRA51tC6tYL4kEpXk6UccoNsFE
/cLYQyrHIT1/MNAA98y5aPNjjfN2HCgcp3cTtv45aUCePKMRansZ5zZ6WIWZ
Lgk0ReXe73EHJCLCYSgrQ3vA3zt2k+ZnWSzJbvJzYbvOzyJKiRjzOy+vHsfr
erlXBCWq5gGl2SYAdzjNajW5WN4/1TiHfmRB/bpJ6CviIWAiYZHhvBxx9+/N
SkkVt9fUGq8+uBfpErDaePYfj7hl9R9Xkfk18AfIOYwqAe7eGTm+HrptU9ch
jPmS5TLoczkKH80Gs94J085uwhSHlsOUFNDksAjV6awzQJY5FjOlEW4oE28i
g4ojxMpdoORlvaiTTaxBjQNwQV7e6yxGG5Ak/0wp9L6hS4dfi2ydayTyHkyW
AsJMIHvQ8j4HaIgBdJbMzhgvj4k6E6fKc7XNVbQi2P2oY3xfDrhO6t66V/4l
r+W46UiOqaHarKf4xwkEcX1lifOQrlcpA5quKNuvezcIvMPLYB6GFZXK2y32
MlaWtvd/sb/HAqUNA0LpemCkx8Giuorn+RVLD/naB68MF/gxW7kvXDqS8o4H
aAtz6L4WonzBTUbA1J0o0QXv5LLBZsNhsByGHyemTFIaPUo9ldRoDLkFBysg
CNegbzLS5M4TcBkL/5o8GMIXfvdvmOp7m18bi+Nss1GfpwXSbNOtdmiI4XMV
ZqjLnnlQcpSacwnpmlU1p0u8vsCqnNuF9PAwTbemnwZ8kecrvMQ6Zm39q0Fb
Klo26bLi3j21S8Y5NY36dIQm4omGipFGpCwOGHC0+iHGgXu+VzEm4LYwK7X4
71BJDcoMW5TWQfcnlHZSqE77m0ExIIjM11bT5ZKxW9nnnfyN/weqivHC8gez
55/cvwzelmDpg3Et20ADgs5OVFXtXWxWsPWTtO+oNadWlxxqfCLSa2M4ZwCE
DUFLH140OGRn2e3HuF/o0X2XylNvDsXJaQdUxqPFIdrPu78oCjFfaDksctJH
52tU9pxTYLLZAglSqt5NxU1XckJFqEbxB5KW023KcW378qMCNcBKjY5IS17u
o0WTCwfMs3VdpgXN0Npk/XKK+wj+a+05a/luzTFWt/Q+iJ4Xp9+Lp4GfsrHQ
6gYsCc/tpDZD5D+KI/oS9ZrPSbYjs0ky7WF/7NaPwP7cdd9UYI/Q9IBS5oRr
5YNom5izvDPCSEwqiQOP0XaojBKe3pVxlex57CTj//e3KtGL/DJUFn44e5oe
n441OaesLnmfHISktrZpu7IF5qVvRL4iR2Yi+wd1DKL5tMyQSJpkrIRyrF8D
y9E3IQBeJtgCQym/r7QNJrBFuY3KZCFk01yeBZn9as4lwHqAwZLIymPCrvt7
6S7ZeEdBbDIm46/dV4bJkq4c7mAYJIEvK7C5C/WiqCnVyVzQ7Lk3Ny2AfEB2
zeMl4xu4gbkUm7WdaA7vxmNfBHPjiBiGEpOA8puvfk5QA6Lp308HhVhi7/Oe
0nH2ZV0Re+hfXjdrSB9UBE05UyL6ry73/krFnX/pS35TIIFaiWuHpwz5ernq
Dzg3FSUa+zdMz8i1wqfdg6xMwUFVp5KugfppiipH6As2sUMtmldtG6oG7U07
cc3EzhO5HQayVY40EqnbtECyw1n/oAowr34CjY/bREzXf71aK9nLWns9XxBL
Parwa88xXfVCKd48kKA0owHS7d6PmgAl4V12lxZi0qXYxTmALGc/TNroh88P
uOSaFr7xius6gNFFTHvS6Gmfr0V9ALwLL8X48LEKcsor5JTH+rE5ehPdA8VF
4kt1bZcOWnx8xft7LYXyJ2a+/uXotXi83Z42SvH6F+JRgsJyq4L2boR7tGTk
yoJtSID6tBQHbj9hPDeQpKj8OHFoYzdXKnxWwvNz/jdBNU2yjxDczkawugHw
HKRYgYWV+5h2yeuuNw9/osaCopfxAu9R8G0hWPmKeNNASNmJzIx0hkZ1qOHL
MYLOsOxAhROjJjgvXzjLSMtkQwJcKoXu1mu3jT72gLRLvXfNMrMEc58Be7LX
5LFz9OArZYi978mtD2BDVhGpNckD6AkqzyUHVUO2qEEztMkPTa3mQr9hBJqD
lc4YPqzeYcfDQan8KzK6O4QL5ziwnGLnA2PEFBfT3SBpR3aARiDUjlaLaxnP
TuFzZVrf1V9dOKDlGoxGciWvszqdHeMeXBjtTm0f6aLIhBwBGON3yQZTldVR
Eu01cTcdCsmDJgeRwL5e0O01/aBhTHJTdx9bJredLcyh0lFWgDbScpjGMzNN
tVczXofZAKGYx7v6Ee8qsOV/YSoSV6GPf4DfRtaWDEAf11BANAWbgILHP3FF
4T3pRWKiXwOgIY+oLd4cNHjelAzrdvTFrEqWOJ/G3ptciBv2Lpvl3d9cK5ds
Ps3RoQDA96miepJ6L/TLjA3GREobrx3SE+mk4zEvcMapof0Bdnn+6ItY8n3g
oLCSICoekRH+DSoInFxKaAK3Tmbk2YdGMI2FnYyMBnLSwCyhG6ttOx/orjz5
q0p57CyBLFZGLsG9wBp23QJfPjBlaqXnZuSV35t7SVeyRl/D+v/6FBryBaj1
kAll8nhVSaGmL9iwg/ZvwmPQR1iwkJYC1t3YbVqJAKOqHLBTTrWYDJzDuZti
z9QlY7SCOcNOH9ku3zG6ZVt1zINS3gJZKu7j7KdBMaupgPHTEPhCMWR+AzS4
Y+JgnAKrHFsnD/G8752KBdottEp2Xt0tTd+1e+YeOHrfsBK5/UM986MR2f/O
XXV6qQ8IS5ribRkqKtFGCFOo+5fh4N/9eT0Ud2qN1FzyLVxhZxcdFkG4R8qj
EzH1c7OsY9TzPrkhfcA4uYcgJJOjnElpI6o2WUYUZfqAaDtMXqd5Xc1CUdr+
vKBkL3pk/cCb4QkQsT+45Lzt5rQWLSurko0hMEjl3nysx/nzL1toAB3fk0Ck
znlpTGvJvnEcVwRe3rv+ap3TFHJxhidsJdy8NGGQjt9krX6zhlZmw3YgF/lp
HDRiiDqFUH8oJoqiay1+H+C5E//lsfeRZ5JMxDeSqoIlQQi54eN89ryq9n/A
FfzBdxYq/tREPcGcy8PBTMDrsivTqMKhqp84AlmK74q47HkBTZEPZbr+XZ6G
3ocSPZHmXSEfdLJof07NGrv+wQEt5RdzV9WJ8dz9POCFf7rteyzaplFarpfJ
VXcXMmkaDYYbBQMa6TG+HKNQmW8aRdUdU/rUWYCHsohVsXbMfYK5I/ZLu+ey
ecJA2BuIv8r/K9FBFaUQ6lCtHlhIP7ENOsC0g3EU/HyNzoq2OJnqPrqCh5BJ
+3Loc5WetJwV+fhpjqfbvkRoX3BMcKGXpuJ69PNyIZ6hIK1h8Jlb6UDzNC3w
0YX/HiFl4As8D6r9qvEKtptkn4kHdTVwE0cZU0Fkc3SSGaz4LXZCOc4q0wZO
6yCm5AlVVFNFVk3xgTE1/iPAJHAdQq6/tvURae1tomGQL7Sl0/PRpRmovbtY
aq0mhL39nRp4pm1KVNS3nfnd05xK3orbY8xcWCeehm2BknFOwqEIrowVCDfT
dHjNC+gY2Lsxfp97KKtT/7PmUMxjigYSOQ3AneZyQ3kfb60ziiKomh1X53CI
Gal+0oNhkummRQEhlnyQ9sBb6IVkfJI0bqUOtRsLYwUEZOWXdMf7d8Atl6Sl
HR6psL7T6Apk6u54qhjISiWhACYwqHo8msBnNSydQ22CKMEgienXmJCPLuOO
+dDdw2An+xgULPslBDy4iQPfWoUWrDzJk3KV4UcbSMJG6fTtjjYXxzgKwY8i
K0Wb9W6Fq2OvqO3wn4mCQfsQYV56Cc0yJTueju4rgEMUPyksAwHML/ucdnzd
EqMRmqMaiGqikJKPcR6TuJEAI2QOBzTLYIANwmJqNWMHW3/SwqMaq2IxDXTV
lXlKADuqSbUWLlXLlsz1bu1dFuFnETRpYrjIkg2DuO1AO8vtAzspJOS2VVeE
+/e84OFRMjLSfxEcMSbk7HVCXXEKngd239prrEB/ZAU8AwD243eoccs688lT
KQrG9mwy6UkV9rinD+0wyU7M3mPYJPieTSvckezqKNkS392INiugjvz04cHh
ionMWFauPuKP+uo+s6KkUwfMIwIryDyCadZAjHL0CxBPTtEHYk8BnQD/3JQQ
Kw4isRg8RoUpidi6+Wdlr6gZVHGv7oPsAXlo7uGeq1iadIkl4xhLoQbRFPDA
oSF/eiUze/IWINg8NZ9xMIKZ3qtFIHevYaZ9ditS07MYSWpu9yu9uoaP5h26
/s7ocNrqCxNx/G9xl04cS3nAkuAIKfJLqvqT9WHodiN5rO7aajxF2lhdb0I6
2dVPukJceTxOEuu/l4K2544IBp0dfY+Gfq3WFXdo9mbaBLSe4WPvnAvd1tXW
lVA/eGm7Nsc52tx0FbuYEy54kCjb+DCYS44uJO7Bz2lSRpSVoX5uQXZ2wuwX
tVkCKNMjQzJCm9vrkQ/VcEMZIUP8M26LrL+0ylli9GZ3UStciVAkBsnYVIOY
PNYUUiI/ywQELMsVF5u0FLUWnUsvq9frT1upOG0uUGR1jbH7/QrEhAwxxQb5
Zrsjb8Rbpn7nFVR8g0iKmAsWbystkA6egiZj3ZpMhJosSxUhrQ9hw0NEaVwn
absHWnUm5gEl76DAadZJTFVvnLGO7p8eu9e2az9Y6mJ1IfqUeuxCNw/+HAgl
VBPJdY2iL4UCxJAmMibldWao/PwrnQAK7mDZ1G7fCVh6QkBgKti69nQIGv9x
p7qbUyC0+OKSwlkjvv2o7B286eDVibG/lf7tWm+sPOmjDptdnJd/tbGU3uOS
/Jqh87vnepfKWW4QNbPtyWYJ+TslMTwNZKXz3izOkZoCkdj0rAAw09tH+eI2
iQmIYcnjFW2nGJeBytbj4kT7OYv7MH/7gUOgRcaBexMEK8nXIFVfsxn69tl/
TBGnsOY+ZnyEImvMo1Rkxsbsgv3rULqKZ1YqGKE+frgFp91EvmTmTIw6QwZH
NvCVY3s1DMGBgzpXjoDcAzBT8ONG1AOonw380jrO0lSYsOq9l/xQamJXDG03
efL0SvONto1BRSTjzZdFabVszTNnPI3X9KeTSa5Eb352b5bhDUyjgUfpptXa
QJ8sln2pzvwUyxS5zPOb/K+dvP/VQpohY2KaB94sAz/PnTEx+r9sIlRUMDZN
pHV3cn1xoCzvhVyOJ1QL9oIAofE4/WGGIAbAwd/83ZeAW42IjeLIhbjblQpF
liOaaZ8Q6+xN93fwB/S/fW7mEo8Fd22GacYVFoFPJud84Zyd96Qe6vdx+2ny
/i04SKVMcEoqDGot/qrD8E4n6M7Ii3sdoU2OnmDXP3K4ZkJ+1DWvVBO2B3ed
jXCv1V+M/w5UbwmVNlmqalNq/WcrscrXO83IW5OpR0f1SMWOsvwSci0lTNRI
B7lMtnAtFqOrCbotnpEL7Va7eBerEEk95UY/wydTi9baMFIYPrcXhhHvBYc5
Je8RZgATMaplrYFrxB2Tuc8bbY5ob9Cfw8k2PriFbYUNRVXhsS45e/LNBK7u
lfuAT0mVmt+PdWp7kNYGV2TTBgZj1Kg7bZCoiyCHHmy6Tv6gzfzr2pG13RsF
sLZq3ch9QC4p0QB1ZyXfcD5EeFmqvpj2Xr4t15M6CzYMoh/mTAZd8kW60NH4
MWE2LprxCG3g3e4AHA4jFi7moLfirV0Wa2Aw018rMbUXmyjcHywsHEIc1gDe
a1RSjwytOhXorxd5AIKZkARgjbJQI1qKAKVqgdyYTThrEn7XW9PvnQ5NWw01
2U6me8Q6QptsMYuKe/oOhhmm6Ap1VxW8b659NUNwTsO8N1UASkQOtoQwQCIE
YccD3PaYZk+sJPovS2SN4SZsX0oOMSx1XaQhtzs2XsOr8qxq9t1m+k+ck1hM
bhoIXvQCYX5tVDyY9hSBSRRzHKw7joPvBz3NyvbQTxtIPKktO7ZreNBOl4iu
Zs3gzlWL2jPc/iLj7IrlqD98hjX+YKaHiKVp8/Ay/lKdPLZUuwne2WBc5DMR
L9HrDKybwJPCfpjqkyQS+14WyR6s5IzhrZEbRXH3ju+jLhU2PP1cIS9ZXDtW
e7EQx5p843SgRNbfFjTMh9geCXl3GEMEuuNQQOKJcDzJfsOBMQ8i9k0GIEaQ
K4xIZC6c4jboAihEXzr44dGgU5MstN4GK/w1rA0YuwLpl/NbCcwlEl6doWG1
+EMbFdVtTM1hkoWW8r5dMW3sAkzGxU6b046ExtaRndGH9WjGOnqEJPxuT2DQ
8K7Ap4PYxel2NuBZpCJPJKZHDlNGbtIYRsbZBxfRiKEXQgGdIopT91DIjzrU
srea8TMcnpdEHyP1lktuwL7w0/LX3SYdd6YS3iZ68OpWXH3OvU+U76d0rBAV
uC3m3Rwh79FLAn1D98ZOb0/TG/xagJbWuEYAE+F4vHxyyl3fCKVaw9TS9uqn
n96K2bq5Z9z9GG3PvH8VJ98tm12DRGQ/DxDL6dh2kMM+z2zX8Aw9WKXfFC76
9tZqlksjTUEBnix5Z8oZ98AOxvFMIPk6vGI2nlChkgwvQvoUUb7H1diacT0y
9hGgk5kPs7MnMhIBbWqK/YpXNO0OhoIs5zxcmRFypdn8G8W4S+6qjpOn0f/e
uclU8yg1bJ7ZOkPnxr7Lz+r0se27UWdRvtqCjbVCjgwoUOYqntdOcQlup2QD
swIA5H9DS/ZC3/cJqe1mQEqrHrarn+pNm9jppJNSK8KaAErFg3SgNvCZ0EYM
Ty3HpuaMEpCfWedYHhYmmWa6HI2j6ngYMArABzjQ1NIFlk6ld9rfVSWzIknu
jEVNtojlPOPeQIM5cvqMEPMg+96zS1W5j4FULcr1LdoTgtsuYrhvX3Fgsji/
RTl2vZ9LhD8LsgArg3Lwzr1FbBxlIWuLDQKuM/El6ozoyuFydgILqP/Ymtjo
dNS4xYJqSWZ2nVXgzPhlZXrULxUv9KITFnGiBWTjXTxcNBk/Qp+SFXik6ppW
zwebv/ubS97v2AMlss16OKdCtb724S0X/JRzpUfKecOIkdslV717ntEI3ipa
0RNqN1+3CrKpEr2kPVYsE2SthQQdGKJgq6FfCyJt+bCPmY5cL2JEuDRbqWRo
ox88SI8CGcdbHj96XyYSMX7WgtdvCFD7KW38Avor4bDYBdvKBOo3wHa4OeZX
0fDlyPb1KUAjU+aAWGDUduqSuehQZJYVGM8idJ+CasEE5Nr0dsEY7ue09GIq
QIB+PtdmVxqx0o+cKWOEn7Q2ZsMhmGsg9HkHMqS4kENrKFy0CKjAG9dLf89S
maNUE7/HC0uJjVsaSglqZjOIyZx1z7PJ6h2UsTHt2VVJpJjYHEb+T/07+iPo
ZT5iOGkwcsRvy43WBbggOOetqpPpmf5VQ8htjlkO0yOrs+wJxl5i/FZhxYFO
reI/cEm7JjxQwEdPlb6vE5agFwdvBh3R5GpggDYtQtF5oB2Bpev9nWyj2Xtn
97k1TP5ZZsF0738vzDqkROtFJ3C2lF/J9gwIESgj7TIbzqUqcv+sFikBkLQb
VhEWbAHC1O03PyrdMVdUuHR8Oy2joiss7QeE9LxyOIcPgjuFy5ut8a+Gho8/
nd++kj92WRKzCK+KmXHIGL2DPuOlR8DdyuFX7nsjS8wYBnKquRWgNnXaDDgZ
zUOVM5IeLixvt6sVrA/gywpQcU81RE0MTS10lF7LcYu8ge8JtgA0qlOxwcAU
J4Bl9FdkVfpWdaGbUTyWy/eWu2Wr8BVeGsqkhk0Ifk3/hYwFVbavzRqYb9yj
2HS2vnwQi/c7xe/VWDM8IhncnNNUN47St6j/DcH8xwK9tFwi1p8VX3ncPiSQ
NRO7mh8T4eDs/Dj0dlezHWQ9Dxx2UeRn8jXyChWOJbPVFaPbsu2M0lYsRW0g
gI7IW/+ePncs48DBMU7PdP3Ym8SOOG+rWUuUbohaK7JEdtxmRgfZA5VBHZX0
mEg/GFnguzl6f0pPu6+lpdxDkN8uTU3g5tj5AL2YDkjDM3Vmh1RSuR3Q2iyw
YbcVQpm8qRR5alK1FuUd05Zxf460ezhOq23KeBC3aDYhTKuCd9GMbMaUpabj
sUfGxSeQg4emwRLYWsQt2woP8NB+AUnjEp+/H8sMCcQZ0wxTKoqIbjrLtkcX
kccq0OB3B+HcZi0MXorHhTmmkkAe5YU5rUycxdhRI6j05jQ4RJy2kD8MxzIL
fUHx7OaeqUErLccNMu1bKUB7qYfVV6dtaf/b5mADfL8Ml0oyVkPVoUP06xc8
yLJ0jcMsxg88m5tWL/8aSaMX90eu9+jTnmElFV+n2H7e+ArKg4+rz3ZIs5p2
TdRjQiEdwSjr8cOwRzraFOiDYIjtXzuMRnXgvwyWfD9bJF90UyBJLhWxs2G5
WrNs86F+5M/1X8IH/+Usv3BvcyZfXcRmj7/3jMfwJNjFkuU7v1Heole4G5Hs
6o0TNGdX2ZardUg99APTz84IKsSlts6ElcAdS9EyGoDaU+KxLWAXpnvOJm3t
h22T9wEU07n6sihXG7hrLiHF09atxe/arWFWCAJ2Q3+dWiCfQZ8ICVqny/uz
aDdUTMkHrxKWPEXteVOuD+ju9AR9sCs/sQeN0cjMcw2ugNTd9qlIl1xca4X7
5TdYn9BrzgPNZPrXNOOrk9F/Ltl3pL97t0/sy+NYJueyjIbOcUhHMa2D9AW+
TcAF2As+QbmKora6+wKmUdV2V8YeFH2ZRF5/1KwXdCwYUX1/fD2t9shJbvmp
CLbP8i+fSL/sxZJpAfZpzsgXs25bVWV6giLakNCxDb3Jz8AnHaMch+jjCUjb
O50z66BPGjydBmCWx6XnAPD504skE4POMiK3rImRJmWhEYkqPGr59pcbZkE=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzeHNP0oF4pX8a0FcZUpjQe+i11HDIps2MH2lpQwSUko+SGEoOQ9xFzwgUXL1HCQVSqW1WZZpQDhkng/MemBuSp00xTvB0/lBI4/7guCJCDojfXUWZU9m85xwztCdxoKMjHUafTRWHdiSCCB+tgm5nQb0WYqrHC1AGOt44CJHUFBtk2532noqWx88Mm5FR3mPSf0ZrMDZ3emgHZZZpg/JUK01uRT/u9D5cQFwduo55IwkTRXxpZpDx4Tw6Xj0K7gnUgA1/Jwe2qBV1UFaujhu0DaMnhMBoN15PELkY326KUT5k6OlmdzRDJ9YOY9+Bxz4ktyCkg8rzKoJIvwQCLnzbZlfKB7K8yNWopdaeyFSSJlMlbF330gvAhktsvUeOIGxiFEof9Oyn8SCmXGnVEocuJ/38DMk6quDOZW/91XYXfAiacaGT3gLhExWjsJavxkrG1QNjBx7mdhj94eoMXeMEJfCt6LeDwh4VFhzaJvZxFLzCjYnLuNNRhvU0bdWtWvJoQOIiN9hAR13qx8lSnTF7933tk1Si0pa5IXu+TmEX29GESCRommSNN6vywsolqU88VGoI5WkBYhsOi6MumlwyfvXNnmlVTyAVWF14lKdqekQG59iMbBmp/YYKOFLMHsFex6LSoWm9HVUijnIXYd3t4wOHuTtdG0xSlhDg2BYQpnfFKTNhPRmChQTPiu4LUyRtes2OI05BAg3W+w9kblEdZa62eXsn7/wnNxKnBRR4+y+RFsFg6j0rP8ao2hmikgbCpo1CbOiTj7qrqpteY8FzfO"
`endif