// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Q1O76VIac2G0xW/djzHobCS6p+VA+XvgBojj6pbCMJNdU8swTd6NN5XfBd7L
tgzOviJwYctoyloayCncWEFE5p+ImjanYWQh4ggFhyCcX3deiMdsqUogtzUQ
1yhckf1R5MCg87tm0D6sIdBdz8Awzkre57OToVjGt5UBz48Bl6nmCIVfmrSh
Bu7KsXnsw6nqV8VaOhPCbf1sZKL+3Irgj4SFEpu7t6kSSaZ+CLq8SnvFIZsg
M/YHhQ0le5AunY5HnIb4CzhSjQ5IQiJD78ZZAg0ng8LdTwVsQRUg1hvrd42m
Xnp0YvxNBC8wWQDN7SynHZQuV7JR/URRq45CeAY5Wg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Jl9Z8QQzy5cc2WmjEmwJzb8A+VP6CbowgFXHl3sUJ6F1zwM5Y1yYgB8PGw+y
e+n2E+FoQMxirSAWBM+69HfquzWu4xJC1gwcL3ca6nl1QWSuZ7oZg335EVz1
p672Tyq0XCnavnkY/pjF/+7UuvyBhkbV7A6eRNIua9aJSRZtkWAV7PZduw3c
wt1rd13y/Y/Q9wf99SKyuJDstKLSz2SwzZ8yIIfQU77okp2hHaOJnEnThIpD
iXcLS6Z/QP2w+sWumsLoQ32TKAIAwN4EHxeQKm8xmqgGL5vfEnlQ9dmSNq8x
I5fJ//YBKHMYSYt0nfGRbEIEG0Mw+6jfOZEHhjn6eA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vXPORQYlkYib2AcbFfkyYIKbFmwvgC8yBVeTR1gxoXemoYUJgVVHizL6szGK
TADqd69rFZRIXbQjsXI9RZy40OGysH+oVMBYNykQfCVmWngZDiPMYwU/jCww
cu3XgC9RMgxi4vhl3m8boEXPizZKIMRiOn3dsUTZb+Q2bs04TEG0qT2KjoPi
AUa1/ZWjKhRJnYGlMi0cMvB5x4oCi8airTc6hoDklaMQNmYuHfhk1B/IeIAF
5Ifghy7RiVHrVb3JbIbD3cdhoGNkqA7dVq8zBlXk0GTntcFItdRHZ+xURF/F
Z3GchNQdMYuPove/bkZr5odnJDZYbTyvWTE6bM4yGg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ctkhceUJR2KcaJSU/5wjD0ncbCotKfeq4epYa+FkgVB85gERbfXYO/tLmTNL
qVtjZyoFsb0f+yU9XUoR0lH0CcGv4zWwlWOe8tOs02DXNp/Z/cbEsQNgbUgN
abv8a48w/Jkln26W3D6dwL8B3xpgX2D6khULEBEDIMF774DyeOCajW/F/0Wc
BWYhKh0gD042DHI0ch5HkWgKHKMuPf5ohQEvbl9oN/0jt3ii3cD4vsdzuKu1
lDL7n+Tqz2yZBWm8QUv0X7P9NwEe4wfjasl5LEVMO+jFVEERUvzgfyE7Ezak
3nIa7oOi/EZVCPkKCkOAxXelEK5FT+aPueHveID/jQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
i8iOvqJftf4pCwjplv5wktpBzrJpv8H4IfTuynMPra0lnjqEtLHxwqf1zhwm
L0WJ63CvgqJ50K9c2g73Snqzpvk/MvgmSwIsgxMBKbruiZUfWv3hnXZsk3qs
JyREbRAQveJ8fJsWzjbScbPUXUc+IwPGBtC2TcVosB5fMMLOYXg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Y+tB3BaiG3vwgpwiqom8Diik9P9WTmaEhsRf5EbYtrxtWzmqZ0sJ5cnxQES9
r8zZBTzHn0xnd/EXITma0XlTNrUAJYdBWurFjWSad/vhzzG2+1NrPW8uYIgU
jQHBKmLzNCS+WTzO8KC85WBAOCnaA/AZxWzyA9ZA45P7aFcr781r5BqeTP/+
JzTvDG36aOPGgIsY2iOFsY10UYMAD8fyJ546e6Sz8VUsGwo7rdMJZJ4s11HN
OSMPn2bcxrOuDb6Z+FMG/7eInXGYkmjMK39dt/pBTDP7gRO1h/RQ8xoVIhVU
355khhfQPoXb/awX49RY7c19z5ImnWYEfAfeHQvvo1I1Op2l9hK9gceM1cZx
TytbJwBaCS5VtPoal5QcUzw8Ed7l2TGa2LPvOTkvAczs3LS4xqMloOpIox+U
6LUrEsmy13c6sqaM7KXAJmHJ0K3iA7lHxr7zrYKiwF65gvZ6Vs/1qLKtjtZp
ZBLgMcBa3Aa0b+KT/1g0n5mlx/Zq+mQU


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
W6SJc3i+UrF/Jyv3vPcqxoboplGYEoZuQXoc06ly61DMw1tAbXx+jXXFmeRX
UBz6zAgE8TbWFQYW7VEb0w3WK3JQFUt9zgBhBtylT/HoaLhCfIKBhoNn5kXH
SWtqDjNfPWvtUI0sDvGR55289yvuMm34yyopPq2yvVO6J91IpUw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YwU+9xbUqDpIqiqqahT5TVIMTJkCc2UNTQbjynbJjTOLbgC83Za0hjSvyIt5
6T8gbNG/1AyUuLBhf+IJQpJOaMIJaX3R4hDWzaYXsDBzI1A8TQLSIYz0PEVI
I1++7E0jU9GeIZTr2A7hmUcYXxuIxhWY4aecTjEZf5nVdknDtf8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1472)
`pragma protect data_block
2CewEEuFk9fvh77lfwe336zm4olPkwtX6Rxrmry7PUD8/Gk/1XzaD3l9OSYm
wLRNISMzqPuE+ng75hg0vTCTEUrb6lfKFhc8/5BZZ6cvMNKbfXNvusf4s45T
RaBY420NzT7Kp4nwfTfzDm3AC/8lv91gsblnHaVUulIULU8MNOl9W+46TQ15
B9V+RWu2eakgzZ0Zf1TdK8Ow7XeBo8elxfZo+NMqS4vj5/2tRM0btyN0On83
QUxv0vc+AlItKi+EP6UQ2R/THDLJd9zct3E7r88JKfh2B6iQ+8rj/WoJhH67
oucVZiajRtIBtilWUoFcCUp8rVRqIpfI7R3pBCQXG848ilVbYjSPoaTxIaiZ
01OBMymeq8mixyPuo4Es6BBeUPs0QD+Ujy5jPHx9qwvs9Q+v7bJb2OK3tENX
593FNWBmxNWA6g21vUNBXFzL+WpppY3K66Ezzr6FX0o8l6iwAwt71hzJnvt4
colgU05IdaPxpx4NTsnnDzbUWgNGYMnQIKKhIVqZlUqCVg3aEI4eN8PHAXyk
d/eiPNzQ4glt4cUjZM/+DFhf3ZooiOY32hLBpk9IQnOCG5cfsX/7d5pWJR+S
vPr4/IdogU2PvPc5o77ZKtzrb/uPYvOLo6k459jr++lbL2SRmasg7tQRiAMw
yY5y6uE3CFDjnE6VhSebBTHpisXvs7wlOf5sf0LB9DtGtnV1CocUg0p22odV
Sx2airPviIu6V6SPvS7D2ghJj5WzMGpMJo4jii4Mwg1lLGqyamMtnz/Bt8Vx
Lqy3oqpJ+O7tfa3ByQwLMmlgWw0PEOxUsMDOhSQQPf95DxJm6+5iLo/5L57v
6UsB6TEfQ53DX96aOZJBiE7l2V+kBnwOyqtqkm7JuZRPsp3yXgZ7F+xwf/U+
Bj79A63xfiU3imTaHnDxMU4rYgdDVaAXjPwqMjgBhauuYCfh7qEQOJNle2Ya
6mRU46T4+li9DtYGpCheMJVeGaVwZ8gi1cfCEA7am/KcHz/LPtSZJyCt2GuT
V0t7f6cUACpD2N6bZkFNegZkY9FLMqSOyfRmJufOcwB7ob/a6lzfkSg4GZcP
rzr7zemgHuHelTQXgTKhtkiIukGDLi9MANo/KUvlPo/ADmVduBInm0mfFKGA
yRTl441WhM2VwcwVOhiJg+HwhGSCGAXtMgImsZm7xHut6FLRruADC2RQ155v
zXV9SEMvH5h9P6nx74EPzb15hu4hUz79DZ3MNWJFSzvgn69vDVQuKjQwNu+M
g6VO98NidGEorp+iygFwtcktQsAW3h4sulfstepW8cyTuZtZBVOZy0n7drMy
cFfQMNsFKDOcnb2TgV6lSt2fxp2CFTcJf/o3TYRnLAuq41Q02/PpjvpEi9vp
r2ud9/1ECoA2iOHJhuPQKGPnTHgZOfU+WTIw1Z3TBXRxHIPjemNtcaJ8bCpz
Ug3ldeCD+UB3Gm/FGBh4ipeLVAkN92i96faxnAGiFUWZsuGHGJJ+POeW5WYd
iYXH6/2YujX/2kqqsYC3lhn9jSpK2XwmnXGncne98nWxltfATv+LeS51n8s8
xMNa9lEDPCAZ/zEqzoqglEkME1k9EeDbS797PRtKl+LzZki+tmT99rKa42Ry
FQrEnSILL37jlrwsqdR5/dtdNx1FU/aOCGNM/exAS8QHrscio71Nw2dKD7RU
hnzI3BRO8avmnF4L4htQPDC/DRRt+OKaAdf5ufifMdXt6uBURxnE4jAcaJgO
iyi3RkFDIjyBkki5nQyd5XSaUqMD0odcvKSrvDxb1xeQLNpQlMK2spohFrz8
bl1jSOfyUk/84RYd606XWcZycpvwu7kwYZfTx8Cwmgh1cm9YaHN7TVO/4ToT
WVd28AHOEegzAXiHFtTjs6ZkFkCRSddhQ8k8xHt2HYTyRzaR05B+35v5xHUQ
lG20Ynmz/IBVoXf8DVFUw+YMDYuBTwgwtC4RehDHtkQ=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqfK9P/w2aE2Yf0Pl3XDocsnslrIcpQ3TzNwgsmMUIMnLS0ZzwIjTpZu0hqELrrRqQ7WgLoUxmYGFOfnhNSRBzUNd6gbDci2nYMT14oGoZUF0eY99ySpt3EJ9yeNlBhyYu0WelLD6LOmAyATE1s30tMeNkS56IpuxTmX4RsVqjzATXN9ksKo8xn+0xJZInssQvIRGk6ijZdqi5CkE2hUnqkHVwoOM2HUQzsigyOCByTcBkGzunSwwyHFBCtPFx86Hf5O5x5JSm/hY3WjiONgTvwpa+UhnQWQF/fVT2wKLaXHN6Xy6kAYxMnruGGObjAmQttuvsje+Od7xAgkE+MSodcJc0FFrL8ps8eKRwpSpEzVx3Ltn1vXhvMGQ/rrXBpPhWryP2RXnFQLXvLzK4Wa3VOdo08G7rH4+i0zaQdfEYORB2Pz43wplpgsSsShqvl5rs1m0NXrV+fW5vo8zqsRx3AX02vD65D05zWBye0wy1tI0Oqc5eM1gbo6azW0joQOLJB4Jd3CnzTvsI+y3DIf64ATHzcnoW9mXduUdCGkZUmlYWFntOuaFxzA+gfR+AOVYnm+2YXpKeqAAy5Q7YUv9Kpb+4T2ymOFln0kfOIrnOTK9uiZtY6VTB8tj5DkGhwPRuE3HYZPlNo74crp/z9jIA1tS14ZhspUIJ3YgWRxPcFknhBphjx8P9Pub8U193ybMQ6+ukYhJcVR5EytQWnfRubcP1cWBUTa9JrWmM8rBdBR18X8WmG7ENCnjh+/UO8zNgYDgglFWs4GgPrp6Wcsjknt"
`endif