// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
h+19EEp5O1SewenvBeWTpmPvm0EB128MjjEjz5ALlfLqMyLtFOqU8Nw4QfvQ
X5OjU9YscFe2yrLON/X4mTNfLxCfdc3gurXGP+soaKzzDMwkk2TByXdgzCW5
gpeS1rtYk/9ZOOfyu+/hXsGIuUnYWo7Vhfs4FcidqZJch7FJ/uXACOQXm2vQ
gt97b1zSkLDSdgHwEmpanZ2+z339ARNmuwWZKFcSUM6DP4hJowFtiCKzaRFe
X9vlBws0meZDoEnHf6ygftihpaHpznvB6tKGnvIm9nmp31nxDcZ76n7aiCKA
XiNDlRV90j92RGMzZBNDRrIm4gZO69nFV1xVimcnlA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kR3KdKCRgZhDvBSvAQP6Ss46XW3dV49XL7Ge/O1mtlByL8ksnwfM+sEfSwr0
xnUWIFreYF5yyrWyNx6auMLk5umFiYbIgZTP/ad/rEkpSoW6xXA/9bbEQQE1
IQq/zmvJVJsY3nJGmKj1VcbPp+SgZ0hRaX+l/baM2tc9oroh7WTDRqffIOIH
2IzmLBbUuf2h8P15L1lxJolc6tgkRfITIwE0s8pIMcvAyuGexHI8AwVqRn2y
bCw8B0Rj4n/pemXG1nGmCO/Hv13NasypHi3fUeo/Dqe0QRtUBwAE8pcr7622
Bim8zMzoWECHuwsSv58zmCJHTNJrG5/NsYfzaCzZlQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
P1yc/RtlHz7HqXdwnVNuZ7Dp9ei7vXRjTP0DmF3az9IUhAL57Bfr6FyIy8/O
tgcBs2GQYqptpoPk0HWOok4idzmjBYEacu5YOtWsQR7sclnFqeDBvOGCaTCk
iJGPtUZp7NXTjhHxS82O463FIsyOsjz9dPKWQXTaXEfkdI7n2fa1axAj5LLQ
NLhx07cq55rf7yHmUvU5CrQmRXuef4yJ9/B7ggRxBJwYVHBkvr9Xi2cu5QVF
p1bqGCSoGLWDqYYhOBnCADWZ+ywIQ5akuxQd/iq3t5HI8Y3gWDCQfM1+SzNy
UWLdovrtDqaPJYS87ZWRHsynL7RcY9+/Wt1WmjxgAw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qYYo2pYIFDedbm8y51LoStiyWzQupdPEP+e418LJo2cDYHhOwG7y/V8rdgmd
euo6GWA16HXaND2uC8zloN6wtbuRzxS230/XUrq3d6AW+4NRpa+zPZlyROCv
nTvFqO9ES1VFYfRcpxth+2sqqNqB5vcbBtO/oRx2auvLIwVIullxT1rH8a6i
VEtXxXG+T+HG8mDLQNIBmmFSQNl1Kg/0WUmBTg1d04NBwy+Q2BYsXjPNbmXa
1uZd7zjM66JKXY1VO0wPFyYug6K6uRXAStCfusKKBB/RTiwR3GygXO0+j7vH
5Ti7D1BGBKibYrqzLaxc3ppE7wZcC2o/2icxFXqFxA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
e+KaW2En8NwsHciA4iVOHPc7RyiILOkwpHiill94bzMTFaKORbTOEKew2Zv3
87fvjVAKK41b+PNbo2XEUSjhzXLs+PulrkTZLjq5yinopqpz75VCiabHquwv
1VbfSHMZx17vNSzM92tixrDpLQ0oXuvmqs1NJ+AQQJjujTkIbBw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
gAsk2VnOBl8ReydAMmkrqKDkQrJjdRBcc7DsTbMRRwQHh82m2yI/jdKShgju
C9VG/f2GzBJRWl8DquetURkcC1fY2AUI10hHA/VL0f8T4eOmIjwFWycstjGU
657JwE/5kA4dX6BxTfCUvdRs/REVHPS5Rz+e9UcK80F6kWjbNodCUgiYuz4s
EmIBoVOWPwv+RraCywJ76ovBevLZUU+qXVHPc9Wi0YptCtWGT1mdEDsFciZB
jSVwi0Dfkow8NHI3JPIt0TPep3pBvUbIF8e1Jn9qdvmpYxY++AgmDCcSnlJV
YLHbB3aJcPXUBxA+jIZoiJ3sydhJkktE8+KLrG5+qmpD/+UssQdcU19SfdqZ
y+YkqDFQ9SLqNNUarPjOfOkm4p6AAvZZ+06TvV544C7BkXzohqxr3yLbRV3P
X4dV3CILR+8PX4SCqlmXA3o6nf5k6PsJcCigC/mXxtDoeCQyUWHS5GVlOsQM
q1svQ1gfXC5SCw4Dl/PZBmoBf3S6sAEK


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OGI57TWkrVTRrPbJV/vqEyJdP+2cY/zfV727/lXv/akaSMCwDtzBmpXMTxdO
k5Hsogb0ETBS6r2pVyG/iRs5Knii/0svvd+liqF+K+1ZQRHN5kZhIki0yhDe
W2DNH/Dx2kjBO6STCtxaXioAa1rfHpwuiTDQleQjJ1QP+HLnCTE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
H1YvdTD4Qe1/eENJqPqfhfFLB68esxkuu3keebloyw6TSh2FsVmeXrWgdYhx
WlqFuJLwBIbDks5434Ao1+IQsnAM2ebBUxi+5+f4BvfNm+YaEaOnAB5qJ5aU
czOjh61vtPU7Du22CKVeV82cp42gelY1P21Gl/qCL3cuJFLh1Ik=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10288)
`pragma protect data_block
d4QM+FzBHDKZkFDnBSSHxmSxtQpSduI9un53VBMUUz2QTo/kcbLr3IqmFcDb
4cBSB0AL+l3FzgZBQy/82f/3E+DjJk7Zd3EqMDlEGd3tfpwv/04Lo4oso1Qa
dyHDiLs/cw/WVh9yAcUvRPRVjTnaCKz9xTdMfFsfviGiG+BQ+XhwC2lP1Ssp
lLmK/NKHHwIzB/jNyvK6BTi37fh9YVf0oTZ+WA8JKgJK7VCpMw4PuhPaJ8BP
49Ie+3NcwuPQ2+jsAOo9uNSHeWw5LlCNhA5upKwLQEzKehE9A36SWmxiDIy7
e3sbwcBBJFBr39ocFrj93wZv27ZHFrZonb1ae3gxDCwtovvT5SkMsCDqLYFI
4lGQ4R0vOPLABydog1ZXWvBf8MTtiqXOE1w2vAQs14kwY+QPfYL/MsLhlLR0
sWOBFmhejXDX1cVi4YYuG3yZ9k3qIJPj8A9Y00S8YLgrZT2KH0+vW2EVd3AL
S67ZyXoYx9D5NP6QqfrFZLEL2gQCHtc10L8z1DZB0KebovTCkxGN4X+xcsby
Bvr4vHqDt+cnIa/HkkGhPHxwQp7q79YW+sI5UpVmsxDhNUl1gqLLjoPAgIDn
ELP7F2hWqQqszb2l2GhT+c7DpoPHUSdcuOqebcP03f3fDl6pqoj0LoQ9r/vA
Qsbw3f8cpMxXB8rD3NP0GqVYBUXckCfn3kWIbf9vsdtcCtcce/r8nQQw1yml
VzNg2fNksjbmOsQPI4hAsEOa0QBYsSjQeVuV4pr4iAhxkZ8iugWrbyUUOkOM
X/9VGNvQ0zi+PgfSYG/ZKcHXCp2R/CwXZ5NSNJQhovdCaHCENoVLbSqqIpTs
Sq3iCryqBW7bK9dyI8XPqjM7eeKkKOGrzPWncQOah59z4QJCLnNZP8Wmem85
Y8LgfTH8u6wILZ6Y5uBznpv+/mGA9LaKWlE1zX7m/ngTWxQ3kqNt7KjqhXac
8QwV/nm9mpRGtoWhwQZoM+VFMPnkA/5xUcdowvXSx3akUnRkXctgPYelgOx2
pkbMrCc+Vr//trUfgzkvknzhu0bbNoGuL/DgZj5Im7u0Q4HH1wsjlDY8R/Cy
6ndyOUjYXSj08gVeGO6kjfGDVKQaXf6s36E5CFPVBH/ZsIZC0BSwsFYNDBwJ
IHqEyQ6gx+HzmOU1eCXY/k9MheKAlEAEIUmkio7mTNF39IcgYOtJCEJ6NwQu
dQvbhPDAbgIpH871rMZg490Z3olVR7dPJgZm8Gzbhw7XBH1cIs6uv76XHvUM
DECeyH4FHpSXMfEHLkT3og65XbthkV4wNV4KOi/Sl6KU+SZG0I3o2U8At6/v
9iDJv76f/RqJPxjII04EnejQSF2OW4XNkBApT3YTuPiwixhoWV6rxIiDWMk1
txBfcHiC3bCNN7m5tFsle/ZQZ+OZ2adNTi1bnXdwpw9Rfe389XAHuhOuInYO
NPAptyTzQBmDA3ZAB2ODsJszvNOl1fwZxwfOOTP0QkKbcRTmOqVjVQKMIjdf
SPgm89HRJo2u8Xl7PGyNycZTT9lCOaJBn3CfyXv63K6vhnz44tF19BgD6W1T
3vPFk0pVklnHK+C8gbTsM2m1MMOASjzUcFHt6TKqc1E3BPx3fv8Z5LXd/hLI
PNVbp/Hlwif6q7UYhXWwwaDUpZ1ArPuC/+ZdeJJCu/ZwwHOV4YxCW2cB8q1Q
QqqiRI/BERZP9L70RqkTuo4cOs9FOx6RlL8xUo7HP74it3l3sMk9HXfa5oIQ
FtDC+XffGWWikaIj586QWgqdx9/n/00GIZLe12q+z7vItAmiSVftR3z2zqWQ
K7zcoftVw8tqn89pSMSEe0glPAL1l1Nau3zuC+hxWbRvcHDhH3bE+Wa/t2QL
WO4s8jDtfmU9El5lQhr/QvC6P8WabkAv7+1rz80BI1AcUEBRXycU6BnyPUEK
feDP33Gz74UXRDl+CmKFv3GBePuNrYNi2NMPc7SmQx8Z49HzzTK2nx5SVahf
y2Wofcfw5/TVG9yolWnTJlajwI25gv9aaWWaDwCeQvqGAs4wYJR2ch52Xwan
4v42GVK1Sm8hVs9D05cundCeSdl8Tm7sQivqDaQuAXJWeySn0b6fJixS7rYs
7KicvTbdFEkjqlqnpLibw2CHLbLGaPyi6Xfb28Li5FV/U8vVDK+SwF3GNLJI
zhWOz1XIRdiwoZ4P/QES9ZxLRnnQnlJloI6kdWSwgUGdqp+xwjM0YE41sIPU
dM2FKBS+ynbYnra9vuQCLc2RFI+IQCtmTkHhzK2Hjq+sw2GG2DriG1Zz6WLL
0fawM6QikT/QPGQ0RKJ8g7CcyEICvGoVcz281K9dXh5xugisjB8lbn++rwG6
pDzopqn8fH3aW0SiLVv9pALY9thOP5+iEl1jtl/Km0nUV/aWeKjm6sG7faBG
g52EMY3890UFsv2Hu1veRQZWsPeHbA7MhVnkHOYbHeqSOC1r9zczdX78hCI8
8vM228uj0L74p0/pJ4KNRUXEDPYFCiNTNoAq3bSvg05kPT/JZlXSdemHBpTn
OwPM0P02B0ZTvhLiIQVXX1jVLmWGP3t4QQm4p7SvbUkELC+7j04Jtq2FQC1Z
9pVBkcOz6SK2VFbMOWjLZ7WI7Ahd7HqpmJLORZ6DuBDAp9Vfqp3kdzQIk/Jv
EJpdzsV0EKixy2a/C6xBJVbnNEeuMOoF12/cYrJaeTCgOccXERQEqX13cr4/
OPCMku/3Ta3E3H9XlvRX027hgY1QdOD3BOh0MpspZ5AJJv+Nl7k+U9Z/tew0
WlavHLSdCPfb+dLzFhpSxDGv+1opP5DAIDmeTvRSxKSkKfru3+0GfqRBLXen
KwAgSsXb2EgLP0EKQN+6jdC99MPzEqa1estJYFy49gjq66vWFQtZTV94xTwG
aFFRF+Zm/+Nkn/7OEivE1agUexH40IsMZQX/RmmsRRQnvyatBYkwdQiBxBj+
+43MUovVuyXBbHta8R1G/QGqOIAqX/Bs+wqx6rJ0a7gkFxXlHpIiJORzH3kq
6hhyrEjgzsbo/l4zyVXAd493KpVjHAa8Wlq3xotUJ+9J3kwd/sYHHl8nQmcw
StokTqCYso7esqWjGczFThlyU0aXpksQY3Q8J3abc+vaHhQNOQp/hT+vQog7
7s0we4fJaB/kwp1n6WlPFeqoFUfHtIIWEWbn4u4xm5aZeeWhAfaIkIhEruk1
BZuu2Yj40btKUlbOd/ht34mA2m1YFEXdtl2RAo9Fr0GhdEk+51hBAQtZOjm0
a+uRbAUxLCr1SccQcG8sdMUqOB28G74wIix0iBkZuy5hp5thH4BrmiowmbkU
K8T6YNdRQbdRnN4gB9MzrK8tqeq8PKXpBCEqzXDaczNjiHbFL5cCAj8W1ljd
H+yGRt/YCwqza/HI/rwofZQRAAwNoKP7+6DouiFj33/XHbwQI2Cs/8J5vkO5
OADdWNPJdQn/3N4eta8srau43T5GHEF5rWzNzhmMgokKHxVxIJlgGV08kRNi
lgPvvDsW4AuiTQLiN27FMEX8pLBmX0mldTE8NeRRGwqfpMexJp8Kh1YyizDz
3543His90x6/vsz66zcMLZm8jbhQB0dl577Gbk+DWJzsGXNF8PEPwVGScRyD
GOjpZQfYZlqVYc0k2/4NgZQf+chCtpo+owXamhBUyD/JCP9lIspVg3MjfM9c
WxgYTdAlSxVCB1yTq6RODvVAgimznMlBDhCFS/y0zh3Y9mH7dNcwoHMo7hKF
Vz1TRxh4vWVy2BLCGZ0QUS33QHZCTOGJ0ZSWq8IaV4wgiQxa8OXlAr0E1xXy
SdldiCbKmTIXy0m779oLsZdCmEA0Tw8JwIhkmTeSu386ft+9yA1jU1Ky4bqH
jVTTf4UsPQxEd/w1ni/UpwBX8Z2XnNSsNItK+qsRL37FeFXyGBYvNRkCvqps
RzZrmyOvV/OFb6BUozUhaF1H/KnwOO8qG7i3s+pIg/JbPAv8WLM7P4Pv/o97
QbH9+OvLDwNvgbvwxYURVVzXGeTogWmLbb01J9pXNT13+Ck1qA1tnJO1I73O
xI22FLrexTnmAcv8w9r6SPtnsIBgLXvNcgNQneYOng63I/vHDYE7300I45Oh
K4nZKfPjzIUVpsBcB19/jMbc++kid/gCtYbumGSsib8VrIN8ztEch2xgSkNl
fvKayXLGoGIjmAVJZ7X5soaWTmtZ6GgHmvqpRn2gZlcPC+5g8pg2WM4bee/w
rKJVgzEhHsTVVvdUVQrM5Ligb67v2P1dQcOmtYNpbuhrlLG2UIkxPT7RaVEs
7J49B1oSo5lGc20ytBvQR6rnvyKdcKF5p5cxvQt92mztFo85gcfDCeKqcIM0
GBk8SfrFG4OXblHW8qJ+j0SHprFz2Pkb8TbRJ8DnDLA7dGC+f50AX+KH1gQ0
XjueMQlrYjJJRBZLQQqWhdeHR4dZBwcwWhhgEeiMdd45igcxhDCL/p5KmrQN
SEJzPbWG8JgG+Fo3WspzYy/jmv9KUCszz0ZfRvCJTIH9xXCC77P4BeaTs4FE
1xvChZ6/8aamVTRs3/dh6KPMQNMCaDDJK4wQvMj3/7rsUM3E7TFPUKHX+OVR
SSXwrtw1l0bb+YaeKdXZiNLxGPhq0rG19zBnYrg89A5DM3OecoOtoMriKiTk
788TGuSL9PivRcpHEYSXqCR9wXy9Y59hjm7mrfPccyjbc7jmhsL4g2lrbnaj
PzCFrR+nuT9dmDSSk3LJ/Xvo5ejdm4M6lQZaLyDnKy+V7AoQw8SWnLE8dt8d
oe8HJJe8csjm/FEoSsoBMTfiDeNwdwq4gNyTwF5WkQxdimMjJRF9s7TSiLQJ
E2ZKLkfBYNE3vU2bmYcsLkKzGswlJnx/wqaXbB4Xzd0oH1ykuQQWWlWgc8qi
MbCJg18zJMcqcg8aMBBCJCUTcTigK/JCXtpu8nU/hgILvk5kKzK0Z7uxQLEN
57uuyTAnh0chSfGHoOWSpt0IcW1xULZ2IjWnRhmReErkyO9HxCoN6rhxvTk9
oY+kca9CK1XZPiP+gQFo5dbp05Q9Z39WI6A61uCB3k/hch5WP1uL+e7McFtx
Pp62m8m66wkbb9su/Lo0+s72PWZBEXVYnTQSEzuA9TUgaOVBlyzviRQqwhfR
SUJTKL6iVFtXtSmsq8modEQzxBqLLMdf+fAXt7Bn/xiLWErd1Tx4Q6agdyk/
FxczjXFp0rRkcXynTRrxdGSMKHiJsZZamFs8zkrNr1ZaB8NYDlW8X2qk7iOb
QpF1JZPOTeL+9Z+dMgWCyknLkJqQEdBbDNmGUDPeEpUJ/2PUX2QLwH56yaex
aUPf3LwTci3TD+O+EOwD0tTSV/1HxUIx5eh6tsZB/ynqdw7k/giH2xPhDYnG
1kF3VW8y3YnIz7x0KzO4Zgnim3DXWBVcALvwrkTb1KGiHll4WR7rAlNAXkXu
R9DjC/2wztvmD7TflBTnHprZLhQWGy3KwhCofE1dgMLsYokvI/PrgfV2/6hQ
UxNC4EhL2MCEsWYXQLJetqPLyP4NGmrUPiB+Og3oC0bbStoCKnySynBQEJEQ
qgj8IVKVYjbWN3NVD0FRGmqVvtP/qfyjX+vW/ISZYu8ETICI6aLk7ZwWqTz7
6NfD53jyN2yz51jIGLq8c/Pxzr7pTbRiHFfPrpmD9VsKihv+7GuKv8Y0xEW8
Zw3OdGf4hCIHyUPvISYqoHSiU3rerAZIADQXdIta2j7TTLlecL+FZLB8TtkB
JhKmjUp55QPB6b+d5Y8EAj1ztrKN7L3PRqGpirzPuh08w/mE8OSxQP3Sjm46
IrcKmyZ/38jdwnyJZzV8cXklbFy+9JzhzquBAf7AIUR/gxgRC/3Ie6jNNdqM
UvJCUHpa/QG38+ObKRIEcoKlAkV57PRP+lCwqmjzFOM1Bs+srPMXFSoKULoJ
p7aa2N1X3Rf18VY0RgQlPl5/sI6AsjMMcZbCSkin0mq1d+U4ZRsY9exln+Tx
qcma7EV1M0D33tWdRgNVzdDHx8grVhVhakDlQ/wreHYPsgvz3ehVxMx+K5KB
eSGKMRb8FQ8iuEBNjnkWAZgdNyyg9yiWxUhWL08IjT48JoyLauUMRtF4i8lU
4RfxcV3ZywdWcVSJVXvlUez4SRuQ66yOsVFNTpJnSLndgPmoGPIaCnvcw/T5
B+H02eleCv9BZb2ERNmpx+TCYNi0QnLZbtRI3Y8U587t7+45r3wZ3rCldmra
QmDXLw5sjCY9cdil2IRV2k7z10Hj/GPKoB5IUaBkAfpH55B0uerUm2Iusoid
pjnI7sUDf47AozJU8nrnocbqVCfL4SJ0nDl7c3MUuKPXaK/oaiZEEeEXlhG1
7gy4Yc6fyWISiN/jYbP3RWnZLCbaMLH/caTnY/BMTA6g/lSaWzKA8Gm+6Xnw
STI573Mvu/DMHsctLwzC+2kSBuxhW6nqpDik65Iq9X38M5vKgPSF3t4Rcs5i
6Haj8hgCAMfejgLeReSLgg+wr79hShdrGvcVRDWZggltOyw/xH4bSIsKL6tc
nRGFUOOHmN2XCptUoL0oAWsI43doH+9Ilm0mi9K7M89oJemdA83Yo4KnzU9h
SAfQDSyB/Qn6/+mEsL4plLlYWZGiKIHbC6rAnB/fFs7QX62Kzrce4Bi2uuEw
rDR/SYYQw8dgu81zedm6oslGUT//96yVjGtaJ/FLrBzD+B2oHo+g4a2VeLZJ
B9DJgQt1xfkZqVznJk9tso0GIJNTpvoaYJ0g2MscJBBeb+HJDbeatuxbWc0d
m+3/hoOyo6aSv7Xcd6PPVgKuWtivDLCIRAueZWuXi/q32nnGsETgoe/gn7Pw
xp7HKzRfZFrEhNp13k3km4xul820HHHWV2QuluKIDcn0p8+kK6ktW0BwyvTI
ARXNpUmySGKUupELaOUFWrFaTRN9rSoPLDJi3g41N1L9CH361ogdp64sAfIJ
7NnQLKG9kC+lW02b+3LP3Kxf29v8jR43ijZurddBI8vSGFyONZbUAjBXGlL9
f/WCQRvjGG5r2LUb+RrYOJfColq8LVZ7fNZ97XEH9A6h+5xFlnqtUJXZmtCw
9HzCD7eZTApgW9hDHRY34YDFGPZuJI+hFexxZ6NsF1RDEqPBXjZCqTKK1M3c
PBdxnI7JiYp0feW2lLNCLXY4M7s8kgbUN6fahUQ98qri76u0YFysSGtRyY5D
GFgukTh0QljivMVxCZUnDZ4sRlCQKzfKJjaYkXacHazQDIKqltylM5CWL6EC
ThUeyOPd+dLrWCKVJ3SSuv0CVGLo2hTjU3Ds8xOkfvBnhYif46+FJdpaddmA
Ha0grL5GX20P0vb5FkSGCpxPkCj5hbl8M2D8RWqhv6wXFiOoIXnuDoemKUD5
auqURsJpgBang7Udm/ZousWgk1nLvBb7/ZNYhK6euNm/QAEjqRAbu15SlASE
1JR/MuEZAu4b3V+m1bJJJz2b3ajzar730QFCkYPRP+woGkPPr2iwq4u6+WRi
JWMwvG9qGzh1Wr+5F2hOs/vDsuWTevz8e/MFPlomUIK3baVlhB4Aqgb9WCdX
YMJrLK+MzRJdJiGDS6ia7YRdlO6uryTmzhm1DWIrPFaT71uSu1fVcCWruxR0
fB5puZfZfuqSLmCG/Ty9AuK9lKgflrvADZ3D4vyEyaOq1+LXutFx/BvWW96P
7bxW5oF92a29CIF2wqWqoKu7Ag0ox8ysECMcZC4K577yRAHIPLhkyvjlo68o
SiLbumQzyMhECjnOqe6gSqArDrQ2be4cZ/d4lrnedypsguMQ/372vV18D+O+
Tl2VzipHoxu2MUM2EE9WZ/MwN6i/g5cfl7ipJY14DgYTIsccM5qG4EETaQrc
XBvllkElIYR5+IxqkcFaobv9VCnDyae75W2niXS677DexCzDrEKmCScPWi3T
t0BosrUTQwU+1i31XvS7bjzrPTEHH2a4nuLZletbcGKURIFpYOBMRWNEuVEr
IizZgUgdl5wLxXImn1bMMz/4cEVrbCtDSPWb2dnkTNySZd4j/FaIkYl4w/BY
dKf3Gwk5Upu8Xl6k6+uwaDZvt0LF5C+Ijc75JS3Rc9zzE15iO/HUz5yqe/t9
Xq1HKefiGJggvX5Q3npLBI6P1e23WIeK8kAfKiMuDdXUfHiC7vVgPwV1uNpL
iAPyRmajH4/YznVEONkKMi2CVRcuG3EJx6yYe+oVXs5p28wSEwh+9/Fv2GU2
4cxS1WXIhPRmcHH3TkQJoglR8CrDKU5nTIuJZkOpIv4oNBnLUtfnFgNpsuNO
lo9lG2Et/ITdj6RTDLVHhlSCoOT/J9RVZR/M8DaEtWlaeu9deOiQ2ue7JWgW
BZh/O5PusbSh8j6nmQfekCoW+PRgF5RcYvh+oeUQ6aXZZRvYRczpBIwFy2oz
ddyC+SW6hbo92zY6dostm9p7lGsqOVzxN78Kz5vQJtQwomjQ2X7t8p5/3QvD
ZVM1a8VndLjY9Q+tQWbVxwkLjj5C4uWQZ+hne4dnmW1p55DNfG3Hc3H17/Cg
jGPdyK3ZKzDAvHrZg9Ea4X2I2nXbvai+G8XePiXguQmWb3hzujlwzC/N3yCP
sVBb5rCBxE/hy3lm3zIUvwIYEFHcNH6rGle2Yy3e2HijInzqPjoQzOO891P/
Ccg/JbcmtaIlqZ23zuWStHqzNOdnDMIwu3Jlg+G1AeRKk9IWXrbmumPOvjgJ
UqEI+GwkjDj5PJ0ZyIWyPDpbylNDwurA7yL4gbQxJeC54tZNYOEmifFDsSj0
XYWzkgL1s/3d3CH5YYpDF4iV/ZF+k5QjWMLsAeByyX3OeatZ7bLccu6K7i0O
xbCa7Vzn8p6LcyajQtEhCBCrs4ZSaU5+TfhUlpk0Kj3HkuZH5bbNHXjKHeSN
kdMRWyiOEz8k11DVCEgGlqiGIjwroSCW86wAy87XQxuOHimQUJyz/4TNWHKy
j6tJf59vYaZG6dhxTWb09T2INetsMqP6w8kAS7D9uEYj3PPJcFBXbAOM0fVR
zhKACDqGBHxs3cecwTZfeI1umfpTDJpktrW399sOVox01MoUl6KfiD3LaNB0
0JUJPGIO7ETIpkPxJegjx6WHVtZpr7AkLb3kkS57Bky0zycrsmx+jvjq3ACI
oU3mixTZFMwVo1/+ZcLjlDGsZIdj9U2HgZkiO4Wr67USbYPmZBJgI5H2+CAq
+QAI3feS1nSN4ABvhgcM+lw25MEj+wTHhlBs5qqVkv1UxZINSEtQrzpamrDc
oJZ2n6al6RNXDR22QqBzamcJVj/Uj6j43IscH05p1oxKiEITvA4CHQ7hrdBC
IvfiEbmWfrKIsjrAdpXOC74yyMagkZd8Ho67n2sjTAzdz+Kn45lLQfm4MlnB
+eOBl/UwdCp3ij90vC82gcJf1wwl3tQWtoF/X9Zmkt8uDwIgutTaQzij1xpu
dy3rVZXl4PQ7195aKLHxTrFgdZ/v/KAkooBs3cNVgPpOiWIYnahZx7bb8XKq
DRDhuB25BKNDeeU1q7ZJDCQNdvqRHJqJ0MNX/ahKT74kj7KayCxAjvUgwa4f
QPmn2ZNYB9uP4i4XrPITZrB6Up4+gMkmcCf1gHV+UIVSOLJ9VjBrKZiu+D/N
p7J6V6XZ1Szehj8Ra2JLGOd94+dIfc9Yv/FD4lU7uGe3/xTwXgeA8iaWHa2K
yv/NyTRL7yfMMN8gM29AmZMcJuC4zEJAYXAUw9k4FMdix3fI1gzqC53rjjAE
pWoJhoMZPOBpbMX0Ft6ADWo6YNrW2lYzfP4SMK0Yjou/sXblrG4+U5wjYHzz
WukE89sIu/7qDwne7Q8jtuFh647ra087WhD0pgz2M7Ygt0S6H7yOKeeUmlcO
19cF6ZM/G99mo22k6EpisTRYmDS0h1x8SY/WOi9ngEu6TW8e/Ek71VdhlHIC
wR8i8bkRznAQQOkfQdj25+h/pjLFUA2WPfdYHfgTg06JpYAHNoDau9WaKXgb
HCTCOTAhDIfESWPTynwF6Rx5pQGXQGgMFKV4dT2KPU7sl3FQ68MKTOuc/HLr
wggr/wGULA6Dirjv22m8175AQdM/56A0sjxLi5yB4UjXK8uDp1SGc6EIopCS
E6wP5Z7NjfrmSkyTRCuZO33HYuewXdcHeQxDTyC1HjtEQoSkDJoQzryBm9tm
vCINyo+RCKnnnV//gwg2JiyCeAht3q4JmXihSurU8tQKZopA0DLeaQBQC5V6
U9Luub/vyIHfGTSu69JOmTVlQEdat11xc4t/b1XuICcCbA0kJgsDi8uqhBBI
VdGcp8ceO5EAfbZUrTaCB3XqAyiBZyzIUZV5/DhZQDV+L+doHFLavmK0RpLl
Hb4jisMwAn6FD9TWtbisXVcqqGVaxMkRlUZ7co5KYSp3gcCw6bgrb7ZgZZVc
I5SIPBKLW/qVX4LK1vt6B/bcGRAp8/O4BLaN4U+RezvBgz38KtjHws56i9x0
kccAw4vLxKyBTCjH3THIqR4ZCH3odNuZ0STPtVXM527ErVhIJLXWaV9eHhEv
zq9ortdGxGiV4IbfwKIznj5yIIjJo1ue8kXxdrsamKNNJhrEgQj5SH1h0Okl
zB7bNhUi0WJX3lykYWSVkVWhnlbESnZHNko5ual9A3c9c9s8gcOSUdQmX0gt
bvs447MfA24T+YodIegW0poK0UY/dKqwk+KPMYYUtkldHga7BUBIAubPIbkp
YUe2PsBlr3VzV2FaT6D0ufQJyZuibn49QrLe2Aj4d8iGsIKe8ytT5e3D4ptc
uBouuKZR/UhC29DhTUJDhPiCkzpbKVIsamiqtCL6tDlZzSKb22MBkRB0StBi
kQ2Hj7eqRyc95gNNY6p1GsFD1y6lDR1GIiissBTADqmU9wK26UanQ/i7UK0F
m+gj6DRc4Tx8BPMFGpRCFJBpW1oFWAs95Q5OBJu0YvF9eKPtMqV8Nq+WCJHa
dhRAoRqYsrp1sIsvXMdSe3b3hnrtF3Hix2kdCvhu4VdyTuY8sbntNnrQHAnZ
3WTQJG6HYdrr5va1TlZNQo4PHtPTXI+sArGV9Tt7S8Vgc57C6+E/S0SEeD5C
WncqGtVWXduUtW5YmPaDCNX1D9pBHS/VN02gwAkwaQX5eKHXMnwAmPZMx7Qm
ysqRdknx135mzpx+uZUC5S+wp7rmd+3P7JM2bnKDBkJ58RtJlh0SWscAg/0q
JEQVd6cewgprfGEyVMoRs7lyS+i/RUVTrINoJ2AjmkPc3p5hK0Dj066QGEHf
MapE2h1qDOOmg81TCHpFeruDQAFvfthhygtW5j2SUZV1ieYaIuKxsOuOTG8A
MyOwJj2tRATqq+RRj4fDUND89Z+rZu/LsjMxN+dxbSGo843qqH/tk96irx5a
FCgRM08gX1G67CluGqxBCfz+iwZ0UZohWQHPcK8HVuEWhQ9r/IgICSX7N2QH
sANb10WE6QseaZhZ+Y6NjECLmDE1C/BMLH65DbmqvooMzT3vDjedu9CuvGnC
6qV/9ml2S75+ZzZhoR25P0uUKF3+n5oXm8tVu3iIucR+eEVPUBTC5HCrk4/x
OASFtJC+2rzrvJ3YEITO4qWfMaB9xYcVuzhORB3goPE2jCiAE5JA5TXPERTJ
DR/M93r7fsbYsyXeI+P3IpPV/qOoymWZoi3cQboo4F5+jyYyj2yP6rmZAK3V
er3qRJT9s7Kf3ioEYrcmIgxBoet7NF4NxRK67xYfym1YGlhiV/4UN6p7uCnm
E2MlqPD9nCdNgBMMLQYESg+AIVCP+wvPN1X9MNKzzDzzJQF2PBQQC5f/Kr3Q
BpELtn2QB3OqU6ER+mWkOBO1gOVYAa5hKjzfLRiDAG02WGvr/euXT7t7uGuH
G/VStNEgpom0DshSTOsh+NUw3QHpRwthWgX9vC3D/OkXEEr9QSl1xSAdzksy
uW7Bu1k6QRk9+gXM0xJhUHf4jMfn3b0hdHfIwt1AFeEwaXBj88nS2Pxtw4bz
DiZCZ9KRElDc7J06wWrRr4r+4q4eRW2No9XfKMFB09Xl7NKsKENH7BHPQFQq
um1/8daVN1K27Zm7Jf840Ck88IK2A7MMaPEiKfNl3Lc9uj9Gz0I+WYy9MZh/
2UaTUBZ2wktuhCgELLICqIjqvSExGSglSrJBU3HleziFqw8WmxvPyA+ClDCZ
GIfuQnM/NumKpcE5wOmwYVv2HW8YBxllBHg3FpiHNMZmj14vpZI66z5mpaUi
sB/lFsTOJBVuumZ5g+Y8XhKIWMk6Io5nTY3RDU/+b7jnW9ZOnWMptAZotA+0
rWy3MyHPhKgTL9yNLODqBDWKFXIsMw33Zj7tESgS7p9HEnw8tA5Lg0G+/WSE
c2w//Dt1euZcZojNg+VPXVErjfUoLdRqgeeLNYHZ9UJsCRclkX/7MYJgmID+
Iof2lkZSlhdlyDavJRXy3a98rTz9PY1h2zD6br0Jtfl5IlhrOwIzQwVY4F+z
g42DSas5m07Lb/ODh0mKr1cp+iVsoPNEGENypTP1OfH5WSFkT6nWwLQj6oRJ
e9Zj8ByJenfPAGftWTVQGGFyndPMPTio0HQbCRR0rCusdOOugynFZm8HC9FL
4CYqhUUPTpOQsAUeAUwg5RJk6uD00XdJEJBXw7MLNlXlwHp/UvsxhP3kdw8M
InktN5ZB3hrryAjmofjQDQPXwF6pYRe+R+2eqHlbD2I+rPzyagyPL8Do1VUc
o6bDx94VwYBWYRqJVdSmZAxx0cWRP3bapgRYehn5I2hUyuSjS3aJJ5awA6Lb
yQDqc+nTGD7irSVTSLXs1aGkXGCzDjG2O3yQ/XmIK3KK7kjyqQ/4ibpMNSvL
dzw2QdjFIIfBdgXRtei0MjVyTuG2p50FQnPoFRAfTRNbttV5BAQNoteUbwGr
YeLV62xSk2iSPUAA3f3Be0EATKRY9M0StSJkfnw+obCNd0YGUMpoE9T/jdOG
sqEplrZxzVztGnDS49xqN7+t8NZxLBE8pt2EMON4oUECcZaFctocsF2YdUhe
msCysSXtJzKQedgB0BJFEDHkHW8n7kLt403W/Z7kaixUC9A4SmGdv7sB8z4R
DAa/wM6RwazLRL6+eSzJqgXtnHlBhwKxOzKQ5zgI4//R7NSMKIe/3iO63Rmj
QeDiOZ32OrgBdlaZXE0byCDO0y8cu3oCl6iBZNmPJeIannFdbIYsAolbwOut
B7YfX7w7LLNPexxKx9ld3TFxnIhYwDSmqcTi+lZAVzWflVR9lgQ1vD+ln5Nl
RpeQDaQJM1qmZ24d23EmcXt2hgCJebq5DVk4iUJF2zvEkcXZgP1r64g6sjhR
j4UP9t3THIA8lVfNS5Wc1xrBFYSGcwk+juFynCgl5QqO4Iir8/Aeyk3vn3Pe
23DmhqXhAXk1RdzRALteoRz1jAtBwdxoDLRJ1CR504eTpUbIEDTN/ESdHFVJ
Pkb06V6Fk4vJ9+4mAh22cLliE+7nl4vuyrVBcc9ofFo6n/nKVajUg0IUd69M
nnvDNAeOeVwAVDHp0iAvrbJhvPMMFNMZOFxSbX/8I/brvEx1C8gGdiLCllVM
rvXteFkFOl/ovrVpPrrRXbDDooOyRKwXceoF8Ap6Oumrig1yIM/AMWXQEHmA
oyFmbiRu20E1lTbHTvIe0B1MFz6fY56TD0kjRv4WSFtnATcaJajz0NaLaXkZ
yqRrxMCksdHAdBQ6uu3XrEh5l2JiahnU4BeHf0P3fsm1QHxtt1XbQcfh9Z65
IyIEZVHZCUhdtwdfzn/RxuUIpiMpntRJSYl+nfBaAuKowkjGZTWxLx6y6f93
Eu3n/4X357BseWdoxEPXPOWk7f+wACjXFyteyQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "9RW93T28GeolckbYRvHffOsKFRFmORm+azyCUYhudrVC3P73ufaBfyRVMCXUVPfCA/gVx4qupGWo2/MTXHrbiqujt9kp6+gvryDIvlW8esKlSeDbKqIxzhLY+DL5yFAjg+mCmTKnMSoiZ9J0N0zgOO806IAkac+OYN9FbEIEFuaO+G41krhhxrcYAZ7qVX+m993ig0jH+TdTkf+bgk6VV++svRquWf4VNDUj099hz6DRTCemdUWnNXPjQwU0QqR1pjqzISlKQFSRF4VCooAeIet1PmjVmzCU/4EKBPOuQkh0pwOccPKrwF/EGJUZkHd87fza4OpaL8IH9rYB/dAXeX34XVSIhBn+qL7iLgtBee7SYW99BygVBqkaO1KqQSFUCytGpA7/qXArd7wO5jF6DKS7R5e2LFVEKqdQHa7FBk/3HzZzky8bPhjoteuMeDsLXVw4GOtVuspVWINrvuknXxilE0T0wmVbbtMQERSPZ2E3mA1bTtEsBmwpt8XJhvzBmx43sbcIPu3aV6lx84AXlX5E6Xo9ioJNAXtkulM/e0z52Z+Qm9pnzCm75TSFAF21I1hovlVRV+bM9s2/zEqlvJdZH/MCYNqhE3HxUN38+ov0Ba+P5e9qsU1BZsIn5UIQBh0bubmpHzvCLnRfR9XATWqzpfAyBCGlNkY2DxELS01yH9sUvyKyUrl3qvG6JV8h4iNb3hJ+/U6VuC6k6J9yUgZqym4bqLz74i233am3Pzq8OYNnEK76Xrf6UQOfR/nqVOPl/DkgrrxT99zj8V6QwOLFHQq59gNFkYHpQPF12cbDOiV/WquNexaOd/zAPEx61AQ0wirAEYpfGG5EIco0GZv2ieZ9rsbyhzmS/Mtww9xVsiZhe6z3gT0L6B14KKmPF2yvNTQD5m8KuhBUtWh8q9NjrMief6HDo3IxS49YdUmXqntf49J4lMepQUbl8AN+amElA4gyzX2hCA6SZ7Oltv4CpeFMjTssupYpqAyNqrp7KkgU4zqNo7cewSyEfApP"
`endif