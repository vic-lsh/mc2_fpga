// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DgoJ1rCwuzpM5cb9OtLatqOIrhW3Lb4Jm5lEfYE2CmFHn87Ik6USGRHpSaOy
A4jMp9a0CuOy5MRDqmrKeZyM2C9xPOk7VsuAE5lMdhBjin+iLF3GAny7jiBL
J5gWjxbJqZwnvli4SoDj54cvdlhGfm6xyxD3DHlFbniFj66LWUNljF40GnDj
LDmOUmDeKK9Beg7ljrV37giQiy6yqLlUIteqMD89J7mb2o6J4BWejp55jhy+
Kkb+m2N1ywyn+lxqlDebOc5UejqHiD7E0hLvdnlbMnOLooal1vk1pZ+NfCrT
Me8JmACcRcoM3RuuVwMS34+gl8X+RfUtgvdazDmZ7w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pfsTXeD6wDNEOZTPkakaBAPzdsMoCBAVMUq27eVSfqaGg+ow1pylf+tM4glF
FgwG8exSp7WXwY5Vu7iaQhcYeQu9oq3vGPcBrDzio0ZN0T6ubQ+Gfv6zUGfa
Zwlt5p4iTOd4ttkppmsxWEi42rhGJljitukyrp+exGGba2cb9uyILoppR0Pe
8DFWJRT4vGhfxbPyg8zNLyAax1UY6414FYb9S9IvVXBdntD6MNKvTTeo58o3
i9hsAM1uGZl0YaiXNfDyk9nhpXgC0wPr3StyhazI6F3GdN8yC3WBxKOR3psS
UBFFDAf9XnU+AAdg55mYjC6PvZ0KK2z647cjfUeAOQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Qfxy6TwNmqVvoqCX4D+NIk6sMJCe8+nVF6oR2LlQZ7X3ACQMYGyCExoWpov0
YjLl7BMfXvg6UujathaOLEUnWQM6pDiIW8NHZ9Che9PsANZtrB8zsCCVJEe4
WdnruBCU+lLbh+VKB2s3A5LY/fbZfG252dvsRWaTLFKV5tVg/Vj/1O8/t3hD
YnsH2wTGKBmzBwspQEJf72OfYTuHrNAAMg7jdaRxq2LHxLGAZKk7Dn86FQpt
7on/tUaiu0xK+0mlAo9Muj0xky5zMnpDb2EOgJGF99eSFlNyaJMlmS3nZoHw
/aK9TFpcwRC4VP6JgJ1C2TRpZ6/zHmSVxrWjCkrkFg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DmSJZtLur0UhqkpfkTS8cQQJCtK5fqKenw/Pw94FMJLlOOujw7qw0ACPBDJn
1K55TDTEtXRy07Ljb9phS9gXeJbNmPGXVUqkXK4dVX/OQB1134JtwZA2WDNQ
u4GZzxzPR1mdMfrPCyQsm/hJjKAHMGX1h3t3s3IgEyz7vlyGmzwctR0ozlLu
7XQU/mBIdpWBFJY+jGqk2FuoEs17fmHwqOSN8trE2U4U7qCrQCEmE+GRP9mS
cTSuJ9s3gyCQd3I3axQBmL2iel90wWFewhoa61DrjE+dkEpxXa+ABOVoG0Tn
pgmXPhes+zr+UNbtD/M8wHVw0LJ1oBtxhZSf/+0bAA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mVXtqLYb9JoCM4soUSjDYrzU7rJ0p9R7x3aiY8K/5MKuSxu6Cx8lKTz9RKD4
0mSIRKYLH5acIB6uWwOmy+0IN7jmJnJ1NKxVWTDIHE5W13CO5llTs/4B/iTN
Ng5ENT2Zh4j9yC9Z0RXieZ7rR78ZvPhl4T9qyqRNOy/wxcPdGC4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
KNrhP102xVqpx9EbF6UXfxlms82a7fMzi762kF4OeLdy9iECPCz9cNQI4V8X
43u/CXUaMBpaNyky25D+P0k/WyM3cKneg7oAOt3CfNpUtg+efeSuM2ipFnrC
SnybbM9iDl9meOQVIRKiUbgKeEEoFIva4+fGoQ6LaELYOItnLcS4yviE1IW6
3KSn1VRwyTnYk3KPQEGm+q1AV6fucFjAiU6qb4+7ZMQ+EdYVZ8MfGst2PsVZ
dxExPfwju33jLSJ7K4LsXGULXU9etCZ6mOjyKFV0xVdb7q7D0XLC2uaFZFyE
9DDKc4OHn+gda/zdjdp1s/FRty1OIfPeDvaT346vKywvcDlQPm4amMozTVss
KsJ8q6h+YunF5khQNejWKYyOVjy6U6Ms+JFYeqEq5YU+bA4quyhSCJBnGF+K
r77vPbu5mjwVQKZEqhualF9msDwmaAF5xjTzFv83xzCsTqGeJr2GxSdbAhDp
ktN10cYwIrtq0kTj45LwJLM+1SsFFwSX


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QON5+HGsyYMpncsp4A6buR7dTH8EYY+JdTYUsxqqYjpPHYSOJLGFZPEdecgU
TuzNNNvmylXQakXHWEICyvnSt+g21a6or48KBtmTpbfeX8Mg7CCI8CNv2PNn
G50K2NfIfUCFsJ5rpeavdDz8CGNu91DHP/b7pr4KNmgEUowODIg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TNX+jVXaKVpDAAOatszmDm8sb12AaVGFRrdppx7r0B68XShwiCrrYbNW0T0p
73QSW3whksrZ9Yz6ziLCBZJK8p9jgq7ZPlR3/EJISeaTXmkoTrYCNYEqlFSL
1DFBeK3b/nnIo8mAoxsuDR+wimxVRJbRXMck133Clp5ngMdqAfs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14704)
`pragma protect data_block
7Bcqi3erj8XHwuxTISaawqwgs7XGQ7tu2GfjgWItMaagdw+ce688Gyyy5JYm
S5yYfT7No5e6JgYMImO1XLt3QLSa9EmuAoxC9AUx8FeeqJgO2EGT9qnGC0US
k0GO7wvDnMGC/m+2lvPHxOgRV/e3WBXK/lFsISPtMRhzBa4RQM/5d2zV0fMH
+kWBXLfJTtsKkhEgcrCF7Uxhr/h1qg6VPbLuVbDosslLMsmxg8qhWhwKCvV5
CqUjPK6ih9AjDferNQZ2WDAlGG5ZZwnCUys/wyLfojIwjVOCD+WHZ9b+Rhgi
cyqN55ZT/wAiZz6EbzPhp40iJmfaMs379vL6LZEpEhZyL91pKPPFMGMO14YB
nVRpYjmpQmViFsJ6ejHQfPZngEUyvttok48kEgyWowoiBL2q300+l810ECF4
yHkDETVDVy6Jq6EPCK6LQSrKFu8dmwL3OJE1sMcSdN0Hfnb8LwIB9btKBEEl
pRihXx1Nd3ctReWpwjyEorh1ctLBjWv9fMn7TG8Afv9bPXYerwW3W/Fp/U1X
UlxJuYr7+cHYRZ8zQ3lWXP70hrd4KOPu2hV/7DQVSK+eUKg7eN35EjS2MqjR
QH3Cdd57RJSqPf9iyEA00ZFsn3MrbuoVJu6zfxd40QF/GAIedlZabo0W2zlc
5kuAg5HRRMyIOY+TqR8EZ/i9UiJsDoNHVNwUSVtLdHJrOB03atavgCnToTtL
KEZRs20mGNyBPUbOruvmXnjciBopkoqtH7Ui9uahMwr7mO0NtOSrtzkHu5ev
WtHQsED4oF+itLqT/4G8ZS2Tb+8DChKUWnZq+E/W8sPVcebxtR6ZwQITF1A1
0n8XHOUo8xf+A9AWSqIVXR/t4YpdkQBHurGWp7nOVQxgRDkWipIEs6BJwwEZ
nwp9CilbmY960asHJp+M4zLpK87P9HTKyDqJrbdNAZ8ZiI05v+Og5RlZcknd
lQm/n5PcJE93ZFO7kb5HU8g1TfQYZHk2WIMnZ2nLcErF8rZ2y4eaccQeLFi9
rmHfppR90/6OmoNY6M7niqAxSQWpvUIU2M1v9d5oB3uIJIr8MBhiTP0xPNFu
pWTXYkyklionCEuOcWksM14uZvyVkQvNN7qgt3EVwDHTlNdkmE10ND8kI714
Uv1GkXGOUdM9KXIFCqkmUfUy0lArWUExOZLK5OaoNr9/p+10tSfOpqUcmu6q
6mlzSknhxocL6IAbUa182q4ZZ9keOg15c85UXb0NsxCTXdRU/nNM0ENfe5Dc
sa22c+WfqzUjX5Z32EVe4TFCiwU90Z/rKgdTCdajrtrMJXVtUhYOvC/0ywPF
ezgSFMQZxVLA9b0QvCaV+fbB5EEfWj7VsXZgYRw/CoVm3Q8+y+WCyOMyXkIM
Uff82wi7Pb4GYSTjTNToILUQY5TtUWwauiJynvFFHkBJONK5esCwV/wgTbc0
ln+IArA8inSvuXaga4cUGFKuYJvQRkSfZpnaw+yCGc5b7fmzQm+5VpRV2OiX
VbOLF2AJzTsNGH6Jnfzxrfu1saFsuQUwGQBDyZGN7LbqGxWXEQPSElXWKXck
Newk5YQNRT0F4eGpCPSSd9cNrrE8Qj3WJQNQM3YF4xAtUrtms+j0gvNapki3
L4Orj/3fSm1gtbEm7U/TXGgbt0f2bcvuWGhm89b/85mod1g/aABwjHXGDd1E
snnl2F8kpoe3PCRF2pJxnNXWvd1ub0AG3hAWlu2jgaZOIWMm32jBCF5SPbGe
zCv7hVbgc3B6psetaeCgmKVm3gr+3/tSk2SOT/MLVoswEM8c0QKxia1aBvQP
pU8qqTURwfBvSghLtsvHC3IFTJrXVw3jiP5PnkR0eX0Op8jOjZhnX0k8u9Qq
eD18qGeAAFj5WXGBejZvr18SIiNtrhqTCunYjvdq1VPGz/QtECd6/gRuHTMX
id801b6dx05+YieKkjCJVkZq/4VpniFu9d1V19MgqpU1n86P6Sx4iFu4Ri+l
I2MfeV3PE97GBupX0oAtryZQmKh099EBDDxdeVb1prOzCAtXooqrgDSy9JqO
aCZHYV6sk7ouDX56nxQXey8fW+5vZePP9qmGLpnQAIx0yX0ClxqfD0TGhPu5
SCBia2D/ICbRwU5iFsRu2NBPNUtunwWGq8ALW2hvYdK+Lx4SUb8mugJDGBaB
alb6ed3GOsS4uPVljSEe5IFbiCDTYikSSrdCLi2mC85ZRF8IJhy4TglMf0QB
wUrNK56uCZvA/tfeRExHB55KwyT2q6Cg5eVIFoHhNgnzIIAm7zSJ5kvj8ERq
zZ+rd8JZG7DRpQPc2zz886Il3ququd7y7AbTG3XG4GEslniCQu8owwytjMUO
6UEpGiBBzrnflZlpgehee/Yy7eT97G1ADOwhOhYhyu0+lW086nau3kQR/lHc
jwha/4qlw6o6zG6PKfstNUm+owYPtHfpWUmfGrj4uMFiZ3KjZbAAk9hCwKzN
V9XPagxRT5+6TiRJ/yZYEuxejHIioLzgiaD7GDjFP/31Gq0DTr2IpbjMSkQO
Ok7et53ZzwocBDlNWqZYBeE3F193Gs22kz/U6d+TkKAjMazwUnIT7/nU+iRI
2KAzTDH6INYg1Ad9ivsp7VmSBetLUOGqVUgoBd7mwZYqYFXk7wJaB94Kl9eU
qYBPkGzCzFQfY5CjWJdJhgmW0Qup1SiJiA1TML4D7OxRlYtkmxBwLUDLGak9
mfxR9hm7sfT0NuA/Z5uSyiEXKdHkim7ISRsE0WL2ph8Q/p4uv6riu0gCEvxI
ASE9jciICmVfLQyNB04jeMi82YB22uDu39q4T8ymQf35F4f0ENT0GOOlpjEr
NZJp3IpKp2qfrTmXaJacOzADJXct00a7L38QdQ6dhlO8vTRI3FJjOD5f6wET
ufE97XtKQP7n8qXG4j3hssrvXI9Je/IrrLRJ56o60mXSUKUNhTq5BeXzpd6s
8563CVKXhmaxIUveMqNZ8TJYnIyM/YfQ3W5IfxHaS4n/bxe8M7u/ekQzLyBK
t2Imp4cfWWgpjfvWwy7SsF7CI7olsNbzSeYGSdtaMgs3FuPWxhIYzTuz1BW3
lr1eWdtYTePLkNKJMziB8W8KwLL/P+gJIVnrgVw4H03ssSU7vmuyB05EJCsK
LIm5q7rA1K8LUWhghfOe/mcAdwmDhMemhVXb/gcnmZY5zXBwqyV+71Y+u1KX
Fl9ge0thV9Vr4wtvr6AfIUP25jEQQ9VkyHy2t+GgjlnH+aJjjGEfgkXA/K/8
zCKQrS8qla6C5EYM6REq+7pO+krFP3kL1U9ih2fEnGdyq0riir3nOwFKQ/Aj
SDaWSeIv1iBmjCC+lhEFwfcZSgFd4aFcFenxBUdHWL6h45Hp/IOewLvjGEl2
UNhXk4/L3EjB2ltGIEFhjEn9hzk0YjSZTVTSX2WkyGgQK82QftFJep45IH18
No5QfFhhe+Ucp+7bJwTC7Xrp6R9bPSZ6K9w644TdqXtw7xOrFdftG+BXhrTi
0ILHdS0Kf+2/sPSk5sevPzcfSsVdXP3hbumLKaB+zQC7QMonU8EW0VIK9AQ8
7kEVTZYLIyujmrmr5UuivcKYLI7Cp2hhcljVpRGNU0C7bp6ZRVUKUYmh96kp
mOeONVTzBkp/JsXnKUYNtBEh7km/x/IOD+mJkrcA6w0Vpr1IQ+zNeDf01ePe
3Ij3FPPaX9OgbDgUSsZfHSa4hKYWaipzr6CtqyNAjqhsO55SCIzYlYDbE9Oe
CnWHQYnC/LHVBooD5CG+Bw1X+ipRW3kXi75EgqbmqjBcF0EHzGW/+BX8VWEv
hjkvry7oy5n4s8beZwBYo79xUou106VTTNlmcFnGB0BrWoeyg754y4hoHip9
wkD4Bip4qoY75fAV9jeX4VygOg2Dw2YDblmK7yIVmHtljaCkeY909mexYXi8
WL0OzKryDHfsEry42EHLc4hNGdtldKVMeEOOjG16SUT4hgZR9sqQSNk92RyG
h0fi22ZWO4KIpZknAD+7KMn2aK+8X1ChQtGy0+8ZibUx1jHk/PFlA8Rw6PP7
+4/hRtWD31J08TJFyTn2eHlj12WtwUxwZfdbPBF1AZZvzFUDEbxDQDfQW40S
UJn8AVRp98/uHRumghCrvmDS6kU3JkcY432q6oou4G4JkhpmB35ha1MS8CJa
ycVBVV5/YGnjvgWe8wkWie2RWLMVa1wmu+hbbEzHb/LnOStIqrjG/4TdbSuk
Jeeu0oMbMfXyEKXG1d/OmszZQIXvAIhHiUgbJ8kr9NeLQg0qtA+YEp93SYFB
OZc4OnkMG8//S+roRoCotmYCHSs0scoXT9vHjFpQQlcNNLzwi9P/AuzB2iMS
+SIniTCcyiktpQ33uKooHoeVfI3VVra9hOaF5FjZeeFYwKVhwLjV0xhMgdt/
8Jsghso2g9T2MF2psLMRDn2c/X/1339jZt/O8egIU/OfOZLBp/5DPtkLQgfj
S4aYRgDClCpFiR2oGeFjYBhV1m1MiBIzXXeqwOObC+lCLaNjrYFi0acWpQ+8
BuFnxAzJHU1ELtbg/DT5cjU+aC2QVKe3GW43/OXCW56OpWIHdvPGOzOtwPeq
HV3FVQUg82ZDmt6FoUK/Vf2n5y76LVlrW1VmOztJkcaGRY/2Alxa3NQ1LGIn
g5oMJRTIBB9JHH4EVljnb6U3UsWmiZWvWAND2Q2JTyfPUpdbrApVWOFymlTE
YbZz72O+GNKvA7K9f+4PD1X+IE/cMykaBdQyZr8jgg+alBU7kLu5pqFi/dyk
N78fG0HHyNPhELold+dE+++sXNlhG+hB9pdP0BLbSVlMCb9b3mJx142E4r/s
x1z53VCoXk/owTumCqMqnBbNiysrBksTWQ9AWC565DAsBe68WBzOetIpj7RL
sLPXK0Lbrep1DfuyFfzdIfA8o2G9fPagtnPXHIiabmGxbuDBm2ZFyz6YdcOd
teqcv8HjCwVbB1n7UE9dV+w7utZzILv2uGk3mEhJUQO4wLTnQ9tY9zz3/Rjo
J0QmYkxUBAKDnDxmVUxiw9nFOXb35R8BRj4RDc8ADwZe+DXp4r2YLSONQoet
/y4IkECYACSW/02g+1Qor8uahitJSvbeQJL5numoZ1t9FjAOj4YQ8DJztw2K
eZFVBVrGzpLobrwRzTwXlCYKgD10HTkXl9Lfwq/sz3TbkAdBVGvtMjplVDT1
KQz1CXk+EkZy+WgTS7I1P5QuR1g5KYLgISC8xsS/0N3xE8f99iNDlX2CCfjK
l8Ztfbfp2t+J/HGtZkdHcpapd4iEAvCpj2klKK7+NLjk0rFQ8qmuzVcFT5xN
3WUdHFJno4VRrKmwMbdb+dK1KlbQFVMffrl/b0SUT5zJI2MjsMWtL/Topi6F
mrMJFiwylS22aSB1MZcHKpt8NnAILCz5DSC+vrz+jbd58jWGqt1/L3ad0Lmu
ZP2xQ6sMqOCWwpIbR8YnMLF1S4UHB0FtLz4hE9RCJ0w6Sa2JyEzpc47vQnZA
QUlS1TRRKsOzPS4woDoAFWl7YwC+IWaVMyf5E0Qxjwf27B0PCtD/9z38V5Zt
v7UBS2z6miq2eBnGPzkWUxUh+dcXD/TbfrLla3QeWME1+oip6aGBPYhAUMYj
9wTBB8aYed8+FNRX+58lp9F+N5xiUx7P8HYlq1vB1tSY+j0Fn7Otl70Ssmv+
qfIoSzbKA2tQQBS+tFTQTKN5VRvJtTaxprZ2BvuYUvSEMLjllql9AXS4Fph0
AQEeONh37W7FPolpid4v1VSmJv8h79MQ1AfCt9D2F0V9MCgTetDxgmRACsha
SoHuUuZ96nkClEdeDR83G+jZc5SI09qJRmrRIJoseiQETKkdsTPC+zacZGIo
GONYRpUIh+g4SzifFr2ecdzv1SHdYsEhVjJW5zkPuG+BzWeNOcAjWpMGkIhc
HNaUJGAFElddSO6dnKMGMoWBbCXO4GdrqVmmW2USgDC8fKHUTwFGTnESBNYD
bF+miqz35fsW+UY0Q007fMTINsobp4NdJCMiWd5Zj7E+0aDlxC1jAo4k0adq
ydeiHmbGqzuKksujvfnSjzXpdNBYErqkbnz2QtrPgR/40C/iAGFB6dkcZ+Kz
rlQUk7Tzrx/FUamdbnI4ZOi58EBCCrggw1ubG6BdB3hxgZAvF+Sb/dy05fpZ
NrBMvZ2Ob6INMHClbSumpTaecAvdCbg0aWKsjDnLX5/diRaYoo+s05bReWBH
fNjzJ0nYqDJWv08i1UcXTD79I0xvtQoYJPY9B6o+m6jWIxKF0MxwXYZA9DW2
5QYQh2yUNVYUQPIaW9VlpGsHS32bhVf9RHCCTZoJm318hx3gZ0PzWNiAVpCJ
0zgWLo460c2p/5cvpUNrSFXUz/3B2VCcea1EnQL91OXVaQ1RXFCyREcI1J10
XKt45oxjHebsoNr8iHuMr2pZzcT6s2rbRAgOayENpyBrLJTOwvtuVJ43Zlx5
Si9+x0gsa3F1zRgDPXZ27lS7oVQ/Oq8T3mn86oXtwdYrDDyovvZ3ZkyVIdLr
FU3x1LoydaHl9DK5KSfd/8A74Dlm1arEEOovwfIzIxLQ3FuDS3ippPzEllPG
mdkVDtWQpgLiQ94CcvCWtLyH3F0sIHb2hunUW7d8eHMydZTpizM2iu33VxUJ
sFBdI/Fns1jSj+23iJrLTv7RcGYFZzRuYUQ3YHrBlv6zENz2P0i2f6xbrk4v
H2sEzEQAeUJK5mXkyVLxR6ErTZ81LaRntDOBAE1iSho5dow1zHvveWFxwEPm
YQSwn7ubxrcrcJaLd5vKji1TiWFChI8one779x0E/FLUpbvOZscLe8/0RZGn
cSibtaA1wq3dcR9BKuBwLVvZwAGYHuERRB+k58hh6/OSkM/IslU14rzYMSqh
mwkmEXJmVK7Sw0wcOwBXoBGcUWeUAhRCST81Y5vLHVyj8Dm5CyRAl8wcfqOd
FkR68BNEoLGQaH6VsCxZ8S3rJSBGnX/py76Ts4K0MTgb0oEuQoUPGT02+g3H
PNpJKvjuKL2zzhH9OUBP60yDV7x5Efapd8V6CXnISN5UUPgpuqpDX9cr3xcS
6KoU3Sjt2LE81KJCS90kW4RER/QJsx530rw155KgY6z73qeUZ4tNQW+ZzfqB
P5sdt01TyPH6IvGzLF1RybQhYg1uPMHKoYQIjdPgp9M6GcDnImc2WvfLIAeZ
8e4XXqVDhSCWziNgYMVhLZfAqaVXrjmV/IpDAFQutGOSxfXPoqcgRV3mQTjv
y8MPxjiNBflYtKKu5YXZyCxXeZZq1FmasFsMKqCmQHgyeL6nOMHx2Y7b6Mjs
Z+37h74Cmmod5hiRJ0FMZ3ZNUySuRsyHQSOYu08dIK9UNcI2AAB0c/5nee6V
oLsvDlln0xJ1gptWvHp0wegAywLhaVBjaOmdm1bddC74hfPORMGusE2FJ5EV
K0dNM6HO2zJhnHRdJ4CQVcUO653r/T+ilzpAjoA5xr4e89774IOLq4O65M37
wzBBcRRtZb2iMAvzHwGBMk1ffjGNxvMG2KxAB4RExpIRq5sfnArE2SdVRzh7
5yvtC8k6h1zvtJtn9YIj4zMzAhrY8zv6OXgB1fZVVJvt8QYZjYETcoVkqIcH
T2TtuqIxdIaST2gcycjS/E8e90gTr3Q4Lsbd84ZZt06im9SR5x7qmrh7tY/W
jz5fKLQDc7yog7XQlhOZRfDl9FZJWaJnzf6RVUwvk9uQd5WuZaX9y+9XVtgS
EAFd+TmR5P0d6PYU/1ysBDO1dTATeaK7J636KZrYNaDW1h3jz1ai4qf80KVs
tD6+ZXOl/KA2nx3STGFaoaVhoemrhHVNqWlWVyz8tVs4J5gwLwV1JtPGCmDb
T6Qus4XsoY3UXYc+f3V1MOBzbzgMs+lJXGgVDfTYN+CEy4OCRDrP4r+xkpOo
BnMMMznyPZoUVcHO84A83I8SEYOFWjScB+Tre3uuRUmH4j2nMDGBLQJ2qiVu
PJbdoIqyAQiqBmBRlhIffVUL5eAbRGPHjwY9JgFDL6ylLgO8b6PsVQgTBRwC
0Hfe2I23RDm7DAaAKTf4QldhopSx9DbpI88z/wcmKsUZu/aI9ypDT3JDauy2
XDLalWvzCR5U8jyaqNADNU0yreK4xqRSDjbiunoWUN/q6ctEoflxrum1G+9O
coLVaxB8S36zlOHi68jzJa2uL4QJ89jEZwSjIOYT+XI+NTu7vqZyiXYwaMmi
6FRJC7XH5wL130/dO0ld0KEJBSXZqYc4hMU45bOwqWhplM+uZoEzp60Ivcwf
2+XlS4jzHNWDPBLLSaN65JOvwGP2RhGmcNLUNDJqd3QjcVtg/6Rhx+s+49EA
YJvkWB/uo1UvOyy3y3riYr5DfH4uVL/13sufqaVD/cJawQzuAOdjgwlnI6Ub
cUIWO0di/Wvzk2lgTQP2grovW4i0JDufR+BL66NLGo2OXlk10gDxoIJwBrCL
FZWT6adGyfMaMFgNZoaHVUUUdg2P9ZovKuqn8FP53NO74lsOD6h55LAeHxro
pmTD8rcFqPPzF42rDcrQozhaGALjjmdKryPZtdGz1FMitin9MCjkRySRyiDw
GleLDH79frX2KCHr5NDyhwMnxiDuAWol880mFdN1vivnQKOzd3o8Qg1hzFn7
DD7J4Emh3d0YFQh/iqT3vFLdWaMlfFGqfNOab++E8VnsC2Tog0NJkYrhW6yQ
DlApJuwNQAik09tR0Sf7HbFhjAiV8YPn3PTprg40f2+pcnzxqRnfJx+o4Wyd
0MZVhWYTUmk6AEgRuSkt7IJTkCDAQ9doKnTS2VD6YYHG6WJC6vJSVa9xYWVm
vfJv/12JeenDhoyhs8ZR7KPW2H8SoEd/IYK1p1O5FuOwZMAdgQZIsQQq2Ywm
Yk60j2DbneRIIK93ZQVHuFgI2TPDioXDzBjw2GvjtrCB/bmygK0614WlKucm
30s+Zr023NbL0VAkOR5f8LAetJhJ28aUb1dbGPSkd8/G1hcy65xNYGat8mNn
ydtyqFNMrJcycu9OY3LqlykOOiuKWx+/cfz49eA5fLJDhInKj6DOnLYfMN/E
MhckCcdfFVB2Fw+93DFbCWoY2j2oAF3BDCmDelho7KwDhwJnNryMfyR4kzL1
KJ84tOt3D8b1q1U3+3ptR8JHIhTK7EIyk5F+bS95Or8fz71YrRADqANkmi+i
F99Ss8LaFPsgTOZwcnTLdlGiM4Gyqi1mcA1JHg+NrDHhnmZmvRkMfl5ZaogR
1Xw6GJpoBGDXAn4on3ViVIjpZwiITMM7uy8F4zYHCkALohE1OcxS5uK76uNb
JVWIfLLcV4xuWX/sN7O3W/+GZo8rjZBUFIr8X7pCI3cTTaj497+YhSctqucd
CNccu7gcWmW2+px6wB+o4DjoVFa/poonXdPTjQnAt30XWuCowRElbP1sOfdd
eeYpM6HKmB6uSpWI191PCdAE19GL3xkMclESBso4U5vi3JQ5Tx6Po78DT1CI
Pf1OikRo2HyZhAiRltP4Rpqn8kYrksX2uDJC6e0NABLbjeDuIasIf1hZdQWt
8xxam4Z1uo7uLv7FthTAO6OUSPuOtaPwKdzXPvzr8G4hBSAXzwloRsyb4cyr
u1xSyaXq8WQgvLufp4Vrc1c9YqNsEuUmlfZE6ic67DTb2zvIl1gKmv8dLyTz
DtN3rTtoidBpcyoPJjjhOLznvVkpHjaVEwf8XMgj2VToNMf/RAtROYvBZPho
1QYooKKpGsfDKp86mknrMLSDDuoWtfx4v5rwGxBorsu+spgEj0N/1uqof5Uu
fB+kCTz7auiOWIRYTg56H9P6Fs+xxDfKShPn2QZy1C1uCvlpo6D9CRVCcxxM
S7W/Q536axWujPrYxIVtB6WPMyeFWK3Ia6NsGHHqgPgDAmz4g30tZDS97c2d
+OGqPmBhMyvg8ZH9P/iP1fX0bgcoQOj2c0dXXwZSCoveoolWjWn3QqcCwUlJ
mPCMx0EdqPF1xjKvJmhVR1Jhn0HHkr3O65v602P0T0hsEWyURCj7fQzBPkDy
hgTh6NNGTsFnY4yxLfLh1pdWLZwrko1344uUuZDuumTePIRCMYzCUHxwtxII
s5dXOKdGHdcke+SuhGdX2mRgOhwy0lF+rEQVYsnaYinhL9q9IztF2WhCigzq
GYDroiv1Yzja6m0wRB8IVLkLsdvAIHCqP2uqzb4Jm5l1UPUJRM0E7dT4H0d8
mM0zzDH12m338qWmAOzyae3wFgPlKEhZgNfhJZxGaJdEF+zjQ+N3KPJwS5Zv
lPF3JFd+Z8iSUFILyP8m3hlmiliAxMz09mW7AIZQeaGVm4HiM623VR92+5KF
us+Adq4rMB3UrPpl5g1lUf2vMpDL5EbbqdAeeIgI2LsJbjbt77q9HOCieC9m
HJ1wr8Y+jsql46KC1WbXBiR+cDNgkT3ht29O6YKI+OmchZhW+Q0/MNMdOTDH
v8bjNKnYfsirnYskrJUwKuMW6uwA/9i9GIsuVSjQnJrDLhy0ptP53/Eg+P4k
Mu9ZEgjkXiszx0/gDNgzkX/NTtm1FDrPjr8tMO1CzX3zkyUlZVIzWYYdjBXk
yz1vkTXAlSWUvFfqId9pg+DVvxHM9KM29o7T/bAEkQfPTa4wxeKu2Po/vYC2
hnxt4q9Jkpe+m8jTsGrT2yb8UcVmzBYA8NykDIcgKMztEO+QNmOvv0GRv/go
gRkjVhjZ8hHYF0Bku7AMlLUWCxAso8atuboal67tA9yJnWLseINiiqtgyJ/f
15mQ+Bocbd/6YGS7AgCqaW/qNVQIcWlV3sjDKi178Qo1G9STpypEgIqhAVM1
ghMF35gNSVQ3p6QP9UNRhND5GLQsctJPEm4+PK2Fepijp98I8764eAXv4hgX
7KZg8Mr/zP+pqajwI4mZDfFuidb7VyxHWq7dSz6BtWKbaRGx6r1cz4/98Kqo
nL9nlsKovxFoK19A6vzEH//16lcXrBsd49DMj3tbdT3J8SqP8CWvCT/unlXy
xvl3dogCe5aPNVhXVZJW6Ubgf6thxljeGj+4dk/zy+YKKJ4D0dSCtAzYSvj2
HY9mGCiuFXa1lIeGtPwo5jy2x9Fr0fNOo5d34kRLDogRkEA82vrCcfNPg3VZ
+dkU2ZV6KFat5D3eTg72jXIIrtZwT4dVN5wg11gZeq2U+pWwgDTrm9vsZ4O3
zVEpLWUs6eaR5igWfn0g1Ubvhq3ZkzlodHw6uzlARGd+dlLN7+8o0SQU7RoN
e/63St7rCbNcza5SSF807moTCY6bBv/n2P6ehJUaFeMMGanZfuK5b/jD79O3
5K2ljD8eCHVr8MePoCPk056TN70v7TzJSQVxWJXZOO+iwuPvU7HfQq/Y9BrS
29hHhL87A4dM0L8t+45KnQS/re5TDv3XixDUzf0ldb2v+FUBfkvpuXwc9rlC
5ErnxEnfTAx+BIJOayBh2oDJ/Ilbl4RHzDaX3CeI+cbMR0ZVCWoYHr1DA4S9
KKk+rOzKG3aplx2uI3c+dZSdPeplzC9eqNRO5v8KOci2H3ChPEptn/OZO3Uo
10VZkGpt1RH+q5yNehYE7MDs2zIhjzK6U1c6Q75iB9dUpZUhnckxp3SQbyEA
lCzKSwONCk/MfPQZHt/kcvDdzgqnRyRqqAiIPV1pmT9UzJKw6SDvmyNiRYJx
2kU7S6BZNu8sL34sW/wHGovNawzroLG2EdkX4qDToMrXPmnmkUS6re/UhqGX
xgQI4gUn1Je0oGz0jiOj5oviXZevTxxPDQA8Vb1qTrus0bm3qPuuaCaSCCEi
gL2dzSvqLltNq2V8mTb8kmRhKJoJ8mRKjwnBnR5o0YjYxDVhSiyF2SvNIcRC
DHTBz7d9ulyyh6K9AAeZAdE5pKcQwAIdMDQKuZ33OKjmP9GNLBBm/j75EgBW
lQ6zQGsoQKx+IfwhtPag08GzGzvHRliCJYgPOy1KQl7aGktpLPRxwSbnZicy
EZkGmpKU/ppepnsC+dHHfLl5I1GZns/RTP5v7npN8RLhn6LVUcSSQyMkW7IR
6MQOnCpEqd01Vm9rflabi+n3ycI4D6v3ISXMZvjyCGwb1Z1FfISIMO/WXTm6
Wkq/Yx4rWrlckLrGz0B6tI6CLlksD7NMBCVh3ud7BdPNmKMjQWBRhNXFiLSa
yMIxTzpq8gQDCzj+KNZvCvcq3RzKABF68Xe2Mw2PN0dD61eCaJhtuvPVfTSc
444lvgGptjjz5SHMGVQhk3Waw1xGbKzGl56tDNWfyLz9tQ/OnS5qcWJscAby
nQtJBmsckg0bTBjivH5TZIKBLYzUt1m7/I/3sSyB3MsnkibMom47LLLTYJRj
9LiOSlOmxeQpW4ZxphM5ELrbyScvA6HEWKsN42VMPEp++/XJelpKAQ/dI1ea
p5e4Dc0gGXVA9EtteGyThUj7wZ/J6y32Us+d1xT2qNVsljWs+YTAVUjw25TZ
qKUoCkj6Ud0kKu5SbYs+cBLP1ewjuxzktNdCALLKz/716gcmqZat4EkVlYkI
UcHOc6FxZBEfIKZJP0b1EOG/wx+XzRX0TzMURo0kNm1t/Sf72IoInFEOvYEq
nJ63wDmUiKi5DNmvghmQxNAN2N5CzkCXanPVdYafnoCvePK5dAIo4Cw4RXBk
rKyoGt6ugJY/Ss/rHAdRtsAOIkcpNQTdTgUEvFlCmUvv0FTVpu4xBtJJd2Ze
pyyX50J84ZQ5ujlESzPxBrHI/QJ0rOskoLilkJm1SRVxgjkeXV1m/DuYgSNZ
3R9I85OVcDfCBP/5wrW8ZkelrUZi3Ca+v7xX6yJ+zndNHQVOJBrMrS8OAsIn
NDukgLB0vIUfOv6fvTtOTYEtiTUAODtK7FVu/c+nWKPgPqqoAkoAwiYiF8hH
QMj0qbQiL8mPij4JTAk5UTFKpEUfZI2mWMoAONqXofp/vvjKTCa3zDAdKN6Y
Z+7I/ODFGn0FhpeDOg+NQfOQlu9Z0JJV97lCotzJcCbd7pmKK5iV0csVfXeZ
dUwr+wjCxscuWZlQASq45yZ0U88sdd76oHF3zKzNltwPMySjhp5Ke9xLmVPz
YyFv6IOYu6ITgodsfpCfgOuwUsu2Y2bVVZbf9GvpS/gNWCEFvCFAU5PIc7/f
S+CnGjsU/RlOwiMD9Z/+j2Oh8WzBZRy5wjxHVKovM9i8eR9F8hyZ81FuNwRa
utgBd6E6mHyx2LQNwuSMWNk7mjpLo+0VeeP4rjv/xzeqrk6zL7Is1wop6lCO
jSotzrpzvfdK0BEIZRUhj4JrArFpTbYJRFxRJFb9qWmmyfjCXXzhrvhnXDBx
w596hEcgCSmm3s8gRjxd5CKMvHzbsNAEylXcVQ1tHofRcovwHDoV2LA8oVSt
mVLwrTU5hEPrZtBMRqROKueUvpQU8yGZM7UQitt1tzmb1fql5dRk6lMlYY7g
YhDKahhMktOo5i+wPZo7sx/gQ8AWJiajdcyv6qq+g9FLp6Bhe6SIjo194/1G
ueBf6GV89Dj/ZJ8eoUG0dTCiSYtxLUpeLSx6f4yybUTg7uHg6mXSswjWxC4E
PLsaiVXBQzD0UM0AtW6/IkLI69GqLgBKHxegGdM2A/UlPDcfqNrXH9s14o1+
C6dizVEIdauLEq6E9UdJoLhmNcIdNTxNhkPL8jbFmd+++0O216ClMfQUOX3E
p9wfoie/eG9YyE96k7Km0aQc4m0lM2HEWWXJTSVIw47dIlwVwb9b8WDwjYIU
pM+X/7H2oF7zM1lASsUU1rrXJrBu3Jc5DH+VnM3GO/hcO4ipr/9Wdepi2MO5
IueF+Jh6WrP/zU6ingZpOOgWfcMCahW5CG8EPruY4m9qbcUxjAPF532acW03
eYg48JfSe5JJSq0LVwHkcaRbOzE+jiMaX2esXkqXdNRWmFbkitD/1YD/PqSW
pP5FKocklPXCO7SfF6jOaesMVHoyTXhmO9nn39sO6QDCqgqawL6nyiJePZBv
9xlecQ1Sxa8K6PwT6KVxWUiwbQV0oEIpZ107A/wcfRQZd0rikFAGRp/NNLOZ
JKslo89t/zuW5CreNYjBgoUtgBMo2cFUyMatkLwB/VoGwWo1qSSkUTupMhpW
T+j4kteV0iuO3NpgXxMQ+CZqikB/jPYji20L0a5umUsoRbYagJkW/qYn3KzR
1h/M3jw4xw8dlkaZ694dDVAL2gYcy957W+UwsPIl+uWUJmEb/kkHpbBniFFi
tqEp29BUIMJ84ypSDekYlc6oo8xm093WCZnW+tzWJ7u1OhElugez9PLXFdfA
Dbyv+54s2szxiEWnyHBfgixE0A4ArJP8CW0lercf4qaXDmRzp96f979q4w2O
capRNK11GToq1zxISrqZjqMNJgKW02pg5iu9I9puZ6QeBFU7Gby7p99hek2Y
qTSTCIOUOHNmFtgClxIbPQmqyoVPm2TggI9Ckz1G2Y9EzJNk3F7vsvfS7sv3
ZX2OdWoz5WXPXO59Y1Q8DELyxmnxkUvCY+RBg1zpWT2RDJSrl0NR3dd76y2U
N/DGoypwHT/YjI9Pv4eq25JL7fRDyJFgaXUSxDRbV1L7opNhMMq/qqCIPeRT
TlIyKsRNgZTqxp1V9juqNH2AYy7jAZnfB5bc8zrVT1+2lrCe07G0HmxZhZmN
f3Xor2sdkHNICKwyHT25AdAsG12iOYDoKRmMC3uIsBmxgVC4+8HL8E/b8aZ3
UASItST74jHKDJLC6N+RfoOFlqqLNx1agNlfxe9/0zAWIEaz4T0FU0xiNqpS
Co0DSpJFZuR7khYIF+qWizv2Vtl/yekBLViZMavK8OnwLkJSGcPsGfNuj4bD
Lsl3PSGmwsD/1LimrhA1fceyFeopyiVD7cr4hYHH9SCzugenTorWIkR7vx2k
EWsMRMDNyHMZRIYYjZT0m+DEU6xDY90IGsa6raK1PWNJUMcbBtLniBuJYcsu
EH5cX5hK4erwGV9GIj7YQWiPCY6wvVANuu1J3lAYm/l8EDoPoQ+zMdwJEm6I
qqnnrMubVv+r7DX8cx9GA68P9NuF7qHEu748PnbP51RXUqXApJMMG7ilP2If
HAP51jTettcfSvUwn9tuK+8VgNshrLd7oFNeRftZXKIBY7POUaTIAZ9cvFCJ
RmFH00Pnebx/xaen/5Uq+BQcDPzjGGqyRXsfbwMJvhnMeMV0D9QIxpB8IKn8
x1VW/tXwohdmf6G/Z4EyUrr3QiiBzBmf3Ugb9zRedKbLgjWdvvowOJ1RSls9
69DBD8rfizmtg/Ee5usWhupBFu22dj06fgXbzH5UvHD4cHiJ5dRBrTghYcPP
sOWfvA1TZjgrSX44/RbZuJAnln3lLiSmnlPAG8ZExcBCJTWjJbnSNjeDzjLz
GYu3Fpdko+LiM31vf4FLFWq1Kw43/QfEsofk/wPmf0DUtW5LxRXNf/u3ywV/
sP05MvR7bKJtfieeHdwevF4nmybHKPzCBMmGoOnJ4g4urAxeCPsBjG7M7se/
IzSHmME9f1SmgrhMne6ZkjIQtTDJmtviPokZXlbF2F6mBCgTKI5GIYcF80Ra
+21so1oFwHL5Ne/sisVGsbvjcxhdGN3RRhWWioVkkUydvjLYx33CeHhkey8d
4OVogoXNMRCzuFRwsCYVBu8N3zDuBEYQpFxfPlAVvmFe/apDudipS5NSBseq
b8w0S07G320WRXjYprDAVPIEJ/0VbX0qHRzBmWqttPw3svmmva/uyLJjCX6B
GhW6gnFVrNrsLveczy4fVct7WcnAVJI9/9eV3tQ8ntNh8n52t1mSLYt0ORzA
/esI3/DwXmO9k69codJrzfCSqBR5UFkpClpj6ckx2NW3igopnW6/MMMaivz4
6UeVxIoh0rQWVRIv7ayN/RV91AvWv1e+auQVjCO7J3xxO1znoHUFiHgZ9xaS
WJk6+wVEFG65qAGQ/zfoCzoRQZ+Ot7ZgyqJSO2KoSsLUq2vAvc4XrjHNs8ER
NXI5APGXcWe/9MRt+646cnpHOSK/ElxmA9XHTvMnhgLym9760Ob00VCTmA5s
75YxYeK6Kq30bIFAX8L9/OCCpdwZShQmUHCepB2h7b/tsVmhuJuP8V/99uLb
URl/ObVFsWRkV95uz4rjgVeaexxpoJ9XS3/k+cfnK+Vf5fRCAl2VsYGItzf5
G8NvAuDC285kZa+1ngY/SH7R46y1uVMB1es+tb97j19f8mrHkP/alql0iB3I
3S6i1U+YBqT2gcawFY5T3UfxDPwLb1jhzdDZQ3MgpniVGtrBd+HuJlEkRIM3
nptrd+pvB86sfonqlH8yDOWYDDU3FTvylZiflSwXmICneTpfRed93gwSd50k
0EyB7VDr3HczmxQSXF2vcDEfN25wda+gTHl8O78sp9PxO+5MXpPV6SNTk5gU
IQEiagp8g6K2lrYSmwcQcDh6B1wOe0o/uYPb7bXnYEifqV+2oE68iUJ1DXAe
Jh0zU80Xox8zd3dZW/LgrTflC2m04LlDDw6aYhmNEiAmKmQY+tmOJiQmz0rd
6VMuQ9ZZeoyV7m5ORIDzVYgfEN02N4POPyCtBPSJvq0IvygbHDwhQuLYPWg3
hTnrxAP+u2pIpnXLwwGd6p7PrqiWUI6wfBbNdnNCH173NSz66dQnxn1jvDt8
Y2KBBEtO/79bwP6EL+pnJky2zUWBdu6yuN7hiEiwhIdwRONu0r78s5dLT5RH
fZhuvAefYImlWFBv8rf2qUWlsY1GsIJdHp5E5QXfpTMoRQ/sLwu9jCyIy3dv
phi8vxwpFcgxI0yNlIti4orJc3T3ynlxufLJr94mypZZzkXlaNTnGU61hKTY
/iVg2QirKrNPmKildiho6sDTeJtbBRPbC2zabl4kw2nJLIN33mYS4z3cBn3W
V4IRSyQIV05J5YbzVoPyfPGU3vrAcTNn1XaView9wqK39sWrFbHmRV4y11/r
PRwDLvhKr4v+0yaVE5w8bKXApWp4HOZrcR7DaHCn5RcOhB4IIYyfIn4MpGh/
6okhVpmrmeBc13gDIZklh/0nWuxxqj17BZfA/EZECMJ0eMAfmJ52SBIA1ULP
TaD1KnNlFQbuVdebZpZvBckOtWSuO9yREtWNcTOHX2jmqYAKPhj4xKlGoEud
Z6YoniPkpKsdDO27zZ42ktAvV5bVgyAtm8+OzeD1lWXKWm8IlFzXSXTBvGT0
C7eU7oq1GAts8500jgQ//eAdtiFAt9ZQs7EQgAMg8xTY7s2ny24o173lodNu
CIlrOOIk/XVGBW9erJsXbNCFRcjYwu+d0zBTu8Q7bmDUDj6zq6gNs2bTR7cs
Bgcorkq1RMn1ge/4EsS558Tkmdjxw+P9eZNXnE5DoDFkJqCHZj4rSXtXKxw5
UQrbaXYvKE9gm2pax4NAPFxKiz4hpuEaoJKtzDgV8j8BCCmHyfqL7dWi61JG
A/JVAV5uLPXnTPwx1BoYZNoEh3q9O3uQpL/XR2t2jkBLlkyHDgIpRh2ONA18
EMoc0MxxIYvNtqIpS8TVm+kCbmHNqq6AZIwLABSOdmGTJdPMDZocDfcQoXbX
Z69s94TF9osfvwtXFeJOZ1yav9uMpnr2sKqotVzsAR6j8EEsfU9s9BmGr0p1
ZrDYe4py337Cwabuvq0p1GH/ZpfIK0e9X2cqbIDUlKf0JJits+bC6tp+PhQt
7mQNS8J8Jc/r5xzsa2TsD7U6hUVQzLgwnHgx+eWAbqJfR+plFwkOJcc6AxpX
CwyUKmg3wDmOZOxSwRqo7yVqly8fMW0S3LxBcH69nUY1wTzuLrn40+opEJla
OUAfS83HJHKNfy8BZmciEgxHSQjlkqqFPQZgQg9mTUvEas7HFZ2z5v2dY5MP
feYkwyMk2i+Kt0ZtqbgDVrd0VcPAzaAMeF3urvmc01sZRBaCUO9fDEpqQ+ct
oxIDx9GbkjSiP9GSEnwn8090/+cX97545AxbDu+hnsOatCGRrQUFj5pjVfSU
4tmrYMOVA7cM+iHetdANXRrCEu/dU/sSifWSKZwB0NIp1JERM3qiBOKiBibK
XqcFUJsBdB6v7Jjw7fDF5kMS+Vj0PWZhUuv2gtz7/75wGxm0b35ERBIX9tri
VYxU1acmW7R/pPrqJeO+KztIHzQDt6knBZ7a8/35FqgEe5a5AnvuU1KCJBEw
TNPwRpuU//yNKjOHv+nKNewPPxmcOFa5yJgqOeSbi/19fzCw+Hon8khQMYe3
aD7VsIWHai2/7cbLGJzz+rPUx9ZHSfRpZRD/gj90jva9Bdkdln9Y2boJtnD8
Oj+Z2y5uwWGGx/oVzRtNUoThJqW1a4qfLmbR2E2eIkCMSO9XMbiV0dkaygwU
puCyWaB3+qmbPcN8oyhStfPOn7g44El6qmmOOMCy6QtiqfNP/RXF/5RKxact
AIxUVG7DPLr+IYLyFdt5q+1mAg4EfteKv/HPq/dWhGrek9WulPcKJweeKwZw
yU6dOOmmcLdniitSeAhRbQpYFh6RRS4e1L+x0Y+9IpcSb+JxpVma7pTTd+3R
TsyTAlQBzgPKYEl0e8UBfEkd8rkCqOoc65cr0boxgOYSsylkaQ5og9ULl7Fg
7StOhEjtJuo5/1aoRBc+SVYWczkg82NWDE66DvxHJlFvxFEiyUr+ShvBW6bQ
Jm276cR0cKw/Rz5CVhKTk068pDkH/16nBnWbB6u2B1pHry2g6kCAAdmI6Xu9
14oHtn/gNkSc9/3Fni3vbB5AqtLYa/DMm82ZUStv4H6GX8tG+L/9SBzd5jHE
WeHjcVWDQ1n2EGUa8q/YIBiYtgMxWr1ayjGraVdiiBpe0mFguF+GmechstnI
EmuHwU1DHgZac4szgYBDvbyV8sGWkdtNYfALdDyQs76DV8pttGmnXXfAvhkm
FeHU7z/2E9RP8FwIaArzsDyaVJ8GFGYD0UGDwGH+qXydMXm6yw8Di6EhkpxP
UK8CATi9dUwj1n0Q1pwGw2w8HiwP9lmu0gwz0TCD78B4SfDWW67YtlTwFyb2
gVFw96vECdkRdgMdjruA/W5KnjaBiRzgYrWyoH+lqLkTphXnv3uv7BgF9bxK
tHw7i3AbP9T2JuvfJWKrs0jqaF1T8veI0ZH8UAklsEhp1Vh4Jfv5fZW6P3Nn
wtmzSGwvO8/gredhgscZ/+k4BQXtMVJogfp0jqghhRlunpG6/GBoWs1dizra
pg6B8h5WCZMT5mBGr3tAA0iylOKDzTG5FIGYAgI4ks1ip8FXYXROXiaS9Uaz
yOYgU7XfDUFJI6xiDH5bebprYVqJKuqX7jJXPNvVDF4+P5Oa1TrrCoDg64cg
PME1mHgZzv/C9NbZTrQgptYfvLwyflxdTReRQs+xhXkdeFmRBlnxFxZO+42S
VuWUPWGqvV1s7fRqOsSuIoF9fQcYmRtwSAQFPk/u8KtXpEm7y8Km9+P8AyYx
bUUsTNSbUdd2mUhoY8MSAIoKVSItGybPIeNuq5vJuAGBstfBnvsydF2UNvZ4
pPImXOEVRGg/QV9Y0GldyvJD4/d3pdP+xhr0NnadNXzkV3D9wFJ5qbKBRKhd
sMhCHLvMEqkRAMnrZb1u14FhFl1Q0+0G1mOeFtekYrVhLqrfZYWuiPUxaiJp
Hvz0khlKHj+nd+XaiwV5nWlr2fqMFfEmxD7bnj7ZInTnjY09lxXi0FUq1m88
QygiaR6OzoHYl6Tv1T2XJPKy2sOozp2umM4QIsgCF0S9ekzA08T2f2FAbE/w
68U7Fywim29+guMGUUoW34q8oGAIUMU88MzH/0QSJ89vzg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1JV74dnZAQJsRfphiXZ7ESjYp5CG9uHr5Nw5JnBjgYz8iJI1U9Uns+VF5mDDTEpO535cquCbeXbqS580erhQdF8rog6YD9kr8WiWl3HKeNMZ7J6v8e4KthPfY7Jm7awMyGmBqYxRRTutDAsBMi1FTKhEdaKuBAoNE4vDu1g5iK4l/ZFAbH9a/n/WA1QvbZPMwgJMEh/et4DGK7kHinnSPsICrhG9Ik4PZ2nO4/S0MKN/7xBTCPqOugLApHMEVSsBctfoWMyKZa1AOqyJodSDPnvnlhhR1tSWVyHQxdrioO+J7JMIt3v4TivjXLRBoJHxK8KqiJN8pNE/RF/znES3ejvTqH0BKgSHvB3lTZYtF0pRucx2ZFqyGF2o9k46VM+taQEi+ZYrPP+b4xhfvh6SB/LT/+75uNXCUycCmmt3Rm3u72K25/SV6gzPC0Gp95OV0eCO0ejBqm/oCtubz/duvfrlMOdBL2IB8Dz4emznkBPcg4GjJDMRkEW1IAbDxR6RrgRAnSjFiQjuDHgugDyN3P/wzdE2c06Avsd5phLhvNIWoeItkvlbPJBYYK6C7yzmEwcMKdUhQOEem0/A3g7d3TMz2prjxMW0CQOgH9YZSQYpSytwrbL4nocDWpGVDNodbnatp4P/HIk8ac2LpqwvOzXa0nVPiz7HIYD40lH2uu45f5fQMytjiCzs1DKo+/kflF2q37HhgK1LQaExXbsKUgu+J4dd19spZYPbaYUzDh4n0G6Bpoai29Ukg5V87k7XYXvgRTMsw44VEg1wEBnsQo3"
`endif