// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NJsgPV0ixQ4cTn+N01Jm5poQSsN+qcfHUJMwuI8XkWDz8Hx0wkv2WLXEtTiW
d+//OPyAaBbktVtY/+hVrkkF06i39cbEs62A9XqT803JIjQc38JDGl30WW+h
z3+MKQKDX5J5b5wjzYAsxLPI1CDnoaRcapJe89L6G/u8AgWyNwhzMBFEvpwS
mXDr5lAOEuXqKicff0iU8ZoYDsXU9vyXDwsAhv/j6drPUsqW3fTnll9HhB2Z
7X1eik9e53/e51CRA1ImiB4mmzjFbVdxn5u6zcOBxYe+sv9wFP96TCcrnzsm
puUIHUntZ3W2oqDhUTNYEcaRZfpEOxVMLY3SXER2qQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DD/9LIQiWvcLCQbZ9Tp3OKgIw2aqm5vu6paOBI0BLPBcVopyJNtFFNUXvGwm
LGZ6hYojP7GDOKwy5wsodgyrydFM8VakG0qaQjDtgupZvoEUHJSoSn88p/QI
FrvF+TnxgTUut/tl7z7ODHRTsQBemaEGQJOtSZCPiCekahb9tn87b9xJ0H3O
WdElPutKZPvPeblPPg82HgH2mKxIfypZxhTMyjD3L1uzgCTsXaymjEFRlUp+
iVbJe/yQKRVB8udFeN47TWsq1UDE/+930I787BzWSPxgqJCQf3plEcc11SD8
40emkf8zAMTw+XnBONeCuG0NLMG7nwaa+NA75k1S8w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bS9FCdczXAg/2QbvFmtWLPP7BlfzJRZZP4S4EiV2JEEaEglGm5U/h2Vi665q
AOrHHRjaBBRjDdNXJgXhEScH7qWxOWS2Cpw6VYEgzkajJDv7WJu+cyiCUolX
4+eCkOEoh7I5EJF8a3KuvrC6wF9RnLK6G+dUimhdzr/x4mL8thJ5LHcphXWy
RgAqCKmIpeyGnvqLjkF18U1AU7ECxf1DSnzy1vIDzX/8Am2VMwz8uXpoHTeF
YT16ydMZC0TozVFFzp690I3dp+/9Tz0Ya8nuONUxfWQMzOmDtgPE/b9a0Za5
ovQ0q4CUqEfWj5wDUvL77l7S5EBvjUk1dwQWXK31mQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KGQ3Cf0UBT5cjP6o8t3BCWJWOz7vYVdZ2k30aFYT2ulGkFMWzrwf+GZafAjJ
Lruxxs5cksENGsHZVJPJr+TtI5uEhihGYeh4fNsxmhyZlcFNDf/W/HEfYot6
PRpZf9ND/HUnynH/4snU75M4HnteyQ2kFTRdGwwddizGBxa0WgpP85Um8alp
PvTAkR1vvSWP9i8J8XOqE9/HKuPWAgfJhRxUGoQCAv8lFmrJNcTCJ5BVfSg4
zPA83rwwrvC2JNL6MoTw4ovr1BhTxDgHiFBIasDggCAJxo8l4I/mcRBaMbog
oBNuiMVFhZT6dcB8Dao3ow1VssPOWNqiGXkg+wbObQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FTqQzClS4b378Kp31g9oDv0oVu3HEMRaVvX9KmoTpTLRaCJengeM5NnpBA50
oidQSxN7bjiPl+B4oF67BiLZGFbIQCESWrq5l0hv7gZr1Ft7oC8XJxZ8LZt5
JOWrS8tG1/93e+ypN9giWirWaIMcFP0g9S6MuN3DTTYpI097Llo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Y12UVOaC/YtpS0EHqSBe55wUH3/osY6gxPbrXEnl7l7qpTriINx1Y6Z21Fyo
2TmQLekDyYfa9X7timLHxwgjBKvtL6eRoA6LXTcLEI0f1VYZcFiLdptjdBeE
127Bpj/pGVPZeZfToc2dVI+MRDyImi0P/UEgeUgPm/YJz13pYQYhiOFzAXaA
yynxkZP28EsxpUwbLIJxGCdCIzNUV1oeBvv687J5grf0nBzVUeTIScOJiUFU
7u4WspJHCnpBY2GUZx+8BlsIvW8V1Cev73ZClWu+rZ3eLeSWMxBQzWanrjE4
5/U9QgICsi3+dqJWufv6TSnefUftzDzCLsFSXuzCHbnf/vapf/nH20V6ZvHa
ti5J11+R0Cja6OEYcGpW5hf9F8M/aen1v+2rg9SyTWeOasZHxNohbnyYAfdP
t1NspOzRaOFrtvSOheT/rQ19O4ls6naWiXar69TXOLh2An84C0GgT6t9RCUg
N2ACa+5CD4Qx9TPXmZG7Jp7tiONM0R2W


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
m3PYJoyQhBxIBIcGgcPM68BBzP2RtFd1o6z0V91M07laX8csWypF4LBYh+Bo
S7bPmOSSt853qXWnWkl72xY/puTiLL0Tef+CYIMW/WaD/dAqtoOYJPAauDZr
myLyUSFE7s0/yKVeUVrSbqG4El3OKYznSb85F4xWEqWls0AiHX0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AlQ4q3Yi5Ujs+31oRNjZ2ms48LENxs8aOHZBhoFF6JJdEYfZscAMuL3CvNnY
m+gsj/pVptlW9IIxiYF0u+VfDe5K6M51bO15Zqx6E+5OT6jyNv9OwukwZpAd
GHSPIDYuup2+WAV337EFGJkR4dcXAyFH11brmjrTcQ/tagrrLV8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 12272)
`pragma protect data_block
jD30h8STUoSzFBUgU8NrcODXUFj7uNmS5EpmAabwlEXvnmi41cDu6O7tzEMk
b8hnnWIg0Cq1CxwnD2KZg6ehgpDMDPSxbl0seKRpzUkGV4PbZvQSuVWCyQHU
MMVnlE0Edu1mj68b/32TFCr2gmEAkEefFj6r4V1Bvc+tQBLs/Smo8ZKHjFWK
tw7s5DXtpT2KIj2/tKDMGzs3YVXIIIkNFsGwNMTzsSArNDr4yy+cvUjS9QgM
hQT85oTiiOJ0USOzGPhDAfpzwQv/qnTqw84BksFE08liYBRzoup7UhRlGaw/
t+mv1NaA9hP2Bd1p1c964LjdVJEL7F59QAp7Wxhw05+gcGyk/yJY8tVPqll/
4W455+fxaxuoJaqW3PduUrsCAC4TMgT1ImGlSwrjs/1FIUgDbVXKXZZFkHG+
DghSF2092V/F9xSB8ZcZ/7ctrbeJX1s9I+JcNw1GQOaBxvvQEc1oEj7RmZf2
wOpamkjBBTGOnjGc9ogDUafgsH/h+XFdUuDhjjSAcbqbljPVmnMvKW1GndFN
xaIK+TdoMqNiHqEnXyUFJQhuQfe4WwER+5oYzNlZGHdtJWwp03Cvh/F/mLKY
XKhNE6EqijR1B0OW1WDxg+hKtXvAXmphf8PnFDFT9EnucYl29IsS3hwvcPL6
EN1AcsWlitGwm5rP2xFuXLU9/DJCZw5jw0W1HmZWhsOQTYGF1Y3OTE8dIGgU
lJlIYDT+xzbsM6iKVSpdm6fJqTDIdl0i+L3jOqkQluUqNYzmOEUze8GsBvSB
glr7KLR/yFaprI9jWcdAT56hK2FMRnDYgREd/MVU4loLUzsnjqpvvy/fje0R
3ESyLh6VahbyAv1k2KM7s4iQDpX1Nw1mUG4G0j44LLcADIQDtpjPSbwhMmXf
HVLlGoCi2sc1xL76VWMieUCKjv9Zb8QyhfTVk1cHxl6RNzMLHOpIaM+e3rxV
bf6bG5H3YBCQ/exHvgDe5xGqF1A0FpJwbz03QOb/gu2uIOS6h3uNIEecqQp/
4OlnBMvK4D5vZqOIUWFEbIywCR04SaEmyfMi11iJFDBgebAGlIyjmQnN9yCS
yO1KZ3owg5Ux7mxEWEBidpZglb5+FS/KjekKRN4HlCHqzMlF+oX1nCZVSwpZ
WSOeHRJ4OVLlsTYtyP2lOB6Bxq8rlKo0myfYsV5CP5rokZ4EQO6y2BOP7IsT
6EL1peS1tYb89Bt5LrDeLAScizXOE2DtYXYa3ltb20bCXukElUyJ/ewl1Ewc
sBrYGhdla44LrEezOM7VI6LJCoDFXvuiSP3+FOXK5fNIOGVXKTJmGAX52pkN
WfM9TAv4DAvMFm8q/g1lzYduXs89JeNyrQH9AE9zOfuJdJV2Myxeac6HfjOs
zfLHD5dq21yHOLUFz+vKS1Uml6nqA1V/WZu+XkGwhlQxwVOxh3fydpgvivsA
U3ocGZNbchqK/iSSOzt93oFcqpcp1vRdRf7U2+bt4FUTv+TEUNhyUpn26gi4
zVxsmf1BYdWSLWMWAMblll8RIJn/0j/3FUBCzecwonbz+PAPmf5hVWVrdjTb
71H5q1graOBohIzKjv/CeBzFJL6tZVEo40S1FAULy+BILTeIER9vWRcVlTS4
l0oKoD7zm88jmmfRZFAmYLkoyV/r9KRNuYI7M6hF9SgBhbHCgDLs3Q6SI05m
IxjSMvCSYCvofqQk5fC1Nzs8+8fLTgr9XULZyeaswDvkH9MX+B27GyFHOQam
JjA4OKX32DFnWjGt+D7y2b1Tb5ONKIcFSD2p7+VHO44XgXzqE8IMKl8S57MZ
oJuI9ehCCIceQC6mZiVURjfL0zpaAuV71yLw/6wS6y95Vr6qiIjXI3pWWtPX
2WC49Yn2azlx//q91iaePseYRe6pRSzKtk2Of5JwihDPqcOuhgp3klhek8jR
9aYIn6BY7evwVzvWbuIlskppo98pcKcsVHtk+78Otliq1WxTJKn9kx4iYfHC
NfPx+4iCwssz/z12RV5wKdFDZHhVwED0WNrmBO4Y7k+2n68LR0+hSPiZzceE
BFNdnVo7d/Y14vaVuXVqsfA6r5B2/r00xljPQIPHG9hbFr9wUEJ9paVctcX2
wseHrSvFRco61clYld+YhOnscTYgloztuf6uGmW4Ce3QO2IOpT7J02S/N5AT
QBgkjFs2IyhEcCaIxQs2N07MMSEPsST+fBOYq2lgjpXS/TV45ygx5r23h291
E1bEpJxN2IfJdthFBo8i7xVMY2eQYCzB+1600LvbOOgybIPIaYAU/M7GPTmp
ZSRFslAnQewqgrtEWJEC7LNyfqpan6aw4dwJlTQu7lpO/wKddECx6kPHO8iS
XGSJnKQYWi948NZrn+8aBxY8mjpPyeqwbbZLaKvIgRr1mZOlpTEbx9ID49N2
Qkf5LvVQKfSnTdYiY1pFj+aIEUCKXZnHc1HKQaBVbT3SEGx1FozCz0J53z7e
v1lA9bKKgduJvedvhmZRfc9WsY+WR0YBPLLQvQu8NFeL3lGHPRGRsO/f2iYz
c94nr13UGGtWzuPmGXmevlI6UyBEr4u8IiNAb3OcRyv83vhFs7OunsvAUSC4
PrBbj78H3c3wSFESGsKGnVXi205mnAlL6zOgcpfW0HiZDFRijspkcUqtMLpQ
uicdW0O3FFtYkFyPRx3mykwuBwgUreMNp/DcHkP/9bfgoFAdnLXAbcjCjxkH
T6I5HyepqVlZzqItTVYLU7P5Bc1YmdHhGdKgDYZn2LejmEpeXayvyk1FF/sT
e5PeCWRbhZXkudwWt99kxo70cXNInkDVVKmPiRaINBdCrnGvkNrBD8wXwVrj
rlmzDmwasCZO4wgJgehJpCHHqLcPP0vbJKCX5fuwDhK87HtkFTxsfRsoMH8G
13Jo8FZiHMeNlJR0WE9oM9SpUVg21x1Vj1o04KK7vXtY01KHZmZz91mFertf
FuZk2iC3vhehD99YFBcUWRe1edllV5Li2TfSYP/5hWKxJ87I6LaQUjnIuagO
60EU9QnGBPZ9Tif2RL1ZAICgVeXLpTN9JqsciAixgJwLz5auVfE0XPezPzfw
MHEpCYcKZs1F5RgkYq8pvz1pFNmzhXctH9O1VhLZPQrEK2Fb4X3mm6l8gXXj
DzvTcUAw3wTA3vg9lepMC/6PXQ9qCiMY9ROvbJ+aR0DTYYGAoHxXwFr79Lte
nCQjmWea7ib7siYd+tWl4Gnyg1avrFerdrNDnRf40xLo3x3Qe/0qXG3PhywM
NiG/hcb9g6Nz1sZCn/If0gEl1/rMzOyXU89YYuKvUR2z73lULIvNK2X9wh4p
pbgFbFAP4WlIqmooAf92ou3D4T3tY22MngpkdJvLMeiHevGZrupffp2rpwjK
y9YtWCKI1kxjOgV6rbWBrJqC17+9bCtEmOG2/1y8hXjoQTfVwVabeCxWRLQM
/OC1IQYRSlUitdRjKyv6c44ArV1Ro3LqQQqvIwzSctvfUsKVO7PvsNs8TgGm
hDXo136fkI2ZVMP8tWoWgIAK0beLBjwm6Amc116RX+TIdeQ4SelJw6YXL/yU
w3kCXrtywigiE7EOIaH5HHMIN3DVtgxagROBbnMOsSMWPeiyz2RhH4ZzIYwJ
0hmWpqhW/gON8Lp85b00ZfHBwiyMEMrvNBxW0TSPH/EnMEbLx5vRJ8AQzz4Z
c8kLS5FBxTIuQVEmpzFgxVMu/8eE+qNN9EO8byLdfBak5nZYh9RHtEI5Z1eY
wt6EJkXD6ZlFoML5z/rrWR3Td1lMaqcsR0XxEq1TZN17zclWJKqofzm12ocH
JtqlSEa8xzNImaRpYL4m++EogQ2rIeRdISXUrJKqzjz/jWYhhRIK3YaMngQ+
29NHr1eEH9HawafdIHppouS7AwcV851SDOoHmEMptbCJ5ZJMijwDksYbXOtx
xBXoPG3WlGEaCUHDYDJcBMCmFSkWp5vRIP42lgsJ2N0CDzuDC1cAVF4MjRcU
qREJ3PNt+zy/VHlLvQK3lm6gKxlKR0IGYuIQkhp3OplsooerNtLtTu5HRgST
89JDK3MjG6cedcv8hZBcDzATEV3YhUFaXHSYtVVIbfiv9A6xqsD8UznqPDML
8hjTnSRQ/c0lyQIjX9eN/a+dB1mH4KzNBYp8KEtATHoVANB0qKMeCoSeoinT
dTlqxVsvhaYFVOmIMHunUTwlaBMMNkYLu3TWTb/WM9QHABolqeE9llMIbZ+V
B7GVADE59uIjn0a00ms7utcQe4fQVNG0/bi2Bdv9e7SNZNf35ZH8OpEDKWi8
tcXgo22PJluqvLxqDVkt+T0uwmt6T+x0xsWlu5QSB3rjOQ5APh9kksw+FbpF
pKY1czWUVYAuzTHLh5qChKAp3ZWtzPdSVZX+lalc80YGl03+EoXqPz3W7y6m
xoilmEVFI21bfXadnfDPsKkX5Og+PZ+QIMY1v0MzmxXT8gyulupI8nOem9b9
1qfcXAKc0V0lWVJ/fKhgzd7rXrNxXc2QXjmujumCfEX3uqtFbFf3Kyn5svJs
PMFQsDvzsfRJj4I5iWhpe+E/vQ/mVKBRrhMNjckJ2zXB326BMA3yLRWo14k+
MQ2940kWmIRFCfjfthgI8h1BsLqRxMZ+KF+0DnJP2fWGAS9LB+syeX7XjE+v
+QWokBj5Wl5WfYgapeqGj68ps/axRYhQnRQfGGG3iRFFL2AfLTonFzPsqrUT
ZYa9cVu8Znttx5ZR/EzZcpJSr6yE7/YDCiSM5QYpkUWzQpGqZDvsU8gU0Hbk
k7xvF8nUGfyLPxsjeZBtPydY/qZTqbcVstDODAlmSuZrYNrpqgGsaPM4Dvwb
365ZjiC6JABIa5h0OM9g2csYRglOzNifm1sM4SiG+Y+LD3iQeZsJIl8gNUmc
WoOb8t+fSN7b20mKI2wlEsiz7kNH3yt/IDlskW4CpTPwmvAHgnB/erNDUXnV
w76ZSGWvyn8CANdAMOX8SNMDSh6+Wb/nAOD6jsG/1wj8s51uMA543SVFmioH
4Wra/Ids79Bq4KRalxSMSXPNd30E02Dhyg9EOKzTsJu7vlQz0td+rsRY9XnA
HMhRiedf23XPQouyeKPhyiLcqZ5ZhDt2CBvTtoNV6eNdw+xxsugj0E1BQkTC
mfMIhPX0wNHFkbSNxcsq0tTTUh/70I1Jr3INppdfrqVnFHMMtBsQLHONeDNe
naBsuOgsCGDQkwAsE2S/Xf4gLSdmalG3RUWDVEz7XUHx1W4DWbnBo3vIEYnd
Rk+tZShUPxqy3sD/MaPOyh1nG7A5GlpUu/AoX6pIYxGAEHYZR4yLGVQ2jswq
I1HPAIziGOFl0Dz4ljkQgsS69ATQ+29hltEQYHt4g5sufj/Cia8QrM/lLcE1
I75ZelYzJ38xTsyIJMqUang1IpwmzWd5ej3t6+oqcZQ777VkSgHLYdpd1UU+
oA7jPwR8O38sOhgTrPhJQThvVX/Qsja+a07c+gpbVAplC3KfKZSBe9aHzjPr
WU5880CZ0f0mSL0D2pePLdYw5y3XV2y/FRh3FdjoB0hIThzxAGSd9MjfC5Tv
V4PHshtPt1zgVnQ1MHWY9Z+u2+eW9PKbJaWEHG560d52YW1hybdG4q7hPzAZ
23URvtFxHiE/FMEUYZ/aeqTLrIIPpS0GcIGfs5aXm0b1VqmudI5cFC58F8gt
m5ql0/RK3fQseA66jCXPrE5s1wteLOrOw2IT58BxdLziwTkmhWx45VnSpsVZ
VcSccJvIzIRbd7OX2HXhmbJb51/C+0CVdbvqsGG9HPGYT8NuNvfSR/VvfSOX
kyxMV8D1Bx4IvAzHcYoye6Qt1Je1v5q5W0yyaQLjMGG8yZYREBuwy9/8wBi3
Ogy6CO+AhD9D+pPTLr52tWMPFVw2WY9ZJi0bZeK9e9LAiXWwPJc+P9cw0Que
NjAxPMV9Eop9C9Fu66jILtAveh0MIlIR4pYsIf3N59otYnsap5NgqTIGuMDK
e8lIBDnyYvcmwcFLyWWAZZDlo7YkYtGt+S6Yiy50FdQIBpLn3uhdj5PkEv5a
muUjcyM+/JqI38+YT+mjlUhvnNfNY+qQ3a3TjJ9eHYaweLnKoKfs8Hs/khnv
sA8fQeJ7+/KnnLwXin7FcX/f2BK8ASgeZnVCFMxU8Iww18Wv5QP5EMOypFZS
kCnQ1+LVmupwzQreJivE2pRxc9pD1VdlsC4O3VIu1A0vSSOF9e9W5yPIsjSc
LDZEaJ6W0OvkGUaG3PcErw5tig7oggoC0kbwIhU7OM96mp9MxndMcv8aOlpO
pqgh9+8JrBi2392J5xm14Nj9Z2PZc+5evP/3yQi/cAmwku/yCPmUdmSBvT2y
IsQAoGc11RTdJ9KFRew90VXL2FZtSIPh8jgTX5g05NBO0g98zWFJovI/n5RG
tEDdExp5fIcsOEafBWAOMyhpGFOOv0VFAiD1ajxZW3YkuF5BAUz3KHTbybPT
OZOfQINPwENluV7Lfr058SE+bRH6GV4MG7noD47356Ib6Hq5jkK3k44VbKo3
67uSEdBoHF7/n2OZKT4uwhXoleJ4d2w/MMMMkawrPqahFZSGBahXJ+sAryLL
uxiyo2hPYJTNZPMc/lf/M+BIj1DEQBbgv9cMMBnOpKjBr0jmJrDbRRuopWG8
X4ixYnroeVvuhvy+MAaLjCfGkawoNSOq76sQVo2POlIp1NOs9nEzUxFEgsDV
IY6loXMNfYzY+mucifhMlkQbFpCH5/u9Tmfy3Harf8Ddsmb5hRCHv7SNg5mh
F/CPSEeW76pcKeP2v0LxAYbG+HT9hCr3ucVbcJ8zdASSaZBCsvP++L95KyTi
JfJHJ1TTiePsaMDEnnCUZV8R64v6GycXos6jQ5I4t9JqECTbt2ZicCWijzZs
CtvsfHHrFo+ekG0eYPfBbDJ9NYVst3epHR9BT1M9OMzc7YrqQESgFNM8jOAL
0TlDItceAt+beu8Qu/H56zxBgfPPrFEekj+ymtePOh4f5n3U00RePjvBKmeT
s5/8rXGMQkhNlQ7lRlC4QkrF4b53exLzHUE9uREbMzOXVtKStPPNPm/g7xav
0yW/Yo94yoJ97uoF4MvkrVQaweaoC/nYfBmSMFcsPZOD3rPRWhoMEv1oZaZs
WRC7iJSrxx0rXxxRF71h8hEKEKHmT3CnNRe36RXVvqxL1fRoKLnDsGzwFi3o
4SYHN7OsDZEelAUL6P5zYVPoXx193PS5CNB/ISH+/+gsKmPMzLk6kDJCWbbL
unulnqzPBmgcdyvU1P4UkeLrMUXA+5/i4uU07EZAdX7RpT7yMu7ZtkQ0eylQ
GhcYGfOHbCopE7blyNI1+rsndfC/VKWFtaFhHVlQPHkiM6s4cNGT9LPEjMtg
C9/+mkauFedTgrCvFkkx0Gi/d3AZ5ZOlrDTuKdCYl0bL+QTmIwuwAiy0HBVj
4BG+WcK0YGyjBh8RJ6J+F35F2P0vdmSCeKPrTQ7IweJk6D4iXxmyP7wbDfeZ
0p19B8OTGlnShV47k6b21TZDkcRwVFEdnUWq8HsOfU62Aei5u43+JLsVO7Zy
sm7YbX+G0rpsfXGPnQ8x9gRNSae3q2gOjYqXONWY5K1J6dsvcCSRpVyIz04i
n6d+payDvyEz6Lga1vPuIGlUJbDuw7GJ5Jwn0HDyrXRko2nxeUQCzOE3iaDl
e27qbFGyzWcRlcuh84YAzXWt4NgppMzRjxdMDninzNHmJAkS6lLEfXMheshc
VZ0x3BAVWZrFseeatr5d7P009OU7XIHUwBKlzfKJNolwSmvC+FuTOChR93y3
15D4MpcqDzydaHOAU+fRjRviYhl18xizZ6ra6wO0feKgcard3vOTvkW/4dHh
M+H4xAl+G1nyB791vKRUAukt/r9sbfDPcOVj7pE3+UaINLOXsVgkR0jK1foV
qe7Kf3RCoa9r67DQf0JNKCC2lW9IgQ2xdOQ0359/sJiZO28M0IuKPZi88ekX
VgMhc9TSshMp1QyatrHTKCMVUNqn1MtWSKvYZTuPbJyWfSMvow1ynY4ekqlW
ltTtY/cSAzVf3U/5GtDUINypjtH+FEQQD5k+LboWZ8lzK6Iq9R0ZyXZ/dGzt
EKP+RfxRgpBl25Xv+Q+KCyRtW6wMROrzXkycnpd10Sdm0sIKDhwopOZb5SNh
b6uztm3bMGKtFSLmr3oFNzIPOnK4Z60hjnlENJZ9eJuOSyzcSPibhXpqHHTk
9f9z/vndunPPOaow/7MmcEdPeYxMEyMlYmfU93ZgKzJ8+jkV04xpSZnTpTE4
/kbRIofcDHmISzLdd6za2tweY7FkTvGRg7J3XEdYkP6tsHhySwQJ17ZbE2S8
/LFje4xSnXQw7lsUu3UUS3ZWAChospecfLs9JlH36NH2z7IN4PzIJppm/L/D
VbF0qP98hrObqvzuVvJT6fD7h10jG9ubiDBJS1oFR52CrctRQk0exYyG89VA
SmzbX/O8+aujM/LDQmKJfOb9zZ9ja6SWY+VWAmy/lcqv0B0Q0f4bnpEybbe7
p3/1UM+kKVwL0imOOfmDFWlrFo3JF4q0BrYjxawN3UrwaPZEq7bztxdL9AQn
XXVNj4RfWYhG/PQIMkGjrFmeGLDBv4oUzcm8KyWV1zPduTDtL9g5PBlCXeng
U4Ad6JiVOsUqyzQvi+8+EgPQu3eVCPVdGBVfTZ6FE9s1Ussz6SNXsOlDZ1v7
bE0MKwC8aCa4wWSbPMGav7G/fIEBqgNCjmIu2X3rUl18DFcNFGaHiW27vhrB
XiDCAjjn03IFIx74K93ZbvlYuW+jbW36RxjN/wnMqpZwhv37oh0Uc7TXX44G
uqTCS6s0wF1CXJR8N6k3/K2bnQ92jGIuqnaYdoIn73yVUPwkKt5ArhO8AMTZ
7VRcbnlWobQRJwiC2aIppwd6NOe4YtbwlEEctskQNg2hl25zU5/7772Oc5ok
eE4dH0ZhZ/XJg27eU4S4ywEBcG9QkYNkuezwb4MaCORefxqLco2zlU7lXvSJ
LbMk8AyHD2IsQ5KpTJwmT3Mef0KbosVfy9VKG34TJh2QAyiNwVkNtBWpllkj
TfXZSKHzO4XlOOK2WGKqu+5B7ipv5gaH5QaI6yD3ppL6DaF2rdg21xNYBU0b
lryhe8lWac6P6YTE3NUoGNj9fvVPajpIWnACZmnEteW1FDzOLYoAwYaD/qir
VhjW3XDd7TBGOj2tMUcAnxudcHgFEzAym/eeGT30RlDHKw/Liv/3pdV7rY4O
LlZPOi9bzoETk5fgBEznhxVW9vVPW13Z8YxbUlfusjZZfYOk9aoz/GkJlwrz
9UEvJin6Y808Z9A7f+N5GH2xWJSlvQfNbCpQDYsnBhUMBWzFbNSsDyKraEFS
n8MhmAJXHUDUOUQtTBw53HQhR4a9onuVi3rfYg4vLPEXcDmwMz//mSvjfIGM
58TjQa1MCKkmMIO5vKRY5uwAodRpnffgkAmLYswz4RMFnod/s3mmQPhtRk4W
1zxyTavy5U6G7XFEj3f8fDCV4tG1LkbxgzyQord3p+cxUaZP/T48kIhoBkCx
381CDtSIQmckNu//zWc3vJqpo3dG9p4OtMv6UjflWUlnvKOfVAPzfrXvDhdd
oCQ4qcI/J2Hcot8g+H3vv6E5P0srvdaeaBzG/ejltyDfkkcZaWtFyaL3yu18
7up0l6vt+XrYaE8GjIlxa24Hl90843rmWqKYBYOTrXs7h0CHiFzx0kFuCZqD
L6YwFbbOaPOKWmyOHwXQK4DPCfKMIpI+dcGJqMizIS8Zm7CedFsBEjySJ52+
I6M/zq3eXAVATAUgzYZZxkPlwNJ2TDS7DGfV6HW5qKGt/y4z59Gox0Ve4j2d
oEuLusBeqblW2WHt9S4iYMR2jY/yKVQPNZGfDfH2eSOL/X2P5g/xvpE0AqWD
ReRZb65XHp6q/Wf+Iih3hrWs90IxQnr6gONAxEJhGyjNITwOgLDMAMhERjyQ
/mkl69MCeAVRi7mewYsOk2tc0CuOXmCNg+nTCoWZosx+NprareqQ3Fuv+n8m
t9/yqXhg1NWd2OOJl/sKMr5KmfDKTmXWcz7qiMe4E3p+tD8ihCY3/VusHfoJ
wlV2UQ3A9ogdeFlmyfr5BHlyiLjUs+kECR3zgjNRrBLu9hBs+m5Q3baEZ9c9
kAyhwnlpMtdrAXQyXDc/Ez/WMGSXLFHEkBbGlU3gDnlHJeZj489GKAb1gkhm
haPmFp26XOzgxRlL4bKi2UcIAfTnEEz6f+Jof6Fje7uYWPUQC7vGd50vQF6h
+QlbZ/kPzDT34YsO0s9N36dzOEMmuuQxzj5EFqEEKTDbkpuCPWYsXuvrVyRI
P/rQmo54wQx7bwq207nl4IRziy0UlP/qCCKbVaZqYs7mQtc89LimtVXv5710
e7UVUTXpFUJnoIo46uN5uUyxAP5mB30oAblVhcxOotJ61gksP9gIqlCpcyHb
3+EeEM/Mso63f1Ty7VDvEin2nG6p7EF9umM4e68aOxn1BoJVdeuA1l4BlaCY
7+9BfDdGpIqMWpyPtBIGBV+BMsHOAtQKM2+JnUVHxyqS3Mo80lqL/khw08ot
0fCY4NYjL1zd5bqrqiXvSrpyBxaFB0SmkUce8/KG4LUearHmVPvLWdJFdpxL
UiTXgu5ijdSTwm68N2zPrLBg6lqoPvvYO/iKQ8YJirV1F6Q/KtKeELzui9Fj
Y4+AWJR3mdWg+U7Jyv/U/ZC5VPUp9wAeycRSLQ4BG9sy9achf7fyu84xCTsZ
3LdR6YMBDuwqESkCnSBB8cN6mUGCSiwbj+oib7ciGih7O/2LALIkyS7kI+po
vW3U2dtNfUDk6j/Ix6SONE+I2+cEFy7xplCQMhHCg5AysLt4fVsqvq2kzit3
9lG75L1UAjqZjkA3DWD4RC/llh1qoZIm85TrIkx+kumZA0Z7Cc4Iwvk2Uc6I
1R1JcnA9c17ZF5OM9wWP39Eo2lLHpCNgjEUIpRuqdc7p3jTzWteB9GXoWLYc
5ZvW9KqW2mVRYrB/jmFOB5ebmiO0q7MpW9o8qkLWqBMbyG/lOvu/BuZ68eIu
CFeP8KrnxU/8rfl9T4WwIWSXwXRj8ls8He9yhGBMv/ObUOhpTLY+w1Q6xlCN
X4VyzO0/UopZPmVbleeohSsAXWt8hpCiNSNNwZfb9Wzv+H793QJPfXcPfCjC
RkK/VrX5xVRjc8dQzMUfEgy4is8mjtY1BzwBlvtLD5plKlP5Szyd9SF4dEBX
aSYn3FkqLVYme7Qo0qguOUuR7+qCyK5VS85gmXjnebwYPeofx2myCIkLCza7
Acc+XY7jWC/H96XAlQatf+pRU45SaaitCo8DXuKwnlumxPC9Z7mzJA4U+Gmo
ULvsfKMhGNLLp7LaFH2R7exHGCcoqo8f/24d47y1jSM7AEAmfudcARMAFlOV
XXo2aZYmiRLPHXg8FLJ8L2bZkGgQu14i5/ZWlvxgCg6CivD8/+9wSSrn1V/C
bjjavPlz2KFQz+/+ldECC8qIXZyvKc4om0p0ydShoaiu2TMGJg9ZGG3uolz+
nBT1epR0QJZp5Muw4fmiIgTepqwMI3chq2G+MXIl6pJT5l+cW+HH0XqRGU3O
GXjQh9lCmdqXB2SbHkc3iMyDJRkZ+k5o4VL0O8DAntqsL9EcWZ0q/5y4619w
Z9K89Ak28pB1i3iE09Aa+lLn3kvlJ8i+GiyzPVfIY3vLEUtq2StpHUK0p43/
+xRWTQy+eCauoA2i9p5KGlmKsqunyeFqyAESUVTd9KZsZ5xZ8NoQH+e2vIdo
vAO6be+fAoy+10DfW0RzVdv2LUjtH6RtkCzREltOCTcjSNkAY3Fv6nJFtEi+
d4UZbPPWIwsfClMFA6s3b94wxZxrHz/NzMIElDcdh5vRuIyoaY/4iE2KeDAM
6phwIIGE/t5SnaFeonBGS4F+FOpMtTQOAx1knugXZ3LtWFPJr17LdL6wq4fY
UUBrHbDSkQC2Kka70Bawv0TG/Svr8I1JUBQiEXHjShJp3zSJcc+rqGqFiCAd
ok0ODNZoElsFF8a3pUD/6zNPPQj3VU93Ewd9768iTtFaTtdgA1xVaZ24trqI
Q2LulxxcaA+W9ong2Qz8KqqT3YIk1fYV/iYUdMB763P22oqBBBEXnwgjX0Rt
apqDVnLaTC3HYyqruJE6QqCVG2lPHlIYFy4VcxF07mib2sOeOtIi/O460gfM
DpAkYQP/v5j1B9GGqSYHKQaUO5hOwbJSLkjRPSjFxGWgnPo8Ye9ejb57WQHM
MOfNaXYQJKXhkpI1BrKJQq39BsHYOS9K2sFBCjI/XPIQD4F6AZsuk5jFG3pY
sgB88aeJcoJvyH2YLVhlUWXsSQJG0nPeyop3x1D+vFB8QZsOgzVWWiYKMbWn
1Vh/aqgd6mE/WBIRh7nrFZZc233qHO2Co13bcsqXlfmy3EIGhw8MG4LPPACv
446p0I7IL6NmXyijH7EiLkC3AMJm5jviGcDQGjHjYWNfwjKxmkWIFKKtnI7Q
7gln5AfVgmKrlCqqnwkD3ruITMrl5fd/Y6UiYxf7EBfd9HQwdujklEE2QP4a
HUpyPinVdFnpztDPCqPeGej0U313bSmYpREJNOx3x9R1fIJpQMmAuU0L7lfr
12tE6P1ce9n5RQYoTpMlkh4kDrtuvS/8Zeu+Kcu4ZF9PN+71xmwV6qJxhs0n
yomKu6OQu7/Ahpmau+6L5QSBd7dIJjDFL3lBnpnfZ1FN19s8EwuIMuj+36gy
aWZmVK9ELRS6Hi5IAs9wDvgYFPw0RSk/D0TJqSZK4Z4YZ3WXXZgu4VUS8fYF
luLyvaR/Qi5bPcR3xHUGL7dLgVnPm6ClIHlanqQdUE4dSZ7Wmyb1zYC3Zifl
qBS0RY8/aXWhZ8WpgfXhih1brDgL5TlmFkrd5vpyl0gG1uvrd4d99vo9abt0
Qp0LT0Ico/FbiSm3xo2cfIHvv9LaBZ9yhz7VIlZx8HUDzC6h07uzEvEvvuu4
p5xKkESOYy8Roi7SM6eV2N5SzKqzO1ROfDZLEGPNCoAdP36P/ha5wQpHZ0Tl
+J3dcCJy5VoOyjv15DqNa8CCmlsCJc9ehWW++VwoQeAuDuU9kqia0EW8M36f
1cCJYSNHE4/T8KkkcqSue6K3S0Jam/udYAK/mL44WN0Zf2ZaufgT1sw+W7wH
4n+jOgH6ruHJqOBi9KmoaTI1eGd+Vdq0bAscoSqs9BT9Xn7V16pMVojGdoeQ
wGr0BytTkTUn6RhufnsJplp2xtUdGK25V2Bt6zdjzNFy6q2e/z5oCsZT0vQd
QlQMD54wkEe5fUFwCYgiJMQFEEXQ9dH7wrcOtdNWZlYgT77IEx+vVjsz8yf0
ID9CIsqYKFaSyz44Kg3g89IMspcNqR2NRrN1PVBYwyseTu6nOVEaoUZjwyyh
lnNbRaATLVZs+4vCvr1q69yCOM//9N/1BED3Dolk7NiqaHmRXaB6bkcuxTow
Z3P0ocHxHFgYFxbE/cTVn5BURhvsjUdV4KnEC4W3pk315EBfO9ok8gBTy6AL
2H+HZjPFmY6TurKuwVTImeCSNi7joO8dtetDCEv1uGNDbkgDfM6qSHP1iyh2
sIf4L+DraM8gjBKB/nMXP+WRnHqCWsN16DaS+5Fa+8bVD2knrOZK/efyjk6U
7cA4LAKzKRWTeFURhhRViq1P7OYL32enXbLAEdHrv6Opd7gjn9RvRiJrSa9G
ZegvOpYRt/5VqUQr2q+aIHK8LEAMP+3SxWn06TNSf9GMLLOSFORDMGZwD8e2
436hZ0Ruc3umPEdSZk0MsvG2k5pKVWalycsdSoMZJaMR8zDvzLupTBC8UqK6
2C2Pj/b2nGQcrj1FI/mFVWU9cOibHnth/Jl0j/QYUEXkC0v3lR5ViZyKpGTu
W4WX3SqbpgXyc9lZelq+tp2XZT8WeqsD4PA30ijzwSH8/lMnd9YLl5/vT4Ez
yT30oMLF6w/WptJUm9Gpsh2s27JM+IcYryWXlcHY7tP6CEC83tpGmQ/Fwckf
tcol/LmaZCpfqgGUPiDRGqCMzzXq7qoEdmy0hWOO2JCaqVk26EpmzfFDs2OA
Q58iP0tCPdJE7iDs78Tw3zLWfDHVOdq2Wmnlm/w2G41y/v65EUeCDsPwpDvG
ZiPY0RTHNOvZrQ8+2JZ1ED/2TCfEFruL7uFQLZg/OobtGNpbGETDCTajCiSo
Nc6VjVNMaKjG0bRdNLgPVSGOd5z8IpybmYvngFrnEwGqZ0w59K0iUqENywbZ
4avFvCl9Bq/CKNqnmsFPaNRR/BVWkxrBCYseIWCfIEyeJQOqiOeDkAgsMJiy
wXMmXwIIyQgMVPcSjsnKY56n4ByGZpLqk53QwqkeAuXyNv3iVBdDrMuokcNv
BqaYgaCsoI7XD7X1AT1TpKW+uoPWq5jL9Xiivi7BWyF9gETwS+HZVvGPNeU+
IoymQAKxJqA+ya2H10UJ8m8Go055g7cdnrRqG0ECvEUg9LGkHKLvR1mRmcTw
NVSAektQqdpxXUyp7sP3IAOaeafNBfBvslyWv05CDKOT1YIKcnEczqlugNar
w6gMA1od1yyDKJDHO3ijBfuhb7/Q1sy4mVTCBQ8PFdEfIhyr1RNlJvtDwUaW
KOooOXT+zbE02hQQYbkr5npK36vKsEtwTZB6zDJlgxMZ/s0I/Xi3bwpZO76x
HhvvbwNGlm8t/5aoKluUwzRWoJhy2IHtx7yA/2yCs6YvSntsxAjlvQRaDP46
KkzaWfk4elvZNgx3z8HnZUoF9syC58jo8KJJPutzOkS7lbcJrRqeikyPw49Q
zXkESzIYy7g/71Amba9fp6Pb2OIBHQC0woRWjQp6Gf7sEzj5vosjcpeELCQU
ujT75jY1xakYPdtb2eVVCCI+6PvpHfza9Thv6KKiHMLqFPji5U0leL+ln5h+
nLbwB5LqghjPcJ3ASJcNHMA/RWRgmeGJWomAXMoXr2l76gfkaPkVWjJ7Ixt6
rGpBv5xmcrgIhkicnG7u0euFgqYY7GeTrb3IrPOBYA5GjTNgGdixLZHm6aFZ
RkqyvSr7gecigEjbFz/mj3+VFcLfoGaxsDz3PoY183GoXPCCgsoCFlJKsENA
JP6qfGXCFnDGbg3qMZdvt9BgcavjU5nRLJ2Urm3L/76o9bkTghYBVP0E/ysc
qE3LHB66GLm84rUGDHFmXCLZOdPByGf2ZKsY84TnPQuAf11tKj7oka7xyU7p
VwJBpBE3Vw0gOhLHaJjSEZ+aNEiR5/TGQWwnimqgebvbYpDIT2VQs1Hgom8x
i0ID+1tbtSws+leF5Rt4TKrsKH9uPUShhOGF/3q0AEf9XWVqaAbvFhddECa9
x2zhTe3dFMvb+maz5xLiwyoajERrUZId/C2DSmQg9ghaZFZOepH0oroH2aUS
vIU2V20r2jqEbAPuS5dg4eruSPh3a291V1vfs5MYhEpobxzkyVjoQ9DR0tQN
ddqGfASDJtJLuwDahEK32lGFPIJRVGdP9m/Z3PfZGeIQACasjTTiUnx1QnJy
vrBiLZJ5tD+W3TjrU+I0c2ubjdvgIz8RIBIabTVbA5aQvM29YVLWuWs9pqRN
HtXBdrRomu7v+O+qohvwt9+ibCt1tuZiuZqyfgk602W1tox23cgI6gR3GomS
xZ8ucSmbqR465snjJnlpP6pj5vFzi8CRflw7jcQf28MaUJV2iu8agZG1NGAK
g4eP2jLUih3ItoWHkeL6oPgV0oj5d4pUdfxjdfzHJagviknf+oxaLbebIh3o
AKEwhsngwgvVkqv0Wh+iWxPCOn4AQJY9b6Z8scwj3gJvHfI3XUmO1ZbJ2qlL
nkWdmxTcdhcAMefTqu+Ys8TBRIXnhKximS63yWBM0cR5h0yUZ5vAMv6LfLt+
uk9tv4U6451cE6JvIyt/ymWebgV3Q+2m0dn9XY6AMx+ujBiV5LGzTz/lk7p8
lcTbLgNX9eHlGAalc10i780lT0WFdK+Mdvkl2w3NAsPlnYlKPBUJEHZggHk/
7/VPBtcqQqKpUlCKDhfqGXMW53s+02ff7dt9Jhw+ohLZ4EUcQJSyd94ctfsB
02ktqIe593+TmIG4m+lxs/kR276kRxd1tZW7vCpxNQ+XYuLa+xkKYJ1/agmJ
3rmDlWXZPIYQiauOHhxcK0avS5c3FEX9jlHRK1FyN947vxWGzuDBjJ4Qdh30
AnF6PICQWGepUQ9QvkTnYSrBCcA67E+kYecZp8+MMEjbj3OXe85Up/L4E10h
p6A1gqY1onxW60O7LRQeg+tCSw09UeR+AbpLYNNnJSzkUrJBWd+ThyDoVM9k
zkMcB2lM7uS2JC5f3SNV5bT6Dwmwk5tCQ9a+D3zYfv2wfzJT8w/H+Ns5d3Ar
OShu068+rWNQWUIlRoQ0YYtnULA1fJDmb+hFFQUZtUmvjKgBY9NujcM5cG76
tq8dcxXdDIk2FDwbUjApixBeL0HMUxNP61pAHvcGOQE=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1J5Jzat9UXXY5UgAKgL8T0x3qguFjq/cpn6lN8ca/tAvxeGlOkEXio90XojN9UW3w/QVSVybFDghm1D/X4xsTfThxcos2ujznwOoVm9AzriTZkk7xaCl8nqlNo9eeHgJ9Rc1/NddK0DSLA6hMuS7Jjuuir2D68Yi4UEsBh6yXJbV48HDlRxBmTGR+vLWJzZnI3/qFifqhEDCZyrnB5Qx8HvY7f4geFnXMTx0vFBsSJye0UODinQq8uyEicFcQJwPnlN4mNpDzTkDOxHWXLNjQYUQ19dwp/w6lSDMacdQy0Hi0KKCgKRfagHJ2YiAslDTaGdjzsLcGv787s29s4rXBhDM0MRehiXg3dS66MZtWrh/PgY/mYQ8dKVeVRHoMKlUDJnwpPEOX28GU6IJ9AhRpcdg0iaoiEmEXc2L+FJqjHwTWBOxguACpMsURsKakY6eAbmtrCXtHLChmuUuPv1p6sM05Yl8VR2/j+fSOYJQrxy6nagAywcqeAubsljfxpSU0fUw9j+9xXMceGf70/tAV5rkgbP0+KLqgPdceSTi9Edoz+3rr4crg9WEVmhhX6YDeU4JFm75hpEO5RuFZGX158F+6w9sFGvpySGmYEJqL8gez7OWVMFNU2Z1oVn0f6eLRKRIF6N5goAmrTB9cKyUJ/j9RiBoiXxpztoBOYKg3LTX91DHfgDwpTqjYdK5lJpKUzghZLjA4NQa9JKoYQRG5eJO4mNzdLdcgB+G/upBRK+q16Sg0M5JOsVF2TwWwhVJkrUNPqBV+AVsHBQg18TfdCf"
`endif