// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jrCvTVFZX581fLy8NQragoffOoUXNqftPuhfQA32Q+6/sYigl4zU4CioypGf
oLTkLzvcWDw0NI8S7ZPNQPgy6FlM/g4WxfD02UnUJyg+TfeiSyDmKUPOhULp
uONuGq86RVgVBIfL/dl+9u+CvYvOmatjqLDtidmEOsxzW7lnc7uNLQ+saJLd
DCkCDlk1Ivn5Utb9YXZJC+l/YFySz9G4gkY2tGRNvgB0Lia+wAX65u4O/WAT
7BZzdM/t77cN669okGMmMLCEtMq7LItP5dIa1Yqz4NREmbOdrOg9qy1V3WRn
UAukxF/LzSAiav7uOMem3PXvP9TFCAI623/yBw1M3g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
az+y69ujWDBOr76C9gtcuktKrHESBGd2COkcfzzcujSz4dNUC5tF1RA32Yoj
ORFpIrQPD2823LEpMa0cuiSHdsMvdCTQs4x/rVJgVKsx0HUbAhNM4LRdhaRq
idBdNCjliheoQlnypFmgpFL9lGZf5SdaVxzdQydiZVkpK7YDAhd/kcdDmqvn
LgKdydWi1m5l3YYjVLVsZs6ypmJUB0UG11d01GPA7oQK8g+dALuxIyp+AdFJ
t0iaEWCIhBqQyLEFeKVowBpmNa1cWHaYFzV7RNNaJDek57o9+6i1wuOPA3rp
0BSVPxvYJxjbBXyyZ98OorTQPAxtQ242OfkLWyPj1A==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YZasXcdOLyT9cghVGtXbflx+pGgyYXA6H984gy+SoJYEHGTu8ltSFl8hvl24
WXhHBfXiGtfGhlOLb8MmIWGPicZFPCwhsgRSBmKsV6z+7TsQPs519UdVu30h
+2ojcHPzF9RSrhAlWkmfITZBY44jAp9uMkvxvFdAfvXARSlA4S4QhKU0gyge
zXpN2U6o5g5kvRRe6Zm+RiEZbxosPg1bcE32xaDDbdC9YoXjrubwEEoC2o/x
GCZ+MFduVmaSkywlKGS/3Ws/z6WW76qMWWh2ztcZ3kEYyWZb2xKlnQ6KWiYT
nrYMwAmMmBf22AwaQBt+5TgWgQBKLcB7Cu+j9Wmx5Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CNCmN5KXx67bBJfxwxIVD8e3emaZUkFpDbOTg9sXE3gsjsmLGF4n1Y5ZYdTS
a1KIjlWWs+WUTPlRhnWW22YatBegWFVkETdhJcJX60Lovgw0/m2PfOoZXS/R
WX6IssTP+YziTVBG6QmFWgnxB5HSLjU8Bgsx0LwzK/CPg2Gh9ybYbMeyd0Ga
CRCBLcPIUKNuU3GJowL4xoaWP12s9uIT8/WljWjxQ52OVTDH47D+HFpa6fMJ
vthAtNgpuNXPEtgHL/2uA1/2IFyu4LDpbqVj8RhOQN9A5CncX3nI3nJ7xe8R
NHX/yaAqQMz+eVM2yheMz2JLJk6I3pB07H4C8XYjhQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
U+CnYp40gVSxIFqneFOY36qTMboCEFbKAnJnycM7wtIXyKcsDz9cY0aCWz7K
lRAnZ9PpyP765ohAEIta27gD88nqR5sW+EKgvyudmq6XxFk8wBU/i/WT154H
hJm0Dq//Tb2KtVyPnprQ5FBcJF6ZksmM1R4xZFcGmJ3U9OdznmI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
tFHmVZFXtsasIWa1azGlIHBvfUD1ELgUEJIzRWBJ5kElXSXz8ipABYR/24lF
ixVVuhkWjPnmmYIhuFUxLjLUEbKp3b10ZPFspx9tki12yZHVyaaxMGYGaEc+
rE93eIbcufDzJrqiSm/wFAi+l+p+t+XLpcNz/qlUJRpK6EKsQS8o/TkVSY3v
fEzYlvcTLJDa6Wldclo9r9YAdgmD3T84q1IGgcU5hnBBGUMJuHO+RoTLmZ56
w12T1eQ+f48cIIypW6uZv+bnIEjLaRaO0t5CgpFav+W4n/9SJDcVaHJ0GZMk
qvCVMtXnZTiO2sJp/s17Y41wO7E7frIDok31liaWWT0T4eJ6xIpQlBDwkkpu
nWvaginGDhUvPs9fwaGWQGJA6IzlToDEuvTs50Cz4D1wN5F97R1F3ItZpK/5
waSPyemZ/IOW+mtKNe7ADEgHKFd07rp6mCKGglcrT5a5jXtmpWXfj8vIUrNA
T8iv4i45x6bCOd+xDXfCCG89Re8n2C+7


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aD3YYv1VNuoSbOWc+Jh5uBDdJSJSeL9UKKMqnv4dvxN5wyApkZhImpuHmwwM
+myLRpdhRIydCK1vHqRGJyF6ub3hQDPIhkgZoo0QzjhZ3ht3yXFpEXZ/AL/s
CYnIBcAoPezV7s6xHBDtm8oqFMtdD+HUtIG6CfGrataox+24i7M=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aA5wkAjkYPZqvrVqLdkBFXCJi/H02N4Foz+BbGDyF+u2eGou8W9hBpu7tZQc
xVaNj4lpJn/dBfVENDEJM6R3YO30QAF+7b9LsRe4mliQBtJNqIo08JbobVYq
H+AGZQ0/5EWpSNHZrhAiHknTmucm0BcZi2PKmkawbtWcQ7J6zo4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13040)
`pragma protect data_block
m43wOD2Rt8PA9W2e275NtzXXy31TMthQhsyVV8S8huZRY/Bfxcx+zjkWmRQO
zrKdX3Y/1oMESDLwnxSeX7Uzm+UrCmFTJvIU5NdB5qaHbZSHErVyQfSWfzcI
T+2iCuXw3bhgXjSYbbE1h19E4AFjMzzJBlsbbW/EU9CrPOStpJXmocXDzOpN
GzrCdf5bYggF6/LYy3+UIktZzoGoKXvEPmq3Z0WYWRA4LGZyRJOpJ8AqkCe1
B0jW+reqdy4vA+xSsw91lTkqKcveG4ggXWEd8DTh3BnvmTOUts2HgEi3ZrA8
SRHKIQhAxdq4hbordMqtFoPj8I3zNx+WIO85FLQmU17gqPiSiIWKh36dK5MO
lNBvxnSyfINso7nZPgZgUnbwOBQlQ8agB4MCQZghNaFNL6MVZg3HhqELrIm9
9LDO1qO4x2O1mx0ix952V28hi7VQbreswYrOutNMuqdqcWy4IJBaoLX5zBlR
SMlkwfJwprzkEmSbecJoc14J0P2Maj/++gEE8YdXKPfPd87K9i38RfITmK8m
oX0bMSB91GOyvTwWcygUWzBeisysRJh8X54Ow1WNREGwzhcGYOPFwfUhuVWz
n1uK2ckqh1T1yGRoGXJR+cctnp6MnyrjabSvyWlfHDydrpHK1/YY+BYFB9YL
BisAe9BLc6gZHa2c/c2bvk80f7y41HOZy6jB1SeMY/YnwL0Z2aKzMNE7LplB
6lM0LNgEXjcJCgZ0VRSUUU3VapLhi50kxCmkrnPMth++FDwVgGu4vmOYcXtj
tLPh8KMuP2NbbYhqLkfm3lUJST6sVPqrLjXGyxWRlmMRQMbDveoG3RIAwok2
9osY4NsXX2Ws8+qQGk4UdmODSPaNQfmwzzTb8hjMgxY2OlbGufJzfF9miis/
Hpd2MO/67cWkb37VLFMy7W1uiYgZnJ+etJ44ZyJ6ctQ3fuf7h2PXwFdYsywD
rHTqQEI2Weq7aGSJj9WS/BEqQUayJbS3KjwOucIiwvtBM+ZjNH8QLOh004sd
O1qkFKOCa3AxwMJgq+mH5DYtQxm1YkILBDux1dUy7sK6l5MHPktBjpUEXJ8l
lpMAe2ByPY+wFftSqgVzTe7vteCDvR17sYsG2GMi99jjnAljQryvxvA4EJkH
YgesEtjIzmkJPYpbILEKppIlKbG4a/iLjRh3EDbd0G9NxWmEXO1+C7SinHP3
dJGatCQV+9cc0Dz6QWAm4YJMjXh5KE/MlC7otGdyJG+5fSQmIWOC83EWzHfR
R15Asvfb9ROJzl8f524YV2NHifkx0FU/iXWVYtprC4z6SIlctArSvkaE9lTv
suVstLxLRl9bhOdNYeMeJBn2Tb4komCWd2M30vnG/qWORYvlw2OtAUbHPa1X
/T+k7cezqme/uSxPG98o9ywDp3xtb6tUNgcRFRkiYZ99kH3j/YAIXkCVCb+C
QZkWGKcmR9lXj9cmoKw6sZ24121QS8yzp+wYRD7NMTa+gKx21gnFX0Xk+0c1
fxkQ1wAulJ7HsuQM/kJvbfayiZfJKYtCey7ihGUR1/CzA5flNVi/SjT5hdNd
xWZb4RGYgqgoPHJqFf8Sc78CmwNJsFIuNQslHvSKXSfRgMGPmmn7nvlF3dQI
8MQNvVNr9Brtq2JCFCt2UOP2zyFNUbctGMhpfqGcoeIfW3cjukZfKyqZ/4X4
fiprC+29d2Fo75qbC8Bwy+zS3is2CjRbejzvpvdu6aKySB1BkxOLSEKXXwFH
X3x3uvPqEE0QjCM8IWYBgKFf8wBEvMXHQKJ4HxRhBA4TAa1FiokhQVI8P1+s
KgZTqTT5ytbFioHpG0vUXebV7VO01vbY12LMKHc1hKtPFU/oHjC91H3h5hhX
xck2zF4fu7sueX/eBmUS3wiI+iMxmxac6CQ223Pbug45U6+hs6ACHk6EkUjh
qXP/j84MbkM/LTUDgZEc4b25ZU0BgQENP0PSnTCD8b4b0t82X5OfsV5Ovss/
Sj5XwFBNnCX3oWUEOWq315RFiOCIJKT+PyzGB8DOvRzAMUeTaW9Wpr4nnF/t
hpykXiU5ZXA9c7EAhkIQ/ZEeS0Y5eb26ufN27XBsVuKSQiAeiKuRQyUDnK/Q
Yvp5w98RQPH3/Hsu+bTcaF3zSjLZJaS8JN3bX4Vamb+FI2aBSDny7ENmXO2y
T+asO6ewnmrVtEgCBOLXqABl4o71d4+NAsRjMXH1e/8x5AgONf88LGMOxw6n
6cycARlrh8Tm7IP6e5bcZZwmd0rxRE/38J/ioeJyVx05oCzCk8YWvKt4QvPk
tSgrVRyDkr97x8kSBxc5LWOTdyhCWlvigZbP8+4u0yWblXTLk4LxvIhx2qmv
KlERP67pUBdufnzGF7X5x+dZ5nPz9JsUcn7BB3FGJvF7vT0V8f2nI87PZ0vo
BRWeBDTFGcJ9Fp0pMo0NI+iBp9hAg/wOGyYCRPleYVlmFyouy2PnaN5N5yoy
T4Tz6AwcDz4XoJ7b3oDtyHj+cpdkym+os2VCUmxKbLc8CViufkk/Gx8Hnu+o
eIj1NZr7H8R4uBr0csC+W3l19+D5sZo6nmiu6GjqmfntkDeHZkz4LdRZzJ+c
qyx/x7WU3Ne2woZo/rUVqjM8cbYBkWrCBZ/SJf1f90/dJCiKjQYj5yOseC+e
XHEvpNVS9LiZD0LO0tRymGwVaK7EW1rLIF5hlk3HxQ1O0YYAy5QSSWTzkoXW
lMqLzvZuNOUOCPZnoZhiBq3ugljKAv/NJSk0X7zFABHRPSYLucjOzSfqegXW
dojqceXO2/Nv8u2GBBVwpmcLHPe3+kUdtFKiaHyA6Cjx42WYqavj/Hx91KlE
v2CZBTZfhxxTYUkDGGPyzx+x46cqdMp5ZTYnY6fxqX3x5mp/26aNylFcMfM7
DGy3BbrtAvxN6w+Uqhd7oULQK6YkSniUTIsWXL2a4YZcB7glTJSFkjkObpmq
R8/LdY8VA0zwjbHxpAAa+WaOztuvSzAJIO6xIbmi79pzU34g1UKzmkEyT4d1
lYi5zvISYED5DIaeJ9Irp05jVToRiYQxnt354NXgW6d52BVuy6BnKHusMtDg
tSffPSRbYPrAuWXEhFgy5ClMJgjXKZZJ1FynXbDXlUXrT/6kwI1wllZxDzJM
BfVH0RV2nM55MtJvTMYxpLwuRykYrpJV3VnMVDeeseEsUQ3byM/GwyF10Uxr
WfFLAVjoyJMV8rz0f6kzUt9ZqMHh2S1pFSYvbFGJDI1+/2g6Qf5a5rCGQlC5
aSaA4HdrSAodgO7iTUtXwNNm4GI+yTDNMuUznpvmh6ZlekN4VVNkD3sveNiA
EQpK7VLz6DpeKUTcN1J98Klfw7n90Tko55f1/LcTGd7S1rp2Yx5rAApH9Wly
43rv2gXK1AnFrVwI9mmsuA1yzZmRJgbZ2xRG3UcIiHA0M0AalZ0DOAbzHjiz
eD0Sx6wcbrh50GjR/YL63oTJ0o4HcRsJIiwrn0ywbTnomvJnsD7HXVQhmtMy
kILxFNNzoUiMWoEOb4Oce/sIxLmPxJeUSk2+s7Y8YIEsthvfyyDi4FpPEei+
2XbiMRlpYqZBu8wDayjGhdT38M111dpsMdPK6EqU/kCYWrR393N9+0lEihlQ
vLPnkbMw5Z5Tn8U+i1npBV/0drwXqX+4XhTaJX7w/k48RIkHYVDvTfSgxzWW
LKM9HbO5V03on2iFfKXTe2qEmR7kcAgzUV7/Iv2JoiXTrZ8AeZKkj2g4seG1
LP/TWgjNJL4/r8Xyk369EZfSzmFvUXSrnmvAm0YmR4tVeuAnAaIjOEw2BHto
fzJVDqycsEb2bPMhBHd+dVnZHLPFJIiVhYgZ2T5/nr3jOCdPdOCazb0s0/qo
584GScrm/NnxYrUbTRdHDK5GI+4ytCbUBJ9PQd5XFSAKW9dhKPjZM2TI7q1f
mykmrqJ/L8+hxLWSoeKvE5UTJvS5vx4gEmiU9alcchFP3XJuKcqxvpIV9tDY
q+dRkY/f9iHP+OED07L4uDHmbUrrlQ9hjG0SCSyCmrBjqg1fEOHU3B56dd5Z
ZENRw7J/Q70tr8oRBhr+bBiPuGX1pYusG8N9lhcPq7jRQs//cfFkYwhlq5Qo
DL/KtVynrKUIVI3h/dQAeSesArsc+BXJB6S8akS1HeNXd8N8mbVgNQeN6B/O
Ynm31qTc1OIMBCVeXHV/6vQQeAgEsza2Q7iOe7ACZjL6j5/56gx5p6p0O7lM
zo2tKIhoB0N3rtA5FHdVn5CE/6e9zxpZrY9j21igMQUvnP3t+LoaARjiYGHu
mfEiWJrZMvjrZUOkcYv5GfvN6CTexvlEWr9le4fQRonDxrGiA07T0RBFnnse
JgOm08KaGc3YCqXLuJkDTRA+YbYWO3X0gu6iPHSv63Bi+amk6pNP9S70/uX9
aCs30IDA/hnddIpzghKOpjPUdsa0CHg6YPytsSSiRPk+KxvxJNQTNha7R4Mi
SuYqO2Hbepw21X572bNhgVUoIjDgYKk2WLvQ6bFLrNsRhY7rO0Iwl5/Qhn6M
W/tZJGgYUCPmnqr9xnySagcgg6k+OsPyytYG/ulbbUtJ2X1e8IFlCTp7NEDB
vLNMFEhA9sMZlZiWgud+ylaVPYlAUYf3az+QPwSJt3ebINt0HJM2QJ/VVswi
yLVDPTCxfzaulsjHLRvey3mdrwmYywtv/Tesu0kkojeByc8YSclvOyqJ3ezS
MS15i0hWBvsRxBBhOEbBBLZ6Gq2VnKVEOccZo26BtIAPbAczqkWxco8r+Key
cLHmJYbonrJrEv8ONKbnwzhQN7rqFD7V0dXsamGVNfo/yBQKcjOx/tfAgy9i
sIPiKEvBRTc8iDYJsm/JxQAJKPQK3VlK6gRCBopLT0JzGpPxktJM9BBb5c0w
WbQ9s3xQFIzU6HETqtjsQmV0OXEr65RwNRsKWifsllPQFGXEIVEVoszcIRjz
1xFzVLWtkp7dl/RwVLePYSoMLfWeISKIt5jx9fhTr9K1wuQSff5fZ7na9fgO
GCiOJdW4DyJuY1WyNwN0txzr6NhD2uhLL7gHw41LE9V7OEnUib5NlYPegSMF
vyt+O5Z5fJqprTmLTU6by56n6EiOjdczvuQ50yDMO6fFJbp4vkUEHR5KqTXm
mKCb4V9NpJKtV+lRRk3SC8N3oAdDi9KLzM2TckeTDKuF+ith4I5gajmyJtAi
TMkgbP23mHoUGc7w/AgY1Ngx7T9/321sjRcRRub60N42W6/AMwhqi77H02yD
7IUpH+E7mhkZMXhxFpGj2xSX4prQiasVYfOo2opx7g0sWp5Xa2gOjNbu7Rwm
rbQaTFUBn/Lo2GyPiM/q+BBv9yjThKLlUN7CStk/AkWy+Q9QL7B5s6bJclEV
fKcf/M4/HBkSrHXSeo1/m5ZImWEVvqrm6v5jFXsu1YmusAk1Vs0SMAaTV9xi
6Lv5V46L1eUKM5DiUHGUT8Pe45alYRR8GWgXimDU35lmdiIQ+lLuJdMsLS9u
DYz0Z4rmIM0EMmm95SCbGZuNlLNnkiOcijJZVbvQbPkitIZMFuygyCrvqlHY
TjHqtxm5+X1SxHp/iR9Akz15Yhst7YJsY5S8D/ZRIxeD67LOk+FjnpVOcXe9
ohAzrhl6XUmug8IntUWaMvffTaX+CXizoG/2D/ZsqQpJ0eZlv7mlpbkLmNsu
4KseSPW9KG8yx4KewRSuzDeTGK7ZAm/sETn8/fza7p2ZrjnFrGrFrMyjnFkN
WgjRJI4cmrSiuJ4MJs5XUCDkVtDmzUY/Se6c8Ph5FBGtDFS5CVyBfUJw9P+C
4iY6bvaV/6YO44XdPIhyJOm+BWMUgObMeJ76z++egSvBSwgGZqBSKmskyDlo
DrXWY3Njcq0UoJKMklCLT8aXUtIL3fJU8EIjto6KlMAKPsXSwK853GlUe9oN
7FXF7+6vujR3XfXgWDQs9UNuVtcAL6pKR7j9QSgaYu/2rm4lGEwL/jgWxUXn
Y+idhduVWiUkZg4EwbopyDmrZVqahzyKeXlJppD9pFm5JML//OejsRcrVPML
suAWDzPZtZTq1e8YlRKx10r44J0UKpG2YmOUBcDUzl2ZqZ+qzIapqNhjXQIL
9nzVbBrWQMx/ufRnCzQVahlyxQDVxgx7qqgJTE1aixhem4/OdFgF2YI1A9Nu
K1W+FgU7fbZIo1yOQEYUecuzKCI/mrPHVFT/CPAAKtYQNB0Z7ba119wxkg7R
Bn718Hj86rBNC07tZHz73C9nfW2HNY1rri/hIiemmYD2Yvaul3hSqIpzMqEl
oek6kcmixfUa55qSkLIiY6ZYYj/FBaNcYMZ6Btb1jDX47hhFgoJ+wUjR9p2V
bNeC99T/FJdYE+EWo0LJjplBfd/BX65cwNxEIG9LUUj4hjG1rqUJLJbzeqhs
z5LtPD29N9AujIl1Fxmzbxj6kqDhuGYnpc9V5CYAUBJTobgjiliaI4yPZh/L
92Y/f+fqCCY7Y/ZpOGlhPC3rMY/mKT2UeS3dGTazKism8/lxfqFr0xDFgYW5
BSBc7hZ3GJHyfGIv73H7g56YPQyGiqJ1ApVO9Ea8kDmGLT+NH7YxLEnwXH9d
l9+ZMShrv+xtacX9MvMw19xIIRi4vyyBbIm6CmM4dv/EVeVfTW5lyuY3ZLxJ
baZ6XyAMVazygas0v8n9Whjz51bimMp5itsF2Hm5BBNShqVkGiPdS9ITkelf
bwq4lmWZ9OS40gheNdzq8q1n70srtHPsYYtE4DC8YIa3I2kjMaAmtrsLyUiB
IsKRm1y+6RUpYITSV6Wm0d/VcVX0ZDfvKnwbOI/IYCeDTEKLHuZeie+VSDzv
uw2P0ctmD2tgw9IJ09kN0vg0mYl6Xc4zRE6NKLtc0//Go8hQUhKS5misxaDi
zQJmMN1FNB548HblDEOaIhIoPIPno/xqEg+JYbTyZ1RdgZdtqsFQSABKH7b6
i5HRBy5uS76e4ugUa4BUKB1mZJajkainKxBPWrgLYvNz6AnziHvhksAu4cwV
cdMrtaAq1mRv67F2k804BU6IRSUwJWncarnIAWkrC/7gJWz9S7B07GqEliDr
KVlsKGVWcswcy181JCkikhzuRdP2KHa9fJ90J40Z3Wn8re6/edD9DOjTfZbf
TqtAIuL1dE6Y02wWnrSmN3FmEfSDRjPKipsWegVAaX4n0f0qh1XXgSH6UdFi
r/n4M4UoHTe12q6vVvvdp0gWb3yEa4I8fpn39MAIBSLV5KVby+ftO4VeRs9e
38+h0JoF9hDfbmAFlyuJdtwvg3cb575k2MMe3iCJO+tTusZr7jB+nQ/YyiPF
HFWritd/sxhYV2ggtuOIxvQ8wgG+g7emvP3dd4rC1C0IEKuw0S6rkrXyhI6s
zs85mb5Bt2HvYRF1AVU3vgST3KVnle2INcl8SY1MbIDZU4GK+AFAfPCJCDtD
Zt093GUJUQ3KSTVQoUTSGnTacrputSKH5Zf/cekc2o6YprTe2pC3V5PXonMS
z1r9tO6LgZNV+EehPJPvmtiJxMW4jgRZ7creiAJxN3FGlMeBv/JjTKJoARTC
+HEdcXujjqdGX+WzDZiUHZob4Me24rPqyXW+us3/G9TPKhc3Gnyu66jrPg9f
HQXL3y5UKbJf8Ll7zWrQTVVgraMZITOZy7xgqYazFOXpiSZEiWr88c5XWROu
ys5Ps7h80+ZfPesE4spWUx7byhcEpF6rsLznGsSTCLNF6pIrxRiQMcGn+bmw
SKuHLTPtBDDEpfCJ5uQJodAjB/3/QOFmW7/cikW7yqiHZ0r4edA29jSygN88
DrV7cEZNGMVXAOKWGG9SFpUfVFfk9UyfymTdNDI+6iwbl8LGZtg7kUXb7JCP
7lDw3ZgXIiPj2A54XuCaeRgdSpZH504Ahb5sxAXZvCCbmtledixI+dqHrSUb
xRtJeJOhtb7DRZD6kL5rWp8F9z2Fw6dKho+j7PevjngGZV+6k8c7OPQXH0xe
+3GlXq51HRdN/AwHgoBI3mJ8HGUCQ7p5Lxmd1p9Nt4AQ++fpO+ERBc2K5bEj
fz7TOCVeB0A9mzNteRLm+eN/gsef0grFKv/KLzzwVfv5isqb05DlDj4GRzcr
cn67QbpyjvStg/xip6Igvpp06ObdWyMEqdGOM80cHn/by48MynZsd9zdoDQD
0k2nXTLOxBBH3Tl7mQxsUKFBeXWmPatcneA81515Z4XMBm/7HzE5K0fRoMO9
yqBKn+UKGIQ9aXgxcIq5tw9ISZkQTajOTJuJ31+iV2qwc/rG2+pLMmyy01RU
Kuv6lEOAa/Q4aVvnTSs9aXY7Q9i/K7IljJHqV56lkvdUDLQ+pJz2LIDtEfGW
syW8YHhXeTOtBso6L2n1Pmcty039fnmEArfMzx7e0pnSFJw9T2BocAgy6vLN
isTwrq4ztD1LkSzsJTQMGScs/+dk8Eeq0bBbBdbDeT+OxXYXDIHy/kWMQkfN
1ZKxesBjbfQN2jItskiIMnZn509ED1Pu7fopcqKlfFeFeZgyy7U4BBtT54SX
MG1CksI81pepzo3SOHPh9yRbupLNBVkGRrIGIn/T9jf2A38pn2Q6yxWu1rBn
pYVaCtcyVgd+YrG72XzDWsVLZWxZ0BMZW1cTtCR4a3RoiSO+0/tVt52nKGsb
C/w1DDxcsfMgs21awnmQJsn9KWpuW4mtYUTUFajH666ypclRBBEqn945/syQ
v/CEXCfe4Wt4Hmxz3pp1cwvn7aVPAMl/b/uMH+TCRTaF7u9I4eUSxyT42DBQ
b9I3lGGEyhXqDCBjh1OcVrhfZkPV3TSvUE1HhYNH/uVNV0vmexBOa2mthwcW
73hJ1DQM9vm2OVGQr/dzJ+rYzGjYWq1atoZj6ej5ebA4ON+wFx4T9ZWzMziv
QlQBTav16P1A6FWwrx+yJVqQR+OpW2PySZGxZH18ufXZChCawYQsz17dle4E
CK32pmxMfyKBOcnbmOtD2A8z8baFc3dAJetCckbbiFZRP+1Tcbe/0PKHv/e5
u0UPADfQH49BkCrqTaReGKSs88BPd5AN1yQ/e+Ek9tJ96RxIwmglSFh9akk0
yYlU7SqdyxmO6XcISooS2dlP6OPsjAq4aFOB9LzjMYBOjSZY+PeegaMDeJAH
IaMA1il2h3VEKmDGxrAhLNEkXYSkwwl+4PnK+0yGAmNz1qSousWxH+yuM5ww
r09MQbi8Hm+krHeB2iZCYS3yOsYJSMlhUhGNOKOMIQV3ubC7q7q4STK44VW+
lhsF7sxvVcDrAGAD4ad/4efhfWSC0j1MTQaxB9pVgSUgM9uxxcJdbdl3eLj7
7LppzGSgKZSLHB8oOn22yDBxfsR5x1vmT1QN3MreD5/PNaP5DXRNoQk3c+0h
oaJTfaHRR6Mah5btAJR5u29+/nLiUb+fZhm9BirXbAkr9sjEmlqDr4rgmQQv
Pi7oNdXVt86qSL/iPYVcmUT6rttGjsX5D04bxq19GlDqIzRAmtIq15Vk8rS9
fcqnhOGLOQdvliSwD2U4iyTc77J6E0sVl07IiHi8jPIJSSeMaIH6SZ44U23Q
ojzPLkmm6wSL1YYjV7kC9PMTDfkB8b5SiLINdeR5DNSdGrjQaNY4a2s7E0Bo
nk9JyXURp22XOVVNfX67pRyStu4bKyzcns0EzTqYirWvJisUt1y34qVkf2bX
TLJMZfOl3Hy2fQyFw5qWiySZxre/kp55GuEkJc+00i/ZzJWXadcGD0ub8usw
Y1NPanKZZ6zkrcaScUXYA/xGIZtA90i32iLFoTXrtK4cZCBhGYAOGnoSzui7
lpcOa5XqzNIQyj7FFRYgWa/Cqr+MTlzDjkfy73YbJ/yXjvzgw065l+MQayPW
kLVxe62WVktWkAxPS81IRDXYomzpoinplm/0zOU0ew7iBoHhzJ/FLSFyQ6rp
WHbY786G25c4RcVORJ82BavpEPyY71NFACpWhWq8KE3Jqzh9aO37jpDSB8TI
Kub+qTVNXZ4xnOeNibbgKZ2uEkyN84lujw9P1pTjNaVVQbH5frL+cZBXjNR9
mj8jqHQMgUWl2Dda9z2AZ4v7Ht4KWlDhpoiuE0ROF3+43O3vcxBcl/JoAys6
AGUMXTmNbEzmihBFV/pAwyUZStN0RWZyxeAP5B2yLmwNKdLg3bzib7SGHdur
tc6kXLm+l+8C7bEw7rcoc8qiubLaLf8o5oJipVSa2c4zvH02a2hQrAOibN7t
xL1SuJlqJRpahrz0Ve+GmFMZGDFRidk0a8czkqNLr4b/V0emUtcEgp/qgQie
NwtNkyJAVL4RFoESY0X6qJ8ow0IXPLeuhT1fljQtRnPYAIIJl15Ar5tl/JQg
HnbX0RDAy6Y9SHWPvwxZMDd3OJTO86hSbrZZ/qMHZQt7RLJTRf+/6q1ZoDZ3
FxJow+QFoJq6iyFIg2cMqIWM5MhlIDqv/8aVnu5uAwu+wv+Bsi/Kd2X6VUZh
ZPFIZzhmj/MXAthBZtmCPk62DRsaNNYEWc5sDIHBLqGPRC/M1fCQr4jxxuSV
sk1SDkYP8wWbyY5bbg4auOP6TTrbfHGQIdVFvrwWXFL2mWjSM2ubk8oGltpo
Con4zeSA43maeY4r+5bixyfLBqCAiDwRfSLuiw4kP+CXoSqw2vPed1O7+sNO
dBaUTPR5wPgJAi1blD8L85uKfAaAddiUSnUpGSJXIXoBIPd4xYmTHdE+XQIZ
lgeCnuXMtDn6E3lQ0+FaYCChR1GIhNVhyg32w5oXfjuUSUvFnXa4+etUk4mU
PkXVs97XjmH9zCOsJd61WEKqdhaUwvwTrDkb5pPChhwe5SqsJwyi7Db9B0A3
oSwfvdU+++2fk0PqCaUM4fHc0yBWaiu+83X1btMFmHumGgnMKxUwGOfVHtXI
iKWsy2NP+tTciLy1lHYi2uiP5LW5MO5zxwbFHTcK+kzLonDUtxhQtCyQbqA5
72XQn0Ma2qtPwAPd8Xl8FDU0H+hLYzyCfIjnYsXeG7wxa4XXVGrTL2uS+3z9
JYZkX0uSOf8rpBlXDxqdFldbhmJQhazDqpeQNet2H1XzOLYDi3BJMPHhohPU
kKqKkNtSL/2SyURU45SlbyQaXeOJI+KmUMy/f0dISwVFuYUjDhCtfVga5TAu
/TisEAs7n5O7EpaX0PPRNd36uy34/nd7NAjoJmThPemKXrxEU08b7/p1baNY
txwOW0Iezh7A2qOpHFjdp1cBP3F3lbdsQvFrKufc6D51vwXZV5hxNLysNU3M
ObHeLVZ088FnrHQ98RtJU06oUVzeJfwSshFKZ8Am1n5HTcaJDWJQbWb9w5+M
SQ4mHetjT4ikxNENWhwb/NFXTUHYFkwbwuDcLccJJGzQJLbQTqkEwIl/OJ+e
laJEPaMNrL3rRHJ43qOf4m/DKMp2xmDWmnHGSAJiWb5TzvKtWYrImZXl8kfY
Syx0h0Qt1i3ly0pOBOT+bdrpnyj7fIqp78bFohy7q7aYrYkR4NNcG3fRw5hF
+Qw4TJTB3Iv6QzG5v8ylMot0V5KqPWdNySFAxmjyUhkUHoQhqT/aS9biP9yu
kC6Vd58CFqV8c4w27IUrEzzCvq9xJRS3UVbZkjWr6CC0uLIa2yXutcR5RN49
juR2H29McD47iVaNV6p/CqUuxndY97vyEw/FU1veOSBrBH4r2s01cCkBYjdQ
L/lobBjQlvhji/mLutQVqZt5Ty7XVxwGi3858G6ED6yczs7Doi4yX1fUMxDr
9XHG5i7Ge4HLekCTkhdXg4PLEjnqXxTyFKn1/dwf+UzHyogvPBLd5zyshWew
aTuio3oAR5F4DEb9ane/5zta707YRDVIAqsLF0y1y0gOtDJ8Eqkr1gnkoUb5
dSFwqKSEvjUZCnahPcZLVVxsDK77R012a4zJWk5vdHkpRbh34vJpVlEae4cG
htro2DcrkiWl5O+GrI65+lztlz2GTnbMSqoP0WUFbEusxSS3Dh21w/e4IwLD
XboYG6jCRvISMeH3gQQyCx7D6E++B+ppNNlPSpTv2E2H76zoLoCYGFcwOxex
qNbae0EA6oGGplKADpF6N8Ig7Zey26AdqoYsMdtmlcFd2dL6HHRZasF0Sv59
YKu1lv9CgDi28qAmq0Hc1QnB0m/aVZoSUQGhUIz6onqs0ysiOv1gJ1iPy0bG
KHINoFgHRlRtO1vWg1Rrcrb+JEkInTqiQKd+HMRKzXcA4SVKU0IK1FOhEP94
mDXrY7nfBtcU0ITDFgijCpulYNaX7UnhFFuQBcBCp+Ni9XJTQMWd2ul7KqEh
n7eGLY1ZpqEiBTki8OqBWlACDyftVe4IW3NnB82Mk1RrrN2wHOFHihUGPXG/
rlARhKSMbxhrGaJm1IRQB4TkcvABdypShY6/5hdLi5XNZ8cBK8+dbY2dfUnF
k8pN0oAE9zJ8irVtJmOO9Fn6eSjpf/RrXcoMJJHH5qmwT8PHQVQLky4t/iNJ
Suid2j4UA/MIblczxCoc/m/7PZTO5HKSZ/lr1yBPj/8d6Gogpbq9rYftVq5L
rWh1ZTYUh/A16RrjJ9xTWAHBE2ZULg/roHBIy99vWvwYv6wPudqOEMtVRMMU
lOFOk/hoARcADLKpuqEfso3xfkZuu6c5SCdOva5nMR3zI2gotX5S13kDprta
dETGPTp7RMG3EOmRQUDqEcjzVlkr1/KBkLY7P+fnxmpoXwXyFx5vtUa0Q1Vl
C80A4Dz3wLJXVp4QvIOKaqC2LFrWFK+0FVQDuLUnNmDAubJjL10Fo42WTsTN
zUJYzie1QtvALQe5h6dWl6tt6Atq2cCxy4epGddZAkE77thVdaZHY2yh4uBb
2k3sx/5vZo1+qfM8/cfHE2ImoVBw5ot5+6pkYNDX5epiQLLmSyqGo7WAf1Zi
1Ggk04pjIAPqLwBy36aA01twcXjMPURQfKwYXyt7X7XZO5nQBk7nKwjPxihY
7B1slNI1PiPnXYMay7X7QO+U7I5EPXna4WpZWWabJYQkqJCRuyf98By07kLc
cIMXjnfcxUS9+wzOJ0pDq7OVZ5TonMggKsDJ6cg+knG8nTCtoyHPyR5gOPfv
3l9a2y0eQ6GIZ4j8Opm4LGTk3IpgFxnz7mGr2d3YBMJAJ6Os8CoYlihfnCmP
zV0beU7xaJ1N/CpvdQ48bLtvZX0miEvk49FUThbBP3Lt73aQzNDRBWbcztZ0
GRnFV1TasWtlnU6RF76dJXfLJKCkqCDDuS62Y3JKVPd67LFWMbJgZ1KlpQ4x
fpne8XCsJRMHjIwypFBpCIx7VhSAYCgahEyJd1aySfNDQIJJXOLcRIQm2F46
LeZaXEMAHcaIR0N3Z6ZyiPdy09jcmXThWUL1OOG4zC2D/+VNb4s1qehtKsNS
3XF3+nBQzYEQhqibZH9NEnS+5PUYRveMIkJc5Ow0gahRuBkRADu5IoIL9vkM
x57W8B8dU1CAwCA37niVt5BOKZoDMjQPRoEKA7KWheeUuBJ2+z5IxevUeqDZ
OInMfQ6Id0G7rtJtgqsTAgPbHiopIxofLUFeJCTgb9FQwhtS559C/rlUOpVq
scK69yxqt5kp/33ShaIKdsMiVX1ZRnHbNwAVohaCe2e372CBYY2o+FAlZ9Hc
1DSvoe8jhyDlKusRc97dYaDrzG1J8jg9L3wUXHjuX50Ul43/gTqcdsQEH/cx
AjjJUBHz+8Afzh253crj+9megEz11tAbvQaxG6DKCghMd6IRZWKR6OdQdvIs
JtUg8N17PpVI9Uj1KwadybatWeaIXnTH5bDm4na1R7pLIBgLREIx1i34mnSh
R7HXi3BEFxoO/lOFb0mT3eJHFA6vx7JOUKVDBrjF15PdVQ7y25tLcW/s4eQI
W3QVrQl/7qgkIeRXW8c9nIqgsO/3Pg6jVlBkeZG5YIXM5FLkjYx6dAxjk2+M
arcn0hb+PkkukUTGQEu8+A49umouJ9prWIYHvfkJXSSvnF+sxjykdS9Y3G74
F+z7SpKlXrPwVRqB2FPX8HJABANRhRzCPx92g4nOyL5/YMWX4uXIBwA6wA4u
Z4QjoXTUXPDdfZr/rMLyW6YE5dFcD6OP9kkynzciCY+RtBacAcQEPLERdVLz
UJO5IaRcNw6cPqzQF3kUoqqX5X+INdBght98xJHYgjVvj59Z6hU9iI9g34Lb
EZKgvKDne4z1GiMRlsSE1RHlxy8iARWKPe12uDWf/+x6EOEKteVq4PunJBcB
2mSHx7N7qkxmZbT4Z+T2g2neFzrGyEGfu1kRRcUXff3uOkAXt5z30oBiw87Z
2Hk/hgww/V3T4p6nBZNpa8A1rLHbXPm/mW+YXYMCaSoBE0LMwndmg/+GMlcy
53VJ13q8jJkvqPYL2tTowmxIAV2I1FoIiAaeBc3blhOibVffhUB9nXWblJpY
cJNRbNzijNW7RNjLFXYS1v9nDK1VZAJWBwxLV9dK0A2wJXm+qr5Xg8eFH9sD
QK2h8XCA9C8xIeN+oFTshSjig/Sl5G8svZY2WoAWLi0tm6vaVJZ9BrXJAJJB
qydP7/9X0v3Fz6/wXaTEehvYX4YASBFj7BrQt339X0+tOSuERxhctQotB6DP
Imz7JtUthrD0AFus+78TPRJZpHY/wSQ1Rtmk9GBwIK5C4PiGeJzJanynLbix
tAmEijVYyB7mVAAHKkyFh4RsqkyJnxuXS9upxqgD0fedNJxAgnSRh8wdX3wd
Br+v9dCOVEQEm7YnX4aqTaMHpkuP3LUmAxTP5FPm6otPS/q4UJKALZRsj4VD
xHTEAN5n1IQ4U9ny6QwqOUys5DKM8FGejQLye6PLyrMVBZF3C4jRgQeS3fdf
t0efxaJTb1+ksKks6TgnaqAHAYQXFi8+xWSK/wWRRQ8uvsHJNbBRACcHqk8T
cMV8DBC4AogZKDfN+i+KKtk39wjuR99mCQDX6o9O1u7ipjETXWboNy8v7KPP
7eU3bGgWbshsWtIkPBtywG1PV96Ch8+aAoKv5tlAVN0p8xG3GN1DQ65RJTFs
VhEL+6Sur0yvu4ROdiQGF6bcpuX/GwgzmRQfunmarDPyQeAS9oCkgsxeqWjA
A52ZCqIQPxOg4vPO7ixBTZ5JGbO/Ug6Pk93Zpygq3XffQWF2YwazwQdHSuPU
75EZKp5OJfu77RxqY3qiHBxIiztSjdOqugAaelL1GWmndiUG0AopzvJymhGA
bV4CXCxw5L1X+cjQdZbNWHREXIvKln62gX4jn0BcGQZYJO42+sCY3aAMm0r5
KVVt0IXw3zP0qPU69M6MZ/Cv0d1Xi6gcSTNq7VvYdVrJswv3apPtslVkYb9O
vovJdX1csBrPiYt18NjJTr0AHcQtUM7VOvMaNrhSX8GJFuRqY1rUoAeFc+Sn
qj76cuMt+YHZ+v0Zazhzsn7i3dfPQVrOZzRvqaTVNZUsYJ2wLgM9Ry8Qiy+E
WICshU3SKFdbanyD/VFT6HhtRpLYCO0kPUVKzoKPTGjOuxfKcDaRfcYKPNuO
IOvTYoBQIgz0SEDBW4OyjwFeF6L1+gwy8NzSg8upBeH95I4g64ZN9P5Suvk6
fyMV3McSWtQZGJivouwOl8KfgyjwquSy2LE85wamNCUbQjkT1nlBx0MQXwL7
cjHqaBXhfCPYocvAFDUute6+uR2uNllWhvOEd19MEBuh7iyRoA04teYqtMF8
wio1GttKScWVtPgJ/rK9axDa/96rX4PHxNnXOVUHrNgkjlZXUuxprzS8bUyk
1SlRLj9xuFU+2h9bh76FS8Ak5UGlQMz+h8gRczmfeUMqM7du26UFUyJ5k2JN
yPTeqxODBthnxcVb9rEoPZk0SKXvqX3nybXMkANQEN8UN3HwKqYBMm3zG/Wu
+pGygllDv7BR6S+xU93cIE3D90NwbJZRjz68njoSCkYQZWvJyTGRn7alKyHR
RBB3yCKRp4W/Rq6peoKOoEkP6XkuyKxji6aykKrOno+3b5ln8mobl3KlyePv
s/jlXtE/2SqTqQ+Ba5/73ywdpshUuTZcsSGZQp+B8qy143jwA0M/mdGSLy8Q
88SnNcukfVRO7w6sFeSDKPpPI+HgjjIZmN5e3quOu2C/QB4sPUqhjvC8nzR8
U1Xdk4QelirEjnLq/0YC86J2EqfNpE8RgWcxULF0XoRDDXmC5sFzyoLzF2XF
Rp8X51yeFjHNJMubxdh88ohRmgjhaWmabn0lfTEluauimDCWU9ygfePkiElV
5Q6sXZKqT9mws9xuiWZ+8q/BFdQpvGPHzLFZYrxQpPD2iL0nhFunT9lbH6sG
C25phNoBBc0Zy3qOQWDBers9bXvXWpg5LygIHC/ylIM7R6TkU++ungfbvD1T
/w6lya63fN4stYQZqjEsAbMA7pVqggl/dffhQLpuk0CUcAuJxPS264yuLzHm
xORLAm8Wv2M0FjcQsy1ukudAVY6FJ0yj4H8UFj+F6mWgaGPf5pDvS1VTaaMG
SJZQunsUbbIfkg9vg06GrF5OmAS1mkvfdUXg/hiw8JXC/QRF8CXLd/B07bdw
W1PvZHzxXLs7N+clm9TCuAkvIcgC6QLoSFYKrLLxl/5ZS4umL32AzeHXSYXk
ROtms5GCdRAsr3/Tw4UT1w4cOKF/UwihDtBf8c4UD3gSw1tY9MV1ebsIVisw
LI5GGvXxZwhIZo7AUsa8/5ziZxhATYlEnRit8uNg9yJ7koiT9Z7F/UIBuXA0
KCDq2hGK6OkL/QStklAp9e6yQGr5sW/FTeIy7Oay5u5RCHvZC+H+l1Qmb+Pk
0ep1pxBkQe9kLCjMUvx9KecNf1oaOtHCz3/pMmDd09fpBX656wqhuf+KwBFV
I421rWGB1MA7gAY6KFC58baNn6SmTLvcJ2HX3g0loH/eQVf5NYWhY0KBTfej
NwDLxJj8Ul3t9SpXIpYEilVCyaKuZUibb29PqBHqB4t/QB6rFetI5PVWX5nr
GQRl7z6iQnPQl90Fz28JkDCItJWEJ9+4y/AP4+LTjAo6tIQ/485M+C1cq9Es
4FK2/O9eCBn76nkwb8qmG8b3ES7AQO/Z9Dzp6OduwlfX2VLSQPT5CqN3/v+A
IFFZ/72yrwJ3Cip3LWY6NBNFIuva0OUD4JKAyJWBOmOzM6eEL17PjY8D2cAv
FDIakLOe/K45Z2DFWYAahuzGQJX9RETRrfOdeflwTSGFMd3E2sPB1qsJb5C5
FDar5AUufI1UBvdkdHMWHl7XaHdMI6E4527dlLCPMTFllqr6lv1vBUKLq2fW
+Qgk9sKaF1v2LQU/TgmvoDRNxhc95CgV6WMco6Vqv4jocblH3vV3NaaWmVKL
3P3vBkIhdptvuuxu6yWKNUTixrZU7i4sUL76V+DQ1qP9FSIqkR/hoNAewRLs
3ae0W+qnlogiXDIhSU7H/lbCfO1+wB2IgeBy+mZ4rr6Rw17z7ZKBUBx8PjXS
11/DS76Tzv5sJoyejdKKepYUc2zsaD418Jz9hRnSv1miLhg30pPmB8S8Gpu4
ZWLUi5Xd5aRjDoDy85KrE6BixSCd2maVIYBJq8urjxqxUjA=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5MpeipSvxHwLPsefC8lOWvCsGO/Qz4JV1l+ewW5Dw3hBL4pRowG1kVn9vHqh7WVxqglgvl2TrptStl9eg9ffVMFT6tk3INAHy1FsnZAELyJsAZDRdIYXciDj4e14DfaFG/LvJr4gjn4oXtKCaEkbxXD7vr2sP84+kmTMBmo8LXvByOSt+FEfbTaFbW1HzPzu6eaCgoUm6cWhU6xcBWx+9LdbtzzSG4AxGtzfZHg9e+hDm6esheuFc/39WkiAKS+CO7NRjtb4J0h9R/Wt3O4mjtgL6DY1bM8ee4ICoyd0c/OS6sApB3GT+RyVnxkwIAGWotaIZu7EC4aLE43G6ikIM6THT0yl2/bc5VCHf8JOBJkG3Fsm90hpqmRM6uwnZrmfGfRW4kyNcxSWI+w6moexqAODJ94vu1+qHVnu4DqeVC7QXxSHBE8feRXQVPE5zYK/RPf5YkgdW7RkFrveNwIkr8gInsIfhblePttNFo3OSpAsHuwH4TgnbScuVT6OEixUjzmplNATk3cCh8PidY3u5BcVrjAG1/JZe5a/dk90plr0pVG/J7Vkm5IE6V6q82d2h5I2k4jynwahZ8MSjlu/HxqOxuxEJ41j81rqjtMNcGOn9Curo7ZWlwnrTG2nEZJaD5oc6IRUnt2iQu4dtpg4nnF2p/Sfyj/nlwC6IwDFB4fu2X+GUMK0MLHfJO9iB57sNHpm+mxOm4oq2m1SCxk6c8r6+DYEJfG7hQE6bhmhnEW1vB63RGsSSIsewH3CeN2JlqHMp35OmSqvD7CaCthcBzxhjQ"
`endif