// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
1HBhoycnWVUnuXQG7hMePhgWTVIafiqmXX1+KV6KRRC0Gr3v4xV4L8xCxQk1
yV1zpXUUzATkhMrgX8RAgoEpHn2fpr0n9zsKGR2UZV9v9BkTlRVDglLKOc6+
CsZXj0ZYve/wSNeuXJJBILceLIDOaU8cCOqIfYxLypaLY46nGZDMYrZntJ6H
EA6TLfKgkOVcFRn2krgG5cuONycYcvKJwoyESUtrmXaOJUo/mqKFbTMKyjYM
cq1hWZPY87nzlSgwAvI+/kUlzHNAKoCmQZeOtMff9kitizvkRgQ+BPWL/dC9
e9u/Po2CNDcqQwZybxPjOA6wMJGEfewYZXTbIPJlIw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KHAfZ8kMC+os48vUqLOslKTAdYHg66R+63pQ/6AE4UG1lc9sv+uw/qJoAbuX
QuykylEg5XySFTthnh/0+h1x9c4erw6vffdg+u6Ac6toSZZ1M57T4FTlMD8Z
QJZLbPG+4SAT2rISTRV066HsSJAbl4PW3vrtfyQsdVJqefAWykRwY+FpIK8m
bVGpZiRyGgdpDmTPkM+NDXcLp1m6u1aR+6oMNbC+QlnIouImONTMMLQYkO9Q
tQbfhOlf/kfIlRHN4Zfh/hKdyylpcjxGaUvp323ZMiQO5aZucxPlxq0F3w3t
0hoPRxjc2rRaqxM9Sj1O/aGoStsqFa2vqD/sgR+n3g==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mXQ0uDzOnfd1iXx6se/FN0yH1PVg62iccN/yo6vVPxYe6y39T6+33Xnbd9G8
KfPC0g3N+EwTrVuaaySbltzGnDbBjxmxLU7bH6if2q+m5kANTQ2vQpLQ/Uj9
f4x3SKsBfDCdHeQGPlyzw5Ajhe3/RtZqF5z9wM7k7Gl9mDSTM9vQ5HQ+/P/W
7RJuP7nSI7PQo6Z+TcNrkXl9n0jxpqmIhGF+VfAiiKW0u0Lgj3M/0pU6UkDf
Lf0cfC9EgvFYEKBDGLVtlSfh3oP+7kw+9CfI4S7KCYHpDW4w4pmx5jUu1ruc
a83olFfCcbufvj+iPOfN4RbhRZb6f3LxQpNNsOEOcQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ATyyBBnM1DmPAWkDmJY+29OZZFpd90Z6igt4nC+I+FEdv5oqP5R+qbbFUmDm
ciJuepkqqcqihfqS6E7+ruyhwydN4stKlSw1QallpF2hTtCHMsIs7w9xmm35
7kvg3niQ48lzxYoWDRHV77PpGFb/2AB2yK3ss+NvloFM6jTWBZSWoswfsYHS
76olKD2iV+5AAjigJG1Krl2w52JUenNqnnuoGQfeQzVxgPmdlqA+Xlq4EnDx
wifK/3qHPuCG7MEDTpPRLw4J2q2C2Dxzleg96YkOlmjZlOL6cNIyhpySd0zj
GKtZ2J0rMy8KcR1Kf+gNL5Se9K4nx00XNzWO/a38Dg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
M+EZECKJa4wRficykoCSS+axPvZFJ9qKFLo8kNm9hhmrTEKb8A7EZNKrlEGL
G2bOM7TzZCFmmpMEGI2oB65RD1x9DNlH4O9fHLRVtfMUR7vIquRmSFowfFhc
0zXRdHwfttQC+yCMAV7/LxCwK3eHGN9dr3AkLQ0ce7cZTpUb9CY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
idqtRG0i5+R2FA/FS4ab6Z402C2zzMRbIuLCoYaK557i+6ttQ2JOYIMu/HGB
OspMLLi/rfNSA6qCdp8VV2a2iCM8kgTJFHydSFKFMdDSny8AcS7Y/p6DOKJe
eXkFHiOtDt+LRnIM3RsngijIOOSXg7b9OVxSc9KdC9EiyeDsezX6h3kcd4+O
tELWPPirbLKgQXWjDBhX1rHB3ZrvyWVQD/tJGc5O9eA8lknxmWGrPPPXWzIj
d8ZQskbXioKS+QRZ3nx8rdqelOs30ZQVtOgfrViZlAx4XS0gcEpRsL4eZtxy
hpdJfkcJM0/VdG0OVNpXVmGG3EDUj18dqVEPe8Xk8bkSh8P776gUiFdNyArN
Q33uPC5XECdixYwCDgfEHK8zm6BQoGRi6PctONeKMEAp7bSSCEo/XONAO/WV
n1+v6MGQrB+UfmOu0RBx+ImSI2KtsTeGb6axI+jo1V8Bwclw1Lg3QvsHTo9K
s55jh65leoB+9pHZ6dO5fA1eIGpJ0KIA


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
e/5NaxikujqN8K5f4S5FT/e3wP30hSQlwGFs2m1ELjyd6OxYl1AUTTqxgtFb
D19QXAzkq2cwRTfBHOfQsUOUNBOQE3dWMVzDtV2iO8necFJ/Di9dISvQXaO+
WsXi4hhea9M/74S8FxTr49FJGfgSzy2s06oXhJubQSDhYMMIxNo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qQp4oom/VJ2uD7Kuo1mHat3PsTAUNY2CW96T1S9SOHEe02e890wKj7xMJnEL
aLHNTBVHUFFicF6SmLNoB6vOl3x655dp2skz0AJxTeVWsRKKeIngOJr1z18Z
6BM04WzBBhBvmPs2FknrR+4T78PwQag35VLle1aicolEAHH4OwY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1296)
`pragma protect data_block
OMxXcjTwyc4JqNk35uHwVF635izEec/zUWqau0o9UvlAn4K7ftsl8VGMx/da
6/mnzPPDqKiF8m93E9IHWkvhNNSPk3OBvCCoO4mbcuu0Z/mA8ReemqSEzLVi
1x/R+Oydb71OrDy0Vi8WNsuyOYPHl/Arce1y1HAVYJEYWn6Z+5tConpL04Yx
/r2g1aaonqG9iJ/DgpWGhtH7TutPrHuEakS6/AAm8cD5q/lss0/Xy7rA3gFG
X+vsr7IWvCTgE4tHTcHTY8t9SXhqODXEmL/nWltrF4XVwy8gwgo3BRczHWGx
nNwjDMJ+ZGG3pagIyl4k19p+kIfF5Xjkdn2AZEKEoap5LtVm3DFlxzCmO/3f
KFxNA2/5lVKSd9OwO52ZxFbslLY832irTjN+M5V7OI6ccZxNNNxRE2AKeVqn
rNOQscCpY3fb9nApzCU0oMANM2HA9n8euYHrHfaqcu7dbQQuw/CfvVT0DOYi
m1SkMA350HVBGqwyy6YDSK0Cx5IpY++mUHJH1I4AP8JmSUT15h5JpR5nRo79
uvB+6VdjVrgf0iutu/12SXtTH/U7hzmrUnJoDij67wx9MzyjC1GXz1lsZJ4W
8fUKthWfYw6Kh/0GA3+DZ74xFds5WMwidF6Gji+C/+l7HmrwSpD8r2PLTaAU
08+I7PKWkiKGnCUyztv2yjcz4nZVTX+xAkCypNyr9qVEV/7+sPgWZwW4qE13
8ad1d3nEvySNkWXe/waLvlR26L09xRI2pkrrbjS92kWdGxUjQGJzvAmFrtah
zf2o1cUNfMEyyxMyti4/U6UjQRuvRNjrRLv/kB+kR/oWmoQp2Vn60pceFCD+
DsSqPsQOuYwizC6LkWxcwazlBJEbHKV7gioNiC7ZcqqpnvLH/Na3Mn8nlhWU
8WTCIpoviYW/4NihspM7kNSgpoBmL0MRV+ojGwqGTa5UEVGp9ak0Sf/r2EZ/
qXezL9qu0mPIK5+x6LSut9mFyyYcG/HEjWy5H8zIR9wsNwAzn08pJnceW2SB
m7ugM421yDc2YToSFFpGhB3oKoIriuJkegMTeUKvRo1cCmZGf2rRtDz6K4CY
obeL1asGvyuYN+yiDTcOgRVx0PEiS57mu/bWo9BVPyKm7fwReZxR4tGyscB8
zorcv8yGNLD7DmzJh7kiyGxU6ZZ843jZ3IBD6LFyb4AuPcqt/bWbvvuGOBa+
sci1xZn9qsm20zQBdgtJWAAkb0lcEVzD9a6vMGOzVim02lltBKEDs5lxYhb/
8qzDnANGtobqu8d02JgS/BXFYl81NGdyZsjx+W04VFu+HgPO36KJ87FJxgBb
R4DRN5FNZc8ewlo17sCmFSdUdNQU4rroTUzGkEmlIYRz0QVhhzc9wDB+nSnA
Yjh6GvyVCaZIRzpTefouI7xaIEVUwK6rL7Yhsjmqs5cADLrEjR+1jGspcq3c
Gg6wFLllzxu4G/BPfz+mHb9RBh+KqUsfjf9SaoihqsHSvFqtBipy9VVewnnF
Bm8YVqQeYt+cfnkhvfcwP/JKj82fVy7zPC72VB3zUnS/U65v1rKLDME7wA5q
4Ei9VQsavYF6hs/7k78T8sxTv0ThVyf3LYk36rzTRq+ur7FyhrE05u/Q2CCZ
85lce3Y4D1lBpCHz28ek92wCSpyqbNOopoqktUsgS+aq8m4A8evw/QOawSAM
AjLZgNxvUQxL41UbD1vo2jF5ofwPbuJYYfvZEFg71Lw+NPpi

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqcALh4S+TYz6rI5B16Dz3FzZS0w/LM9d9SeIXfuzMwDi9cIfNvd5TBVwLRRwHrxE8ATBnAXSZu4o6DujnvtTiHpkA3AkpcXAoh+KaamzPT8KMPmr6NEGJzAmWMwYfDuV/HdeaMQpt/uAkNoBxkNGd3fBLnLYm5cVQ1MhwKIK6m7GShb+akcUPQilsmAOMkJs12ov77rRhvAuFYgjGzrXxhyebK9eVghpm1qYdC5Ph1Uf/u/ttbwNP6k6vxVSwsV7yI+G/FOZrm3Q3fbTVhfqJzzKFrBJuJWEUU4IfhBmDnRELJVRzEEonjBYOPQ6hx8bS45eQsyJVYVhu3NF5Ar4GzE0qD0DvXmHueAzezWUo8NDTFqjmoXcA2kiWMfeECZ97pT2yN0ajsqy/DUNnHIgs7ELvR0H+I1SyrVeoPaqx2cCTKBZ2YtB6bYSM0twycyAWLJO/aA2Bm0s+FEQ9HmYn2OZchBl+w3LfuiZ8Ndwihog+j2+7ljjlVMxWuydzRXEcb1FLUl2WBi1LZi/LkIfxT1wKVH3D8AsUFM2t6leYg7OP1LOVnVkAzoROrC24EwJCNh+3Zyqsbo/tmfAiRd5gFH/ymJhEDT+Ws23RFIrmyQTpNFmK3XuCCVsECi19e1EOPzoAoqlJJhhEs5eQ8sogpDErRfm2DcJ/0+EgKEtxntBoOIBtBHrb52R6imWoy/gdIyu2+YuvCQDhmRxjF2wAH7UwDknn2EFk5NtHP52T2TfiP5enPG5unlXeH5KHrLFP+8uJxsIyksV5sHw0Muojmp"
`endif