// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
o4EWDTt3PYToYatvUI4Guxv8f2AplkmfttlLnQWGj8pWxZqLLmabYCnmON/b
i5YDnYpVOElr0n4AAs28VLbyJpaNxonlyX0l6jBtHQ2q1D3An+B+DyiQ73oy
X2P9WTbIDj6+mPCwewLCZA8JbxNUbUqncI45nIt3AVjibkxeIRPnLf4FKFXY
JPg/RM2IMf/30BceZOOQKVXH2LsEYlnSkLI8mn8v9ZM+fi+toMYg5HXs/iQW
jgBmdVNMpUWBBmdR0j8mghMrIxlMvTep75bdasHmESibsWtq978s3X5A1wpT
jN3pOdW3V6wbbcilX0avRMyhjQx+VRDGjfqmz0aheQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fQRvq8ptnc6MM6K3jO+6DUgZAREkIUR+tIGLVMtCnKZsQrJcsjQIg/FTDqYH
KiQxpGIjf8Vl9tfCW2tcmKQlCHRpljwNkQGcen9NX4SUhygnEdaikPBDtUZF
Lxext2Z+5+okTD9kvHGaTCgA93GGqBWwLG3OTFQCFZxCFUNELwr+FFdnjy+X
EoM7XBkfS3nw6IPh0QTFmY5nOpXaE5nH2HLF5rtoYEXKvCbqJJliZkYJ8lkF
P0VvHd2d3cl4ychc0ONs1OF2KVd/rUIYhl8lbAbdEWyLIdiGriElHrDUMfbl
xaUbNMFgIeXiac8EXIEAkmDi2YC1V9ucY/LrDZYUZA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DxP+WzABgqiROO4jzaVa89G0wPmn0AxgyvXWy2aymRIY5d33jTXFj3c3fLmo
BO5hwF2pM9xgRMgPie6aiSk4V7KwjeKl2WVES/7SZmRzxi5Toq5nKLE+wGOG
5h4JFSwYeEq4XeBVt1h7CWES/xF3bnff8B1SgF+rJJ6t4CsfwGIrdx1Svc5X
n+rk2bDOQ3C1QBU5UPbZSSkaAK11U6J4KtOdtUEpVxrGBHyVScqb4SOYuk+G
DnnXA5BZifx08hEpVQeSOZO9RExmiTOMQ36j5eWNPQs7+qJQYj4+4BBLOBvD
Y/wrpZKn5nEyZFoXc7u6O0nKYtkqj18f+0NiIGKnBA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BcNv12sbSFUp4ZP7zynQ/P4+mUqDtk7JK/AUD14ifXU5p9ztfJequ1PI4yi2
ooSXXlgZo8dw4Dt9Bk6mbqzK0ZjOBTRcF7VXf8H8z1xzW2Bb1EaXBPQDjq0N
ENPJybeDrcEH0TidhFqZtuXWYbVWiqsrniEh2tv7lRTXxJ0gUYwEG9CQ4Jbh
LU00o+M94XkcPMhYKsKJ95cTg8i5INte1jxjX+hcQ31gsP4b3521YDvOJf0c
iSaZzQPrmkXEsc3cUbgnIqzwumvARksa7V/NR+8+fU2mbOyRoPCFnLoSfJ6j
MNHXXVHjK1eledBydGKt+6ceBA5u1Z7q+E+s7T9fUg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cdhM1HxhhYh6KDpyo6Iatd54Y6mhSZGhzsX3/UvpAleQp7wQV9aJ1yW5Sm3t
wnmGhHIFwTSYIaPzTeJKx6iiGEc0/OgOwprk+0VqqJ1I72tm2xWEYKAZpKHO
Yc6kK6LJaBbx9HIzXKvgUlaOYb8WlXOsEzU1nHB94ztCDdDWMhM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
nVcCFDbIRc3GR+xzSRR/LiCZtHSstu4zayt4vGmLwQkYus8Y7iL7FXKNsDh0
lrFOYImLvWO2dX37rKkxv4C2IV3ZLAn89AWWHIK7S2KOcSz122HsVd2PRv1h
f520n/NTq3DlIooZFRY0SX9RsvB4Gc1ykG+YUO70yNIlY/TQgkDa9gYH2xhb
tJr7JmOf/rXK3uzHrtsx9IhQs6jzp0FXI5GvaLlH8nzUT+6GRkzv8CJAu+Lt
gB1pbBd/ekvcnoaihzr6Zt7fcJ+R2gwCi+dy3imUignTZokp+xAEDQrANN69
vreT6WLpNw8HoXxaBrX+c+3lDctjZdG/GGGeR/aJ4RBSNvX5HqysRTr2FdWq
iaCFICSrXoYy5uc7zYe/jH5j+66haUG+mHeOLG7Ep49Kj3eZ38NWv9pl+tgY
9niSj2dNhU3zrteDp4t2Iw8YtDvjM5Dq7jM9SR39P9tC3ccm2zMvKyIHx+kA
ORKBATyBlhbYk8lg1vV2HTGscIYq8WaG


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XBMfAgc7HgOdN10RvBd4gAuwGuqoLWJcvH7Wzv5cs7feH1fFx0+/EBLrLVWf
GSj3+v+DpkYKvdTN6VdeYzzNUtPnqp8QjV6HM22DmrNyd2IoYxpSVg/UarR7
GyGbmP3JJmCw7v5pRo+46AQF89/CdRi4bgK7ft2AnIA7qOOpMNQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Q38dQ7aU20fm+//K+nLU4VRYm+rH0lkOUbNxdKdulzOLkvLiHeQXU0SJ9dZr
01Fj0gJvL+NCFsHMTJsj5Jb2pLEvnYouQ1QFAXtVfOwRz7yfSi2fPeDMtPdv
Oh3XclPoZczH7yu0entRvD2NmCK4OeZ6UtEitwmKKtGNdkS+Z2c=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 48800)
`pragma protect data_block
y5q3Vc+hOOdlQRDlY06wB8VXAHJ8WboK+ed1Ks2mIRVVFTJS9N2EPSxdBmU0
Z3q5zhW/G9abLfe4EV0ywKKXyeRy85l9ovENRUSAciOFC2XemP2RLI3ygH0A
EWuTVAAdHwYL9hFKfi/tux62pWTdQ3U90gARtGdggki3hi2y7noXx1IHv5DG
4PXpA/mCwvapvCqNhfZ2+PFIa1sQYQ9X5Xvw03VcXO0wzpGfvvep5AbP2Rmz
d2ukwzX50Uq+UHqQMCDXqYIp0XoWsD4Bm6lyTm69o770LiGVo7GCiXX+zgco
3neatQT2GXGFumLZIzxd/20EpFOBw6w7jnpU9HjsTJX0bY4A3rAjUVbi4Jrq
jpJ1xamKGKLFsSYRzZmIKYGo4H89imRVOTtSpIZCXb9ZGddpvQZ4axxCcQmT
R7WmWvw78EWxghVk1dtM4CHwh1Dxt/STmYa8Fuy1/X8sB/eQA1O6Naame/Ew
Qn8EyxF+AOFRVS7csClcDLTF1afTtHsga/p/Gh6GMbLoWy/S8ZgEFp48Lc+a
ntUj/25a/Fm3Vec/Ya3sk1rImM1uPN4qw2Yr6RcOLYAichQ19aZSkekx0prI
rtz/rwv9Z7BVc3wF0MIcUtkR8l//MoF7FN7g1BrUfEDR/gbfb1Y3YOanVZTg
FTt4aRbY/5tLq32tZp1K4ljofzJcQnIsu+Vwhhts/GmIVIImCjVo6EGI+rJ/
H7wE4gTQO0Lhm/rGMh3I441dlHNO97Md2/lUB3WABdRL4uQ4JUxjLBVZlGMz
t+MYwwNixm8NHIn8N2uw5biUjHYyZ6ubcRZj/6Fu8lpZTNEAowrYVIIWLfkT
qVqoKl9gNQUZxLPKhP+YuiRce43iavUNby2DWN8WzKlp8rsy6mAOwXan8nA7
e++lLe8ZbyokCjhY6TQsXcBJChL8zxLrZZCsMfoIOXB4inA8JEGWjtPq3svx
TI0tC2adDFknOgCPZcAWY+0b0rllFENfL+1ibtitjri6QZwME2cUyAJOmEVh
vPbMiXHSyUuoPlEcbmRC9gzvovz5TAguYkJHe2RmAtubLnBLySVLHVeRHeOy
KLrCx36hKuVRBkDitRd4hbK0j436ZQ7L4Q51v95lmxiFR1GpFyzh+5Wg5XlT
mEkHNJUkJYhbL1hiphNkI+g9PG5jNGUieDYgjGIYyyJSkJ6Zz3XPGDaDvvyl
OgXWeGVjCM2UYRq3GP7zNXv7C6Av1qWtH3aagfyrPgsiuIzatarhT8wD65Yh
V9TvZDuVD8DfFRsatMeGMvtlszxgdC+JwNgSR0QSgkEjFHGKE8RCl1YUMPUa
PvjWSpRsfS6XFaBNHo09Ma6QK9bAt++1lWc31TyzZ/3nCj2Yy1aYqy1MQFy6
33aYzAzVr+2kXjqbhL1+T4tZNT1XLrr8bNdqiXMSXC79TR3vE02mtoS5xffX
i73C76kBOnFyhCw1p0dTaiWUK6rpyWeRNpEGFgBOub7FJq82vNwbT72899hO
ILj7uFnFGst0d83FBMRdTsjOjMkMcxsMVBhw9e8LVwsDd0586dr0snVZanbq
ZcxN7D2ifu6QaRWn+1HyYuG3HgiLSgMd6d2HO8kG4RUjed/mJ+viaWnBUEqf
8Ue7BTszeg51DxV5EimlHJkXZzTKc2hrcSCHv6rOme8Z0E8kDDWe++W6mhXg
8ryqnFrkTRFg3mLc3GPL15+9cj6WIXKodooYbAzkkM0Bx1WgMP1fyUtlz/G8
xY9ne3jqYUwliZSikwnWOwRDB7qCDbRfFDOlK+KwXY7t7CcrkHv1ogdfhAf4
x7eOur+2QheMGE6m8sBmYc66XlTmPOZhZVlo6eVFQ1havsbwMOn5wAqBgXh2
yrtMCe+K7H9UmVKzBkaNCF9MXcL5mZZ1HuQzkrSdkMZI2fGSA2FbT5IetG/h
ZKeZMySnAJJUvYNEY8HPxe+HNCgV0kWYdpAitNBZvuIG1JkWUX0bfthJ+zqx
49xEN9UgzoVGWZ29TL2cFEiAMRz991vq/kWDxPm4CBviEH/IIslaRQKvSY0l
cMIezi2p0QRbZ13eJAfbQKCVNjKlumEhMkKxOIknhUhYK5AmABA6N53JsT4T
tLWe07wd5HLdpIZH3kv6NmgcKl9SNWMxJ4BChuaiP4MECiLNAtaPbcran1TR
fXRyMZKKb2vj9LE4ScxQs855ygog6GID31Pe9ANdwcuPzZJdzAMplSLHQqjO
KT86eBzjnWYgmCfvffbT6+B8PK1DJAv/32U8ibStW+3COCe0L76Thhz3vC0C
hxasFFROlglpFzF5orp5HsEKOdG0QqhxD/QKg22ZqvEoYPK6CycZApHq102U
egDv+IUgj1ZEEovgkEIWWVU93hdQK3Ccu9XO3BrbXuL5z8+7W8L1O9NN+pSO
jfbC7r9xQYu76iloULSo3jMXLmXQDgEmrwbtvxeouYMTLzKff9YfO/iIp+7+
CXuJUZE7a2qysFUkZUzHqLSR8SxxodUec6+4lbLRXbBVNPolCKueaY/nJgNX
mHl0IXHJ+57hdDaepe940NOvgIiVFLH4uahOe7Hewp2jnH4IGeOvMuIapLXC
RLL+0FPmRfAKIOzyVDia/btXZt4CbNTrWA4r+tOcRbq2qXZ09s1sbkRmldNP
aX69e7bdcXVjqGYtUyAqT3RSBxGTJjng7d+Nvgs0aLdSDqAM+LFz4u0QgvJW
vml+fs8mOrsCnMgmEnhADg1aWQA5ghWHHu/e6NQcboW/AzELsX6naUXZa0F1
xhNn3ZEb6egSH1LCKGU0pzBTohP0SVQxLfuK/lN3XZ+Hez0LSbXwSR3vr51K
ZYfWklkp+R21uPX5E2IFdbPHWdp4I1Tv6SBTLscUd7uCmbvT4ueagCCNMhbn
eUtHZMY3YfoFSE0e9ljj69iGfO/wlqCo/3e56WNCFfaniFtE9XBGCZ/flrdm
2luXoH8nqZrt8tThJqUwDrOFU+BRQDen5V1/oheARZLzx7/PvYO6ecmRVhs1
LcLnj2MXfxg9KOX+RbPkzuz2s+36U60lH/nxiiOCdsEVBN+ThXydYN1L3dT3
jTBgURhQ76wR3Jg+fs2Vlp74N4lHEUv8tblplaopMLGknDnIjBCTiLCPkR0s
cRh1+tvjq/2Bj7gKWq7Qy+RIWONt6JBSMRp9L3JTZKqC3Zi2WGJmyMaYdoXl
bFcVgfbWa0rNP6tRfqd0WGEpwvcSPnZ+q0lCmCSPTSR4KaYdoE18bdyzehbb
5ZS3tIOkpnYTVKcToboJ4ugap4d0Bp41yfl9gFcvrQp+JyldKdYqKtIm32Mj
BkWIDVKSenMqmjxx/sg361+5rXV4U3WkRQGR4ilfFo4TW9RV0DOZJbekDkuI
Kh4kNC3X7klcLBVEWh6pAq7GfVbGiwP5pfBVl2B9a2jdovoYDijOkXly9DfO
sTycHQQd3D8NBIuBnsu3ZZh+8IGwDyqdZWrJreJW8Nwb2d8lBG/dZHobaqfG
DP/Bz6o1FvBlvi1P/heXISnSwzxz9PD1NdVEieiEPVseOb4nslepfqoA/PLl
lQet/wtsUXesu2+47gusDoBl4qibz4KYT5GZYuJyB9qN4FqpWNpM8lRrz8nj
hiZS851G267GPnTzeNmEpETwGH4dT5KhxyxxDnO+Yx/VMT6nFtnbNEYRCyxz
3gMeGhmHjLZd1F7yK3Ee6VpVjrsZAyZ5EGgfOZ1gJ/7BvW/ZMTbS/muFzf5T
Wfg7MiP6aJ0N3OOfI5b4w0NKlZZcL2eIQwbLVnVKQPYAuvNimnJIOW+Xe9po
L1RZyhw2+48JaatSAKx2C2ORPgBKaxWNH71eLWFJvz+0AybTz6yPlfWcxlt2
uJtI6s58GV3pt0hufEgAqxX+HBv7WivVvUhtzQVMBNMp4JV7gEjpn5zcFtG5
La73xPzn/9iKGqFIk5BrJBrDxXyK775TDB/4zNBbmqIgulAJS2OfRmkD978l
T4jxv2XM67L0kDKavA9o4jgtbcum+a1gDSSKDvT9pEgEdqHYpQ7qNZsOUewN
XiyYx0M1G0mD5WK7UDMa4+BbayUFi/ztVC2Ww9gJZi3jRE3a864nftpVhQH3
+qpKIQcbTRbPlpAMNsO80RUcP2T8uDSIhCqY9ZGimEM/eadXZ5arvW7nuty1
2LrfVH9UXnBj5zgrRBU4/OSet07MfRESC8JTWsg+lBr2pOdFib/Ns11AQeyl
m86JZaXtF7wjQ7tr6NADIkC4UOwzvA0qjaOLPMTq1wE5omCl0Mq8vMdUbB9B
hlDjUfOUX6xAu1Xz3W3Wy45sys+0Q76wdmyIsy0JxnJjCBtvVrpEO9n31YU1
5/ErFxTpnlZvuKJSlBjQ+LhQPw3c3BsaK5cJz1fjMlgDnD7yqHtI2ZmxOngq
lf3X7Ico6mZ6+2jIHhYf49PNGx3Zv+sWAgax7iXH39yzhCiDU1J5fT175ifz
o5aFQacuzB1TZlYNDOrrqnMFvs7Zhqg5KkVHRIL+AAKq7ZdVFPn5jVezfU9a
MNgmWXrnh9YP64hSK4RNtHIsoi1f7n9mp1mUoaBLSCwI5wI1WjZJL64GBxWZ
pFl2IIfxEaz2SIf3APyj2cqATQlbIIOzWagsP+LbH9RO/Ul5Fr1KGVin+MU1
W4ocJq/1x9FquSKBqfgca8R7k0Q/Iz7TWsUZwCDN+xwa3jiQbnJ6XG71r3r9
K67grePL3EuRQBGNYtV3x55zROOaoyp36zkXGDL3/fh216ENZCmtt76XGPfA
+e6LuPGnSt+y3HvvIaIpD9iOa+3+iNtezAzWoZ0aER26MJzR6NouDmaKQHEY
9Mii2sgK4qwjZiTXgs+gaJzDbe2NI7ycLzGK0x8wD0Yf95IslKG8xUOBpTTb
0EwLUKKc/aO2BKxv1SwIXZcbPUX6qFU1u+T69/1su+tRkd8V1cccVH6M+y3t
XQquenCxfvHWrqEPfilqQmN0UNv/Y2qHCAWxwKcANuRb1SZve8lcbUBhKt5m
F5KG1TE030punk5U6hoqwA0joIMI3xii4DaRpkO5uKMb9L16f/U3qbu6n9t1
ilu9lSLIVH0osue0NOZZZLA3kLMsYbjU/jZgic7caX53mra0tmmAWv4zzPm4
Wmy95xbqSVMJMvMv3QJ1YO9z/IOJuurRgGy+P76IE3CYPScs+0tQtuDyKbWA
h66BqUi5ZUMQmDBGhdPJexzYHCV+KP7vRwnwr1giHWnCmwhB6zT3ti5R5vjd
Q0j/VleBxVlTUjECQan6gUZ1GvYttjLu8PJzfSLJUhvUL3i9QdTJmBtECNmr
Ljh5G0laQ3gRJNvgTKrQeNvsGFniAUa8CZqa3Uk6jDzd8qbDbkqODJodutc6
GR35dG+FGs7fCP6v9M8UCsUcvPRxqqaGOoTLVTZnWXZtACM/fCA5aF30KX5i
aB+D7Or3PpB1uHnVmcoqiuFNEuSW7JzRmB9ARAbHvbRSfwRmCwqHifqDXAkn
UlCnGLRmk1n2BnDe4DVWeOLq1JEu8feZrrAF8WuykV+hik5f45rcxFDRqJHu
9BrAbMI7/UZ0POmPVOpTiqWGqavwFWJ4VZ+LP1Wb3aQAljkM8pUkwxUEFtWR
FszpxXQ3Mlw2wCxPeILayL/xhXdK94MwIjQFtiSnxJoXnDFL2gAdC8LbP4Jx
aV/53CRBTemxXueBwHsTNivIPB0tkcyLM/BMI6sVu7lq2ynCQXKVzrYQN/VD
zGSGQWV0heBW/WbM9/gnKP84kfuLqu7XtQ3WFU1woehyhRcTLSiYWfpfbjap
WdBNjZSENw/aAO3Bi3v89CW5R5S1CLCxGDZHGATelpn4ye5e9UYV+gQAE969
E0Ny5846oxy6RO4J9luqZ+ZF4IKbcqcYjsG3QW23rc947iQASRW5rOlwIfkH
XhMzK5/9HUKxq/7Hj78z0QiBNdfB2qhnfPa+eYn1Y0cq67LxyygElDujgO1S
sUhAQMsWq9rBU3rlS+ZC2tXT15iN3v3udPrxwdSUQnNi4fEk+b1sg/toNtWY
+w4ljwFpc1AkxykHrFaj52crjhFXuSxzN0c6++R0wXVG8iQggLIEziDNrEQT
O4CONNuuwsXWju29CliqcH2Bd1IsaNi3JSn8TJD2HeAol4d/DmCwM93Sw4Ht
ss9weVZ+9b4unGKcD0RYiUxNAwomidf7Slp7vt3mM9zzBCK9lJHkxz7oCi9h
vvclQk40i/fN7FLWUY1QS4wz1J3CXgVQmacnA+1OUQOtonZNGswfiy4ixAhH
SwIQBpjqAej9H6JptMTAkiuBJj8hfSeNgay8vGVdAwavOoZeZ8Jro5HsiX7Z
93mHerg94WpNznYjoKQM28sUuRhaFApr8f+pta5LZ4GEp+aosTBrmzLi3xnE
lbub6b9AyZlQlXjjbnczs5KhLPAToxQO03wkClZe6te2fulEBdkpRggA5wwN
y+hLKgzV9/2IYNKa7OJ+YwSz2HaxQgh5nj+JGxtLCdmMFuFRWO8TI6NBMunx
N9QYMw1y4/A9tSxEbwydgodE7bfw3CAgOlEJP03flhbFMPH/AK4w9Fh0m7LB
5vrvlyZYs1N/LxVVSQFD/fA+Lb3US0QAruBNiplP97CF2P5SaFDO8yeVu2Mx
oqBQPmdt15LUWK+Y+Z2mvnp7OKNH2KF4KMn/rWWzuc3QOAWRaRqPl33jgUDA
/tkBUHTUtW8nOo+LrTguMADadXBA/hnhx+FzbkikNDPjBA5KS9hOl1r2G8Zb
fBBa9d1J9POr7LKf7JPMOmVWTrFVOpwzsKg8dbzF9yvOcmUfSP7dGZOcyCyN
KGKer4uwy6IyCT6NIvuDTYx+7fpIef5OEn/OrdqqUx3Ov0KAkPVTQsZgqU7e
ng1BwIxZ1EIESKBHYWV0CenldDdvVSwS7wIWum2VLiU98na3OJK7mqZ3FOpF
yOVdayeDLdQ+NxHsdhdS8nY1LM51sKfNLA37DftotajNDInVDCfhGdpr8PL7
RSUl91V36xHw88G0JvGZkxbKl5hqgCMNV6q5c51BjHJS+FFvI/1h8VhpXYPs
iOqvFaPd8lTliCMCyDAKXh/NS6JoBovZc+7uGztiNLkpefsZJ8Y+2R0VKgO5
E2QpNao/6LXG1JSZEIFISAG2AsNi4njBwYBIRda9iHJ9zWKjRX+wYdxQVX8j
k7aUARBqG63EYYXoYNVa3p/q1kftz30q6ABAztQd2HiOhxWmXQ5g1vVh1MNz
Mgvcyk4wDw6J0kfzzrFOMRdIhBnc+yRhGjmVod3qwe8+WPh013Ijeq3o2Qbv
qDDx1vH0pSh2qjdG9LMlviajiqCfwvG2746iDFgMPG7RGcHaqp3YkhrU5Srm
VVYgeLPIpEebo+bxd+LMxp/pB8UiZkbXjHF/9Wfp5QofnodrlZSsQDUmAPuV
/2ZD8fk2Z7433FYJO20VYIQByNf2hVaiNFHXX6dBHZaLhTOpFZTjDhuNBtkT
w7+gWZyeSZQkmdAfh5Zb6Xmkj38lYQjD+mtZNhu1hc4UHZosX+radgqT6AmT
NeYqDVwH01ejM8xDV73hLT/h5V0HIFSY56DNCmr2okRs92XocRPPwwzKlQeI
qqhomSVw7z4uw+zPQf7kQjFqydUG++iSMvmalirOFiXfxe0at9eli38i78pb
BrqZH6l6dUcrGQr38qFGK1wGcD7niTXHLyUAY71M2I2NxEdHs5VhAg/26YAT
/hIXAOQPjNTPty+IbmVi5FxmaHA308GI03RMaQybUmQi1SNeuM94dSkUvwyK
6ufvkNWSGX9d94YUUbCGXvY5wGjdMCS9g+ZKdDaTxHii1JAcpRZ5fOOPcMN6
/Ik0KfEN2rZUVYIaUqw33Kl5vtXYQSD7LJGba6evr8rMomhidipbS89ssllH
aFEcZqS9HMADeOS4ekqN+rAwXIqE8lS9mCwYVYwQr9VDU83zUjLKk4qGtQVT
8fkzDBnHBmzi3XNhQyTE2O8XsuEuM3K6ycIK0wx8atm9ViKEzEeI1EFMZdiP
TRLzJ7YGOAuQ+V5skrojeWscTC6V1jH17K+lBD6g2v/X7ib3Ls1ceZZdDM/T
NojEhxGvl/QqOQDRatxa9vIDufvtkZtZbwF1kcrdCNMpJqaZ/Jwtl6UYVnN3
Wsu8NXBy0TS+HjidCLR9rBVRkIXk3TbUr+nlf2DVNo7CLNhQodUmY3yz3iUO
ri+ERzH2QsYw2ykaI/9LPeGq9tUMgEoO+FXqQtpFk1PTO9pv3qjISreIRm4o
yIkcARvnIdTE6fP4SYqr9HCZSlidrFdjgRl4kD3YAvrCNKR1V5LRWx8cl4NY
acQxfud7/47Vy4BWznFSYoRpDXXjNlhoSgDYKWVQg0u/ZUZut6VCwM0/uOka
UyUS7Je4nlXntQXqp11CQ6hZ/JiWClxer5DBBMb6Jv/RvRpyy8OLamRVEPaW
p19SnLuNLrZ++uA1nP1toHTVbGFeLhFY8fULbNytEsvb44w01dhziuN2r/Tl
3LF1LbkUmJEW9CTjN3Z/JnQjOioXK4Tq51riFUFDNZ18RsTpU2H5k63Pfc7W
sXvB71zFilWElzQ8QJdmYpofYxhI37CvLvpsd739cGVo0Xqy0TwH8szMGLZa
sHWmzLHoBOE21xA9a4QHJZPqnTUXDOBOt4fVCKZUfKghK3gdMEULdCJITtUz
YxBQIetltHNnfJXzfXcLzBuJzmlnHN7QifaFJJTevpsAS75g8sKxooU2SgBb
z3qGmyxs7yOQbjlbYejUFqvWHUW/ps59RlyYjzGJ7PqFTZ0EGNn8/xpPwK8K
Qpd2weY/0NDbQws+dufKNuFLCtAXuLOGFZ0ZtX9MNdjebNpXdcWCYvSA+OG7
5BA86jNuI5IwSFwbvf0jzrx5RFn/REVCGkw2oMrSJ8ME0Xh8xGsBLKbXkKSy
+XKiRYflWXc9uZNCqFXuZS8CHhGRKTGBHD9bNmiXcCqyh0KSIWs+jLiE4x97
nYttcUZSp5ZqDCA5ggveg8DVOXsIFIHZ9vNAbWzgPS3YHgzxCdsoTzXkT3DT
6WQhvKUJVrTuEHtlChb1c213fnDNrcOniqVkNee610/S7C+MAszSzRvIk2ok
n0fyqaYa3eXawVfW+BIUFPMrDbX++ZNNyhdAbpwerc2tIKlznIc7fComZ7+s
p3ILD8ej4D3taUzbhieDEHHrg/rg6NciWILVA4nmBkRgdYY7kjDEeUCJoMDV
1QtUEGJRaITMHqgeKUVsHxaVbg/a3FHyDFCwRmF7c1/asfhHcjGh+UJ+8Vkf
aIvLeDgjojK/SoytjKasVeoovYOT9RQoaQeC1WzGyRngPfkeohQS/sKOMuwz
uvg2jhhxnaSGJi4d213C57PV6QLmKET2pkAyo7GPRSMNd129MpH+nbtoezvT
0BVdzc2IeX1cXwKH5i6LaCfLaQi3akO9/KoisLBMMWZs56QfboY3OnMuPRiF
JPp3dWpiPX/WpRtZvFhpG7+fAfoKbeds3qWHOzmgI/HTMVo/JlRCtMCGNx6B
1K9S8xvdjTbre5QX0116PzGl2A7UbPAYJIp+4Xd6rNmCjBAbT06r8jlzgD3c
+ipKa2BiWq4rUgCAeWl9mMUYg7hobWef0VxeJr8qaZcDJcZdRX6aS29ZH962
d6Prb0+m8cu126h584FqAyRs7tYiZztHQmXR5ROE3Rv6+kVTM0vSuvpl4lkV
LvtXeCTa+nUWI74xd7GkuHQaTbwhjrz+rVPMk+He3gamyVuwaqfTU3gAoCQJ
9Y2YORHEDDuwEUc7TLDgPsDJHJYCR82wF35YB75zOJgS3wbJqvSuhXFelgU5
Vba7ydzkifpV2owtCBDTwhF8IevdnETPvRJePNfs4yv1FJ3uMTwRHj0XjVS7
EZxvKxS96l1TsccDyEPVwCIpeBTkeiUUu18PxQ85hVOiaKVQQIO7clkwj2Zr
DmRtgQR/cSm8lNGkrkSyivFo2TulGVSE4QgZGTv9cbLzqKhpmntyEsKqIgyM
3NEoM+ZCEiVuzHirxRKYVbck0h5gNq0wTfBq0nQmLLFtPZRhergsoeaYXtds
DqT5osG7UiByhFmqWMhQK8SeXNvdeawQrt1YhlEcm0arSnqAqgJQarJu2H83
+h5wxodTOmStLwlYZurTgJNQ3ADoOpYSsVXPZHDDjwTe3ZynFQZpQsq7x0Nx
CxrlsGXyYSARZ2G8RlfIsoR3UuGA/jPcbygq8p3GytGP7sciWaKZ/X6F365L
ZknabIqbc8Mz/OWsbEt+/z4m/6ZWMP2B/Iotz4f80Wrl308EVdsYo9CpL4V8
zTEx5V4hbPGOsSGbEenZCdfx/yQwVG0lhCm8pbmCxdEow5t0wFfIWBZ3wH6Q
fvrcsv93veniDGKPt4GwDAw46zZFmde9AsqsO4kfN0W65/2a2CQo6QRoCaOI
OsDM0SxP3Tpep+v73X+YOHYQ18x4wy1F1pjwBk58RRdUTxhxv7R8ZJosPzir
9svmrrZ+XY7lgRnowbw6Z1NQmyT5j82ymEap+MqyUkVip33jwY3/JJNi6rTU
TS5UHd3++D5JfHEUkxGRVTV1CFWTSk1tTgr7U9PgiEoQdoGGaGSJn1IjMhUj
6WZE6GcoM9/6F4+ywD5/70Z5oXg8M17WikSVTY1exP1LmfKIKjiM0mw+3tZT
GKjIKC9L3F+sIyq38k7YCcSrSoazfM0fe+ynQrs35tGpglc8UY3siD24wM3U
bCdOUbgZXZhB+9CH5qayjHVWcpA4Osy5nOXmUuWFtLUER5lkQdCYstRyfyvA
v58HBu0h+cEHV3rzkqL/jmlYaUO0LyrV25FugwdoKdFmrlABX3l5cw/ZJkn6
zv8macxrVlkz7415LO/xZtOaq3QM7WFmUCbUsrWY3bhFCiWlTKIBzljdvmCv
p4nAg6mrHUhFv5Gao4FAG4oUXOugZJyuzyLLppOmvGinU9mZ51u2B1pd0Vp2
f9+CtMC0M28bMSro1Jm2vnGghEyyf0tlvLKzhErhvfmW5eU4I83ulZ7NkSzL
11Ww6XcqgMkLQyBAxSfkHz9aHW3NaUSklIHZqaleMKjPt9U14iNhwoCTzekn
3DRbnbawN/fs0MdXABRXCb7jI8WawT1qPCLtDHjuRQrcIXa0zG2PUsgjxLsP
7aJ2f5BTXvehF1nmgy6jMERJFKPSQ5JDysP1LRv6yiZJAxjt+6hGWLZCDo7W
87zZnKOBP+xvXHKDzb8E3BLngKQEPeE8uMakvPs84iLVTW1b+iP7pUD4rIdj
DMs/Nevoh+2RnFR/g9zkc0RihxfiQAlGNb437q/abcIDVGYRMfDQpLxyuoxp
qlJGq4BNlhqh9IYEq1G4SaIyI21zyVTS14m7FfkVoyn49y7tETZFt7W8m774
f17Z6RPG7nHeVoB8k9CL5s0n7OuxXMvNl6JkiBz8mRb2REtPRg/uhpsCo22t
w74ry/CyF4B1PRmRwlqCcqVSTiOAiLnYR386ONSVrZ5WHyic0Kex7zq3fu+N
ifbB4Bbgyw9hhJ7TPMWrh7ggazvIpC9LkRyLF8rxBdxS5LcHxelV44p1fAfb
+5814hfQk96++J/DUu8vw3izFZSp6OIIdvdpmRvt1VBjYbudBjQg9PSpNNki
GKQzCgjR544laIfyB/NsGqCEYd2+CmmKOdEf3KXUvhII+QlxwIDlGagUcZgo
kzr1JlCG7ysjs3yUPKz6ilNHMlhEj4YTnPmbu6BYvCOfJdOX6L45ryAgnGZ5
HY0ucxLiR2rFsTVR5SiyznKdYCUZi6HrOq6OFd05wA3kbrDLuYu/1CbZU5HM
mELvMl3oJup2mLWCTcmiK+8E5FGOHgOLJHLzToIWpI4d9bC4fBf2C4RdhzYF
1dRxXKqzXPFGoMeq8ksmr9tgz4dNjWMxmqhyX74EZsCVH2yOe9wD0OJMMpOT
zfz5qxtL4NNA9OR4lj19IPZIZFq6TpHEWtgTlSIOho8Isjm8hvqpKfHaGys3
IhFGoebi6CwdZLVebIIAkkj7aG3Zd/8CgGQuaCSMbJGVEIQsrcQWA35I7Xmx
gtb59CNFHBvhLVeLjm+Xh/5VMUafRhanbcQMM2peGa6w2aNaE3umYpGL6daS
4DH7hZISUEM/G4DV8G0gEcu5En5vfiFI8zWXb4l2RKw/L8IA0Ud+0FUtqHZo
DgUEUVhdrXGFe01Le5mjo+kkQbVIjLihRpxSoUlRZERzk/MeSlMktz012v9r
Odjz2FU5+cXyky2L4335KC+pci3jkeytzyyCWrNqkzMAF2JenhnaBFqNuVuh
hnTM2G8KZ2M9p1k3n49mqNWeaMuvyfUi15xlfuBaRxxFFmfl7cEibpk/d4do
pGYCedQf30B8unpz5oH31O5vAHvPohcuCopNw8d8sC77B5y0AxtCL9pd67W2
opmwsFXlcEbRvOJB0g5Dcp4acPaOrOUmwqER+H9x3YcKVnR033Z7QyNQzjJz
PvUXv41odOKF9aB31HgnVV82+HpR6v50uaTII88MurXIIjTPqhkR4C5iKNxb
3VHWAKVtkF7wIcwAfft0RFLqfl7Oy8bpWK62y3qP8mRWC6OAqQ45J+c2e0+P
8dA9nnHEBP+t3nLcBD4i+l+kJ5Dw4EYJ7zPzLznp9ca5zbZ0Ye4AvCsrCwlz
Qp0C8Z6MYTA9tzLbbujHgNDk3fuDbLMH4teMK8lPJiSjgfQvJ0Ez1F6UBqvQ
UO2PyVBVkVSWpM727xG/aG9uLxQtnGzPr7b7DRyIZWzOAAU10nj0AzitEB9B
cZwVJgGYYgkNr3bxaMrMt42v8ctU8Vv3uzbAekh9t/sHsKyRecIwBuO5VEYe
4STMQcfcMufQjma0s007MpkjIjo/qxYAw3cSPspoEzns6zjpCN0+3l8xZF7o
PtyFOtQgKJ6QzDeg1A174BbPwnhyLSI/eOY8jINBg1X7pCOx1fYglQvEZpUG
1QuOPIHIWDQYZ3QWqDgw3biiyGbxMtb9Awb+rhbNJyj/2D3pIHhTxQhltG7V
ijzvOd1BrPdG0qTQ9lnC6IrXGmlCHtMSWTCs2710LPgen2amSoPSs9zRrtff
gBb+1YCbuAmiNxCYQq3QvFNHHpgzaWmPjQRWRKh8Bbe2u73n0Bcj8n/YnEiV
wJM8UDPPGzgIz4bLQKLa+FFu4ZU3T9BEiz0PxqWx8Rw2A0drKZDYi9T6vvX4
UpH/p6Bz1gmNQJh4RWY1YReUbyggcPKUI6xqXOhvRkFnWqRAoZZSST69vXzU
cXzCG93RRaYECiui+lFhkOnGpnK8DP1kiceQd7k1nFAoXsGkh2dDow6Mctl0
IkUXx6n17OLiB44lfed28DYuj0kiQljgprYObj4RQYWqngqtP5g88Db8htld
enhaXk6OIXFaMv3F1Xk3kVzF/1dSvrMLDqTywLvbzSFj14E4PRAy5DBhAqXz
6Qyl6AvXMHhLSKyKaZ7W2VAEAuRMzzdF8VixiDJ7rGAU21EKMjM8bdSr4fFw
QNVn4Ecv9vTz8EgsY4P/6ZmqowOKRY32Q1vTt1n6BhUX/sIoRbFWbe65vWIw
/RK2bTEC5ldthUmhSdS8TQOkOXjTRpeKLJh+4H1rrN8rYo3u1m7SKDjg2eBG
aO9+dtQdnDM4VL6Qo5IM0662fxluXfBt4x+18wSV05n4ywdtjKYpaNfiE80v
Fy88tuk5kfJa8wg2vsCMO6hwet+7d6a6P/1MKNcJh9aVopf6O1+3/F6Opz2X
EGaMVZelFdNoNTZ5S/a7nDfXTQB4s74pY1bNELg3mTjGTVRDgnzYZx8xxvG0
KTmHe3BbBVjobq2nOin1RPUSozk2CPcp5OrvXup13M0pTzgUllv8EElzgxlO
Y9SVwcdII8vyebqwx/351+mClQELaI/rOG0wkQccUi9jO/ApGAcl/7GHsEbb
XJHOz6OnCDzS6ZFNlY6SldcgijXkJ7px5YPZvtBVq01s+Fm93G3YLhvJBQ9F
VQeDnVlnDAnO8rLgJw/njZKecdQNxOnqioRzsLCsNC1rQSwFCnDPJlKqHHXQ
2MMCsHfAJYj6cwmF1M/uzINOF6SLnIIm4dr14/70TKQkZm761VAjxfWBkQ9m
t4GV7ZmXsyBiPKEGXa7QNIUJ4zdsIGktoNhSNLCwqbxCM8QyVwZgwhAcIUY2
yyMS/NoUSgQCZtDFRdeoCdwqzh+OdVHGgy7JINO5bySLlDY/ax96WsIB2rj1
4aKvi0zWjf0df/DyY3VL8jesSdn3JvtRCBO3uKCurE7egT4Deq/rRJrx5gaK
NhsfrwOY0AhSJ2uGj4Y/ToMWH+Z9UTfYNUVS4j8akMBPqwW2lwiVtZA9zFHx
ain75ytCbAVQYl6sNqaUgDZzSLv7u47WqmbuDfpav/Y216bQMNg2aVSGtEv9
0Y9lCngJC/xExSSEm2VgqMrMywMfvY8Z9i18I9tLiERhxty1VwSasbnjG/1l
Q1OEylNRJ2RrQwRpPYBeqDUmWAixdlCIKTfKDlhoNZ6FU8R5hGujcJuVj5f4
BX1K4WqxiNQqHkJ+KscuIOj6IUjccKcWd3jIz0eAc32C7kdaARoE5Sh1LkYK
D/M6wNXCcuzP1zvo6STKGzoTbI4d8de0it9fK3ZmNopAeOB5ZKLEySRjYA9n
vDCTc5IBYUM1JJR2FFt/kzvsem3+2e3FHtQVObv4wJPSWAoGK7dRpFMoxo8A
2kAe4Dm/XQLwQThG91HvOJPWADtdXY83GqHIHJS+V7KSWCC2JHyYiUcaBlNo
gariYfMsxMCZq+ANdsPCTHcZe4//BRtqC+7GLmtYDr4T59QkZbRvN60iCknG
vIk8QRhG3AsCKrm9RxQp/T5jIDda7xWccbgJCt5BXR5a9xgKKU2snVk8YUqt
20qGUj5ui+sfKnCe87N+sGHqkswBeu5XPrpSlLklJO2A4SewpLwC0oXjygg8
4ThhFd1cc3OJF0FuoAzYsFWZmrYI81ltMHoISbe89UJznh53WYET9ZSDIgiw
+slsVS6N6v510+Gf0vVBJFF3LvEuRkR8YvD3BfpMvSTgtvrkzKGy9wP+wiUR
7mS9V9HC6mB0qivv47CHkxDTYep9gK9fw2fuoK2yaxPyIZ3LWLU1OWjzxKPC
kWgWUROZSpYyEhQTtQezdlfYE7cwHl3cFZyt16Iw1AAhG0ffP6AOO+ftUNtk
PjEvBzTXzcN7TdJvT5c0ceXBVIOY/IXADdA3E6JSgQRwk22uJjjF+GNppiS5
GKLuOoBXXX4QVJZdBq8AQCh3WtVUpJPZ1HcOJKMr/WAiEBDkNh3LG66st3lL
R3BVX8yma9c16WpPHkS4uTcnEJlEQKqlEMybJGEf6Ge2NNaKtuSwJenLeOy4
rBLvu8nqexLJGwXwOHKBrKnsHWnPdn3syDdM7VlSwS2rgQUBechMXhmCesUy
vglqyCiYvu5sljuxfc8rv4iTol7APZwf9mfc8VMaRKc08SyTJQXxvLujaieu
qyJ+K6JYYqV5h3xtC6Ab9CnLnPdreDvwx902HvI5PS2F1/b80MRbK6BdAV2b
Ssyv6z1sBFooMTk/D+bU9ewpKlbAxE6t6xXZNflVLUP7+WZfQjinh8nTDwXy
Wgbw0s4kawe2qp/Tz6nMHGxdag9OffSje/Jh4igeXV1vm5lY8aRd4ntze38Z
nYotszPIyhuVVBmQHE4yzJliQOFwV0OXlQipfFkQHbkfKAhuiqM5OF327EBA
klauhQeljN0ZflRCu0go/9aq2hCeiuqswO6ehW5oUaojo1hpZbMFywn9xX0Y
MxNDPmwzPzPhYoGTGt4Jksr6HkiEmooPBHC2zFZV1Qa4y5+saAvO0nUAX/cy
QJZD14x3CJ3IfwO4sXCKOlr0JJZFEAuWzePKjUOQxn7qGtE8O7iccC/z5735
2YRZZc5apUt9LgM3tU9t8l/Gz4Q6/+UJg9FJtm2wLGypfTPPiM/IhuN7uZqT
JV149pGE6vvWZG/bG0VfTTLrlx7tEQ17U6ynWTaAn7k/s8P3m8K5+nZ7Iwbn
WiR+97tXN31bLoWlBLUufcUTK9fp8zWGdZtYDY8aaSIslZebPfNdsMT3OvFf
DG77MvdK3x4d88ETesO8hgS5RZtXlNJND+HSJ+dlBrneiwc7bK2aZF0N2ZeM
7XTEnRiKapkoR0rWGm7WCHame1Xb5WutKcT1mtRyl3BkwN9khgEhe/rsiBup
oBsXuzjDoIudDHqZ8+opR9OeBSVYlRJcgsr+NjHuY/Vfc1DFSQDLhFiIYC0t
3AnEhwTxbIAL3IHahpbvWtCuco/cHiUVGGP7p3qC3DS2xilZojVfyxlH06+T
C5C1FaOJuBIcx8qjrOSXC4kMASIxa1Phnraq9l45h9EjM9rQlAT4lKeBxprO
CO/aZ82PwtXheTJg9Vv1xLqh5BTXltq6ptFVrFUlqCud2Ybr2m4RiKLYAaO7
QPeUIOE1Yc8AdhrpcQj9B2iXPoN+VvWgrpF6JndNabJya8/mlSUgZbPZTaz5
Hd+I6fGu49kVBqyGq5VGEmZ91oNIHpRjEiee7WnnpvAlQl5apw4paEfh/8Ul
bGt+DI1D9tu3BAYM3d7wDG6E/lW6YSFWhlGhxBc0Dr7gNWGZSNFBiMzJAkkm
XWzcXZfErOWRSk/3iGFzlCWWXB1rrCh3GlxoM2Y1g2LlTyL5B6KZvwrbf+Z1
qMPqTqrFOPrH5TyOwzeQeu/IQ8VAW3zKkwpAlGC9MmgZAy7wrJscuvKSsFw3
MGG6oFul0KtXU8z3Jpnqgwjkuukwi4wTFH4INyXAqsH90ucywefSZtkdZhvq
sRn43BSzhWPXYKc8ZoQ21eikVK5PPXYoPZrwnfTGXgo3/i1kTP2nZmKdZzDO
56xJLtbtFH2w9ykDI9D1K6qsytSBMqU7tb9pUozjoA6SH0cQX7HeNgovcoGE
IYmvZ2BghfWRgVWpZKQnhYzrZuFY5xooZ2W6cIYwUUGPvrQhb+Xhj47m76yT
2dVEmTMsj5H530EG/SEFYcVUmiCGMPf+x8qkfz7An1YYQTiLizlMYtiYfyIo
8DLFykA6vhznrpILc75RWxhdBSHRk4494Pwv2fRHFFmGIlh2NKIbC4Q5vvyA
VzcIczsaR1G+rkzMYylShzDyQhms+QWyAz/bs3q+QakrMbUQi0KJdyacKdiJ
m1GZHdtUHy6EkBGO3de0W61FjsjwRF5ZHerANYK/Vfz29AacJmfYEwNazJmh
xRMvkrTMnCuk2zeElzRD0nkVGAN84kakmw9Wtyr274l3NiLHnpNAsPUCjihv
hHk9M9DZab/NeyFSyH4axDYoX44SB2YDGFrAdRvuQs8Ht8/tayZ3Kubp7gYU
Ej4fC0kBWl7396/UTT7iPXTJD7zUpExo6fh92q4bU8AYhgZU20HfSHo/+YTx
GUW2MkvbXFp7fDWqKTf0Qm/l9Kc73Qklg0P6z0aNtRQWhil/i8Ylcj9Wzmtk
8PRlmpunOhTgqgg1WlOe2cx2pKYUsk+6LiQ8qc+ojvmK+FRAQWfaJfRpBVfZ
nzkF7n+Tiw/6DhOTHPn25oetyB19yXP2WkySsXukZC50Re2HcCJnAWbFW/06
q/bsERRzqYNROkLKQm6kK/Wsk77Un1OpbO86GifC5sLzBtQajOsCU23dbk6A
y7S4ll0SfDGji8Ax0xUh7gEcQm79JMwiTMuhxowjLtth2bSiqiWz2B23RxKg
9yKUnJTEY6UrcK7TPjq+7JW+7Jmn7/Xj3K0O3wMn5fw8+fCa0cVwx+sy2V6+
Ujq+B4C3r2WEMwFNjj9FyYZCMaTwQMc17ggIgp958+5rzZslHQAfbiYDY0kV
UtxBbar2O5LD52ynI2nsAbiQSP6V5a8x5sJxIH08EJfKRxcUhCRi4Vy9NkKO
XKYaC/zqDQweKaPnZ2Mn0J2RZEN2RA++0LEFxHqrLlFeZ1ITvgritJ4AAACd
oMDaC+Ty4Y3XdhWHpOkwi1xgbkiNHwSoNipLXihOyyFs62FtwiL6vWg6fEgB
uT/YjfnnI2MyFBO7qYjBwqlmpw2gue3xM9ET7TvnSAhwqv2TSIpZJEgvByg1
ncIRsQ71HOisXNFBxExK58bxwhkPsEs/oMq5YXcTPHJu1kKClDgOP1rkIbq/
Wf0T81zOfQqH38i9odD3qVcW6gLkabHsLrmt5eSP9Rk1aGDX+3dPgdyJBQC0
xsdWGcdhdKoNCZZNKhNOEkGbxEOcl1kBuMu3vLwpz3FjFObQWY/FQv2+pz4z
RMrjbmtjghydDJjxo6EOEE6LvvxmEvK/vnXJwoR4f8uvyP1As1sOR7mht1fC
zMDRL7abzlUp1tkLMq/hV0XDAyTi3BRIKfA+c0hWaOCOP0E9HCnV+PVzxXYv
BaRuOpDEo2X7A3u/2AIUyBUa9Cf7O9Ski43FdvrI8IlATJpdebwCoWOeG6pp
Eo4WsLwqd4+RIAIWqsXoJLQo2yQ0n2/5L1GzcsfiaMhy/bB+OKdEUGWjzVGN
KiB0RRI2siv2j4EwfNAglcfOmnrSkSxdB5+8AcmXNpUF0sM8tyh4jPH/M1mE
iOep7Esv0SBd8aQ5EpZWXUJM4FVdafHz+CwQk98mIyEPkHuMCx9h/7au/IGk
JZcXcQgHptXYjCArA0hw6jZYEn3hlMRrSExKK3zfZ0qZ99qOckBC1o/CCqUO
9Qzu1uOKi2xfnxHF7ya4rAKOIKvSYlzgUqse1Q9kJWao6W1xDpA3aae7XfMr
j0bfdbd7LcJYbnujqhT6mdTLoYxBGq9n0W363uo01imNaVSPHu07nsWdrw8/
cOw9xkstppHjV4qqpZNCrFgzUp7UjLWWcNWv64zLVad8BafRVV48TYz1JYMl
K6XNUSDwrcSL9whMHMLGxFsc6udNe/EFmknwla64jRa2BExIdbVeOizfx59q
kS2jPIOBEHWCpXTg385GMb2q4RZ7GMz3ou0Ri+NZKO5Z3TuzfccEyCC1Vn+o
Z1PYbvI09xPzXodoYLwXXiqOp75Kfo/Zm5yM1q/DhkCcipD+NQPHlWBAfmK2
UlNfKJnkjH2UmISv4EIUi8+o+bT1G30l1U2TsTxUkGkEC8eZ07SSP0hPgKIM
kxOlAZZz1azZigQKPylMeiInp+Pu8b6w5bWMwfennTpnRXd7TN4+3X/Pop7q
Nabtv4x2EgLQtxvHgqDzMPELTRhHbUBpyWo2RZevJo5XTVL8iP5QPERES4QY
UoQBMtU8c6CAN3NUw4gWSbpLq/0YfPWCViE0oUt4FcYCbMuqe9JyF0J5XTZt
1XyRN8MBbkOwtPvusKaFs1nzbOmXNsMKSgMW4Na2fv58gs0/SIZnXEaoqZX/
j+NEwZJWpCRUKMdm0lC2Ev873VOH/2OcqVG/rCO7spY6ln821IWpqhA0b2wU
wt8hybKCu8nZjNnHhMUPomqu62Hi+nL5xqJr5DN0lgwjfC4bWJUX7A8Z1ZR7
+I9NHFj19nuLlo7GEmEakpKNkSAHAy7NNYP2FcriDmfhhnGBWytyVS6wtVvy
2ro7IdI9qgmxreOwXg0e9TaYhEHM1nZ6256HOvH/CYP3XcKt/fBBlXiNR/YU
lyOJ2iAO0vUOyyyG1HBblEnUEtL1duF3e5X8LqwHdUBARzfjCaVmsZdYQPaq
3CO4KaEzzqZm+e5fHDgAxpWKNHjJl7G5LTJSi7VZeMc+09rC4qCBEiZy5EvQ
JRtGnXjO37MfMWbMYnw90F8bwynQwQHFM/eUB+EM74dH8nUCtAtiIGw93zCz
PMOsMs0QBqqE9UCgxzPLic+viprjFZ/7AVjPse3vfzFpcUMzKM/Oea6H3PBp
cR+HNsIJEbfNoyLgtjx4wfYDkUtI+m4J6upv5wDfbN/55y7SD3yzoBl7m+bc
4x2EILt/HWjsYZB2Iv1z8pxOYVd7CmP9Q6SiQtNXA4FSvSU6Q5APOW7zH+k3
n5Nk35aOiYih4sQ3t2MwYkYjeGzpGDg8yA5B5A5aIWIU66jJ1Iqk26C7wdUh
55afSQkWsW1s4rnNkE3EhoQbaA3b2xk2cQnBAszKSsSKyaFJN0rJlSWzPJax
7i1EugbEYknd9KWjJoZoGsDLLLGhWAj/cfH6hd0E7pNFuR1hQyvQNNpSIoXv
tLJ3irVOZZVQ/1rljfYSPSWuOmC0Xu8l/0aTnYS1t043rlc7y+vCt3JtT7sH
vORM5j59GyRkfz90l9FGVp1opxqfarDGVNhyrhN6UYZdrwELMEY5d9c03FED
rw5JOHsBsyEWuM5pqr8nAYVPglzEmpM351jkSl++jLidvNOAUpfKF1tZqnFL
J9sWorVkVbHKnfP9nXnY0VK6LQjc/bSHeQ0KC4a7QjxuEe8VLbRE2aruz89N
vDOpFJcTWaDBIiEpS1BiLK7JIhGIcxsgE+UDErOyBgdOZbVsl3y1gxTuulC7
bxsEiouPdFaQ+eG9ksA0Ke7GOsGDwFJtvc7P8bcVBGGtB68DH06FJkEFthpL
AOI9WocKEbKG/PO77ZcqSPXgmD15nvvjKWH8mHCpQMrOJTeQj5BMs+OAnJxK
vS+NfWARgc3rrhk2nKIjzX9+keWLd/jwKTD2gFO+2+MtklUS6ASPtHWoSqA9
zn3lzXNzDK6tSSGdM/pAwpB1otQhk8ZpurOp2v0dRKJdZ7JvUXTSQ8uTzSvW
i2eSk3HaxZiQwO8B3zH8M7X22j18mEaKDSCd5WoNT7J/5phNFjeaFXKVb1uI
PeT+KNXJgYYvbv3pkiLTur66rGqld/S4/TvGr0IJMcwrmf24j0J+H7IfsaC8
+gfU4ZW9K6ZVgnB2KjuTNYeMzuM73V69kEzwUs7G8ZaFmx3SP+zQ/sO7xscW
sT9zTQSMrLbLVepmbeMFNrCQldbO5PNIklMmZ0PXJv5MVTUgyZ4KhIpUDnKz
GwKq5tuM/sk+EkWmnFIlqs5dOqtmCJBXHvwNmRAeINa5n7ZnwTRhHKrlOzkO
gIubeYf+FJu6MaClR4l/U61G+/U36wsO4Gu9O1SXeK4s9sv7JBlcA2JrClYP
zRRdVfTVcXF3JJnfMQXLiFYdJ3+vJhcqyFlb49KWHQKqo5k+AoOTyR1ixzCC
Odl3LCHLrWRvJQmUTykMorW9eMKjnLRJkTbUWNwRtb0J/Nn5wzR/e2fgeWwG
q9brcs611hk8ns6MGeMUqdSOvzaJu6KCqxrJXocArOVhN1z50FGc/G4lWB1X
ChijZdqGG5TlLlgSEoQ+LgGWY3+RNub7xPkATpkrOoow6v277/LLwlYp5ka6
Ek9UcMJCDXjdR6RQILwvUtkzLiPQF0AlsH5vuyhPf/yDukg4ot5HhhrG6Ezo
zK0HYQuiViMGee6xIUuXEMNA1/nLRmXID+KZkKLJ2B5cdgiYs3UeGtbg0DWJ
qjAoj09kNPnD9KuqLREHiVK/u+vKBHd4QrgbSP/WNyiLcXC5oeTkYgqmWE5Q
E3R/bz7WERZDVkRsCnRRq954hUi2SIk/AsNC+ssUxasXU+Ks61rwP82zLCR8
URx2RSYvw9+yqtj2pZSVBkQl+4S8S9IXCWCnQbd2QC0mLzpROK+siz1Jzb7U
tvMQ/nGkpe+WgsWmiFjao0D5axqkdXJkWmR719H/JfUUvEbG8w902YRynxDB
V7K923MfEYjymfUQRPTxlZgGD3fk6027WWk350NaS8E9Kom4GHdlsfcOdHV0
Gm1jh/7FXO9khrM3OJ9uvIxCB3BbZnrF/KHvty6ngWHnB+xn3CVxlGDUd/EF
UWkBQuBohxFaRkwZLGf2gR4/Buu3NQV/RnUQ0KCN1Lx0YbB4N+cVyOLaR5Z0
3HUnesOvChnkRVAtC1dtI2MBnVx/8T2sf/XaN8EFEmvQmLJhgFaIuFb58biy
JSduYfPocRRj1bbc20/A1XnCCG6jjfHqJYjdoxqSJE/XTG0Mt6kTxZfhxBAr
PL6C4c7O6WB42upc805PyGiwp48UvlYfPghErP/CcSz0Y7kUevXy+BeE+l7T
V64yEZWwrwa7erOoQmKjNAG+ziE8YjrTpaUXHeiqX2s2v8MvT1f8Gr1jfySj
Ncpt6gI5x7zYW2LjI0gNYypXbBr9/qKfVlr49Il+rHOybbcI8mZ5x5ES+waz
ZQBqN6NDr5xSaMe8cFi2Mf5AgLq0joFgDd/DcVVP/z4Qcqq967EUIYAFA91E
EO1JFZ+r1tmTHAGTUGljPZ7zejHvzlnLCJIUMQp/ESpD5fzw8Wg5/4YHVf/h
UNhQgkvb9j6t55TpwDI0Fz8iikUyPqe8VWaXj0Kf5K/5/6woDHYHui6UhO7g
aDOUi8JLgJgLAI6l+eNWPM3pRU3DmlDjnZA1oF7K7M+B7EChBWGe1vjbrLX8
fmS+D2cYODPK5tb5tSEencBEEGZPW27KKAislvrNXKiWHl3KACnznU7LSPC6
ikuCv7l7YFVUP6AjcHmPN/25Bc8gM6YP0Gygjaah9T/h/nCFzKuZD0d3l949
5xeONnUE6cgx795xsGQiwkdnxEaxR8ozZhIEwaXZets9zvVObvKaPoi/N2hK
jvQ0MjZlyTpD/7VAxUOO7/JA8+uR2u0LP2FPDap8SS3pe7WOVVzICFIX3R9s
Bf94d8kSV7hJN+JXlHAaguljfIh/svC4uPrJNXNbw9pk67YZKDYWBDcRfC2q
AsHfuBjMhZuH4rXd+G1QHq4or4yfaURlewWz5XKW6Zxy6dLP1r0DfRv0v11x
B1Jhqv6EYncMt0+sgf7KOb9rsmzjgLVwvGTQB3YZf/khcLkOXhp3fVkWCQTl
ngjp4FkZq3oSxaRIIuto4ik/eIrNQcgcqzzniWD4rGTVwEygmmhuRcYyw61s
H3zNL4hmnu8XwOSSZ9dZEoUqfSJiPTJXwUeaDYVA27P7UYWdwwgAuXKYgt87
WRNVIjWUNg5OXhBZDwU5flmdZ2/L+iplmrumpi7hvjaChSoHYjPBvzUC7cJ5
Xbp0FLPHBdFJVlig3HoOGskYIDldidNZ4n2Ncqd1mZpIZNy0tUVW3PHLNw2y
h7zyi6RjNFcqWrDzZ4mipV5JJ4l9z1uJoqn+qHbwbjFfHWjZdHzh98hKxzlg
MLW38gyt64+3V8yFrZY/2a8410cm80mK9ThwB6msQWLfSy3fyIuDt57OSnsl
GER35R+Tvpx8Lpwa9Rgi+N/zff5zwh2q8Ly9TIYlvasMM83oaNRev0AyoU3e
oQDEwCdTOp/9Vy6EQDqScASRPv2hwTIduS+rHL4W5bA+uWwcv/rrnprhYHqm
4cjEouWOpFJ6lxszGrS1KsOoLwMEx2qVw0uA7Si9GuIOAFE86wXmJOZFNvEM
3JP8hNfJD07dSwLPMz8rY0YrCufegWX5fmI01xhrAuzOdYbY8PmQxhvh/R2z
sh2AOy1wU4UgUo48bZ7e7g4CFXKCEuVsZsWjFU23jGY1beYxr/oibU+PGPx1
PTDFEweZiYi/gC2cmOocnrd3kaDRVlFpWV5TfDYeisvbZT+uTuDrpWtG8Y4z
+UFOwzVU4otQ/jWFwQIbxingNcZdz2FZq3cAEuhxOuUvExn7z45tkLpiIUxI
di1J2QoWFzlMVOX6bTqHGSoDt3dDCbds4Wlm0i5QkTcDUljwW+fuuQgo9t4g
6pUTKWfymCPYwLeW+IFvTYgUuJwE99dluCtVNZhIKD/RLxLOBkVy3jtdelZs
bttBAeCi8AYMvSiYfOZ3McN09xbx9FUIrin9Zcf97C1QuWqn07JSszxJiQBt
9sxNNGBzzaAgzix+YMjCUR3OQChhf6ZjAT0Gb8pgsugOMNn8G3xDCfwUcjCk
JMlCp4vPBSErTVwV/jmxk+CnIa9yWcVqOVaTqpLtiLGSw/9wUB6NNftUkXu2
5UicgyHP967+beJ48Y4GcRsXYE3r1mR6MYO/xCfkMlkkCRwj8ZTHiQymDKWn
cVtezt1l9KRPJfiDixWfs+mpLz2gtSzAaejcSIPzUAaT8P2Eb+euhI9yktpp
ZhP+qFF9PtOdI/Mdk6X1Ja1pxLjRMXi5nMfM1Uy33faldMbdj+6b4E7/yXct
64gKPFnZ5krV9RuWLBYYZrJZ7xw5lkNbQY6YXUqCXJ9SGrBsPWN2ctwSpDdm
Koo7C1HNKmMq+e/aRfetu3zaIVMOPMxx+L8cRxudhwll0LBOh/pSuCj4TyhC
EKrp6WiqtCit5TrHRagutg0RxoVBUOcjhhs70vjJ/zWiNGVfmGYsHxKknT0Y
8krEmNVXRivQH1uXbYllDRUApJ6G+hkKDFZihxU4d25wBXRo3uDGW3Xev6nm
7gC83kCpcj/LeNc6GiMBSLPK4LmFWR6LzDjjvYsCEnDj7KXWwLaf67TtwwCc
PnNNAzye+Y+TG/LDQGAxlsqJ1/Utvy69LqVYNJhyt/9ma+pXSJXxYGgw4UKl
vt/AFVykQNiH3CQEmfflajPvdtVvXRl/s+a3Mw0b9hdaqRXaB7Ipb2qlkWdV
+p2InqbrRq/CFgPzWC2JlsfESgSlZTVvy+7EHFIjNvO8NTLj7tAWrd6HZLYL
V3AZxoVjNopZxtUG6Q2+HdAd4XmzunE+FM9snRS4S8e/9khz0T+AOEF9eR2+
RYK8SmIEe8yZIzgTalXoFQCGl1QWlrTzVoj0vWV4FRAdqBOU3ofIFblGeMT6
6FtNVhe1agPiNrDe8F/XetlY5hXBSwlboYx4s97WFx16rjSZ7GZUZ4aRxXxG
4jMH1+uYJoLT0WgYrWIysETsg2r1yYaFhwqOZS7mv6jyjj35dfssPJJW4Pvz
oPFH8jeI89bew5WMzwJMcvmu4l8BAHUOEcwuZoMzBiuvEJt2vm+sDTFRSgdN
SZ10C1HwZIi9BmlAT8Px5cpQWsmzqDc5C1b3W+PniwBtuc1BqNF2WdwEWgDb
0NXw0+TF1lwxPlZQvj3zacdQy79QLdC51Z8mMmNhw5XO1oH0/lhyI1loQWE6
5wS+Z2YuJ79g9cptpd//Nl83cIaC7leg6iyqOxHJBLNRZmp1RvxA4rV/Kj8e
SGk2bUrH7vb37nKwhhWdVeVAZpLrnsrZcxptzcOSuwKjdBhsR9DT8V6v1qHg
hxG+EQy69rvOlA/E4MRCbLvS03A0Wx5FW0fBFA/O7HTM7+ROZwY1T8iP+pNs
bHtP2InO+F276V5lTo9wPglPdNqLlyslPgeM/DAQGg/yFOnBMbjlnBSmfQQz
kULlxCWkbH1FVXVEGaBug1g/2HFgY6pbf2Gd1aOC9aysjvNrETDPkv+DkZ2w
Pnn655lcks+telgyL8pa5FJ72eKUsZ4a+MNpRt0KBGCGFz7OXezPHtNN86ez
FF4eb4xWWCbY2opWPfx0Pa0AP31i8RhnqEKM/6pWWSxNoL5IjBCMAifD/K39
7aI+MUHIy0hVuYhZ6YTv8G1BtTEymfGtlzmF+QDIgx6g2Jn5N9ryLce8cC8F
Bdu92eYxj+59imf2fGnd9ktsfJEA4bIBbGGYwXWir87PhbD/CGCMfluf8ksi
7yn/K3TQZBkzXwzZOZu5B30j6YDXnrJPNcCndd+tcKep4FqJ1WHW9TlefJlC
mLN5Ve39LkbztSiK0dBHcBRzqCYEcy6ZOt65/K6AmRwl2daPpTNnA4dUGZD2
eehph9Jtl0uxH/m/+zUuhqpcFnjFimmv6nzOowhyPMfJvh9hoUmMDqkF9sVn
nS+xJPmJMlsHrBMOsGgk936RZjLWsvd8tBq0URGUESrnWupyIinbAmOFOM4j
5x+CXqOYVspVgJ5q5MchO0EznpBd8uEzHxFtkzmjQ4PUUeoBu0KwtEyTn+Ss
eEGGnKWJUbeoyq5Vn/TeTQjMW/M2/uBJJF9oZ81L8n/8F4ptqVPb2ZOtNgCY
fGVKbjMoBYWi/8fqsaYjQqu2UZhU/Br0vDsWBALNcMbbFlON9Ec7a5xJjGJv
MMnw0LsdWz5lT9nVFqSzwIVOj2d8wN8OEMpD7G2dGq/3AaMSYgxipZkkltjl
gCmm8rskeMaHRQzUfwPtW49/FIPuVBbXydFxhYuq5h1UBF8hBIt2RAaynQRp
1wm0vhXhqVNjJBslnm+CxhWwVC0ZHOeRqBbcyz2wCjf9Ge92AGZmDtx2C/wA
514GwcrN3YrCo3U1gnXlXXo2UQfWaRiP7N7MdXWhS32Lha+0x81xJAtwxux5
7BbQ44jbuSKrCDBVyWJJOzX9DlGF8eDprqWAYBdfszoyYAIOjWyM1J/2g4o2
zJKXdq50uEMkppxCMxzQmPS8Zqfod4tElkbmolIyxssrTRyR/SXGJoSbPS7S
xA6QJtH19hXPcQp35AavGp0o12xj7FsMyF7ZDYc6/2qDUsfF+fDfs9m4lveq
Aasy7wVZWQ5t8QOGFJhgYbk8JUh809rS3rEjl4dG6iPO+doxSIuLd7/bbMEU
O6h1wxYUS1fli2/isHGjdsWOFvtQv5CIDQBCLKFm1yMfNAowYuoHdVLA6+P5
aGrv78M5+XXmqaaCQ+oXOq/w6xFeZt6OtR3PiC8EYd6dNNUTBkrwzNu5cI6t
0bik4YgqqQ1OD45wfFtc+oIcb4WRJcNdZ8hkvaKAR1I3RRJZi+2LK2N4Dn8I
8FiZNGzIdPWz7+IFyq+F87S31oJ9/5v44HQ/3Iwz3hIxGM3bKgLL1nJUP81v
ksl/Bf4FTgADM82wgjaNHnB4nByfs89h5jlJ3ZlUqHazBjeG9Re2X5nVzQA2
bXo2ThRhfTGByld8WK+gpE5qAlZhzGL24y6Oth9HfcK9Xm1VwLL8P7g7GXBC
zAACdp12hqKhMLL5tb38jtQY1BGLrn80cLaNX5nwzswo+TVuqTHLkEx5qBnh
u82Erm8J+bU7ZKRWOdVS4/EcLaC3lQE3AtBsN05LAX7/A+v5sbs7yV7ncFoz
MAKnQmAYb/HV4BAyRjSDpDa1EEVnVJ9N+Quvvo8Kt/DDtE37fcKOsVRSMwN+
7ULLwwkIFRdZtgz14IqV+guNFQiQOIviMG+SsodIwcSeNNEgobXz1A2YgHJY
IdMaIDNTD/IHHoZImyKS1ACEMwBN/aspQyxXMNSQx6RKhK+l3GpBkhkKVXj9
YMOgGpjSspzHQydAnU9FLDa78K/f9zjvdtL4mcdqhinqRNXyUl5d1LHqa6eN
EtwcyJAg6Dw3ZeWraNZXBbWBgbi6+DQgCHJjKGKRKnKzH0uapZeC5Y26kmSz
aaHYYChJPTK1rRoCYE9ucNp5qtpmIyYi7Wb5zVBMmnBOlVoC1Lx2KVEh4tuN
t8N8VL2B8L20xI/Wbo4bGM1CEAoUWKBdMbmkB/Y0vZy+1I+YXgvYpAOB6TsG
7j34RGan5pg9qxi0VfpO8cB35EG4EG0CJJogkf3xO3b02++Az64OdmCs2cy0
e/TmTtcdNqT+UvaJydZtCup/yAcw88TDaBG4H0AnwM+KSc9d8jvMo2f85jfX
eIXtzG853xaPohZH9/eg5l/4jnDzH8hyC7LtQEycVvOt4zTwLBxDsQPzCPy0
iafLx/GYs/EbK6mbRuRCW4DMFA+MPnsS/exBFKISITxFPje8cuTSzcnQdIDb
FILt2rFzmLXEaSFH9TvtfA6SfqVU7b1ZgTRjGujQBnD30YMhhXwFV1VkJ03y
RnKkTm39w6XcZm1QZZYWwTzHn/oWupwwQixHe6XoUueAsHkvXVbCyihSzulj
7fIzPUqCurHecB5EPYsvIQ/6+n0AKfCaEFdPNE3ntLEFuv6+IzAKu/J7xNhD
Ma4+g2Ij+VPxs12AxtwGsAGG8it0/62u4KyTJRx/OZzIEiguNc8sDKeWcQ7z
9XNlvMwg+IbUiyK9ePZb2Un37SiDsdXHCIGd6xsf7LSfHE3TvBL2YdkVIB9n
3ZraVD/Ldb0+meIl9UGsuJgKGy1Etp03k4UQaO/o4YmBNa9rBmsYZjakDYEz
ylc3NFtAcm1WHDDyG/HPltBzpSP2QU90uaXMMJ+EAD8iZolIXYZZyyfvrOX/
t6PfNlFNANd9L3Yu3oTij6T5SyEPtEUaTiEXL6irLZD6owYqFucmTU1rBt5g
yQnp+VfK3sU8J1fXsuG4mHHREGMOgXS/UeGfqX3VP5Q/a/efg5TAdlUAXLd5
RxEnyS9RBTa5TpT0nq7/6O5w/3W4EBqQPniBmDRKUXVNzJ+cRFS0ohVoVlXe
7t3dpSc42aydNEknX2abSm3yQOS3izKDV6ivI+gRY9v4lbGPks8yP/rXqiD9
ZOyv/+uJAmdVO1uD7p9yvJk61l6SArApoBZJUqqMrZaWhe1Ub2QYamdeZNcr
DfC+Y25Ol5mlRp5XoK9H14Aaim8KEXconPnvrIQ1JPYoP5RJMtTLIICTlw76
umQxVuITvzb4yUwSLlpKJzhfFGejly1YyiTy1CXRuj9Chb8TJcPuvh3fblpw
/yaBktdlQ+J6fgLdMsIGQQAQ5K10+RGMeLZ1Ec+qCFgG/A0NLqinpVI1NFHw
604gw4dni6GV5mEDQHz8oWEezQrxDta+VCv1gvt4JjkYFbQiqiD4b2yOURcH
E81CqG4doijd2ybSHx0jhSiVc9UJx5eQzNxKDL0Mrze+cswJ4KJs5EGu/uK9
9Fh5GxI6Vo1I6jAJ3/x4XNM8FHIBDiyH3mHRbL//18npS3fdrvpFiukrIE6y
FP7NM8E4IeNwubT4C42wYQgUeTDaSQVrg/1+z0FupD2Kz/f5gXq+vLte9uze
8xfgbcph+fw9K+gXBbhMi6RypaDLFNceCP/UiSmw22BnDUNb+5CYpxe4eQIh
IKhbX9xTRtNTPYyR5RW2zPKPJRXHctJKGath+o4gz0UvR0LpU1azB2pMnMi/
pccCy9oC0Q6+LX3COTNnTQAahn2OXkjzoFfbsEEnl7Ugv5ux4mI5fwYgkKtQ
Kg4I6Uf5p4Kpkm2DjXuKdPmNc2ljARaGL9/X2bzgsvgoQTOPwpzbLXwt9KK0
OFcba6pjV4fViIElmKR7iDHYBr28/xhN6Vz8y2XQmBcOo3PLorJaZ4Mbbk3/
NUif8LJ6J2LohSDbqVJvv3Er6QQXdBafFczo3wI87MKW95KZWZAcDc5PtW5s
10xDAJxEiE1nvoZAzLuz+bX8eAJOjG8SAqprMPuivCNSc9bBFuueHrJYQhhk
8v+jYK56LCxclkMXj5QMix6CIbnbEw1imP9bZUDnD3EJYJfgMaP5NBreKDi1
hAJGZfZzeYcgkAeUvsExb/t4bUqo1gEnu8/DzjdCBfEivNhvtkiyeHS6xe6y
J39+64PBSQySXTrZjLvkLmx4Ih/94UpJy5gXBsLZNHW0TyBnJiY0akF7T8+q
ypKavPlmBMS+AxT68kkhYl0pbweOeVmT+BqVfL0521LBwXSqmdK6DHMXhv+Y
2FPkiXg62LyaqXV9NPAQrsLiumRaHBKQXt6pbWtpfCrs/0LPb/7EUZF0CnVF
m3VoqVGBhU5FOxqwEUjWZKv//2t/ortcKJ+RRqi7fkQUuT4THUxwsYuhl0pA
WJFQNp9osFuSl6auzKXy8BoZTlwG/N62a3DeNTRaSW7ziMt7qr1zCaipeajp
GQT/JDTI2gl9m8g4SQ2c2QA19Ojw2Wrn3fV4iWjGiF0H2r7rVJErMZOiK+QJ
9fT2cY39bgRp3ZVzkbH/ogks+4F+wuaROeyPX187PolcqxFK4zot59fu9YTr
gypUl+ojFPMlVIQTL86FaWKuX3c7+U0A/Sk53ATqnZQPZmzt4vuQB8fpJm47
RbqYnRcUmHiu8gpZ0s3oecW0V6fP3OLSmDEeZuFXLYqzi2BL/nb2Feyha3yn
a6446154mmt7qiph5/9k7b00KnLdDHm0mtxdVBXRmvkSbD2UFZkkAklV479u
xuAPnfWvPdKI5sxTQ8tam5SamzujVOaLYUK9hTrYw4JqNvQTPz5r14wXUrG4
4lm28H8+RoSmPY1n1V0P2iQ+5hdFSYmNtkRiLOrO7eE40Ty9SBVhWJ5/42bA
sATpMdgU5ThREbcYtsK9udhHEwsIklnOAD1Pe6+aNe5MFghSa53y4ZQeTpMg
40OEqY19CPFuLYnavYoyNdi1NTHWrdNQqSFRhaVdrTcMqQUCtpIxOz/ZYslm
4frYf3F1kA3+zWXu1WKYQv0Qb1DpmnqHSTOeWgjCT/kIKbnr1uCr9zu0XQbC
tt+tMPbCqFhHIiUgID9SxQToioer4iGGoJBqYZG+mL4MgAT19qkuFDP5sKQy
pJBMyOr0KhiJZZMNvM6tfzdD/lIZcA7tH7MP3ipVVSQj79WMKAhbQK7bN038
XcqBRUWk4VKS0dG1n2RwVltlfOgTqq4VChzlUPiEvhb8APt78eNTn0e968TV
VRzQea0aO9CMRG/kVLZnxDzkwIyJl+J8j2tHKmd/Age0PmUf6mHNE4AnLGfM
T2JbW3uqpkS7sFu3ekVD3aXnUCHyJsh4xPVNM9GwNmW4DntwLoc0Qd4FeVyD
XdNZVEDiBg+n3pnulhP/voHceaHnkBohgsp3o4ihLCH/orVgnz1gEzsBe0kN
FaKBArHhSHT1UaZ3jSYkJ6SrAhoORtuykpa10UZzgLee1xjSeTEDfH2HGH6h
DU2RCIZTsEZVenRjy0JeUmraJ0SQNaQlwRGvEUC40LCPcp16OMmlirySVxix
CPPOQOv8xY23hKbnLJ/0BBNv7acpSEcaakvQOFy/1TBOtRAPr/IVuRaWKqDR
csbRq4RGuj7fW3fPoQNQTwH4neu0KUa5BWw4j2yLZ/izjKBPmSmRV53UFmVt
ncHjNOSxcNbGTDMcICI7PGiVVlMCTBu4bbJ+ckiGhnQjWdgcNK6ReZ2BUTYn
zgmVBPPeCZcgc4BFN0/aAD7TkPsPHmKE6J4NIe5XkoApl4gG0gbYJKetB6VJ
MM28qCrXTHTsXSlH1WKbyhTtInaG1oI9fYHm0SMUFRc6POxcs1+mkrNx9y7p
+3rtpRjLuEncXDAp0EjJurcWJhknvjKCtKavKZTBX5TH+7Q0gqL2W2s9VbHX
XKr7YSAuZ5v2xgINGKptXrZoh1M9+0B2poIqUH+u+VBRJUfmCTyMeE3gS7wx
Cyeh0Q4hPyl2Z8q2Y8FD27ydrupbl+EkPQzbBefQhmP/2sIZ2GW3yVnyD17C
TEHOfytru6eGpSQR3xXPgbLAHIczbY3oBpA95UZ8VFtG0fGFq/9iV6sM4HkO
UG4P4iba9IS3DsVXNzx3Ju8NZsCG/ohWWwbpEaFny2A+Sd3J9O9b0tzAwji2
JevpulmpU4s9gyyQINlBmx3MOX+Xb4ZJqYgZT+PuiezJmX9tH2KN5ut1fLTd
R6Hd8WRRaSpjb/3tq+JGPYHzMehPZQWQy5dod87E5LiFOA0m32xblo4iepp9
ueMbWUCVmYF/GxcsHKmPJW7eVuk8aEEZKGY1QyrKTPI39MCUgrDlxJVTv/Zj
MQjAmt965eg4F+uGyjHBk+LuCcACrkTynkJE9wFZLdAxFbfihWE0+L2h1+6T
ii1gpZGeimoezfQ3mFyChzZ2F+N4HbZALQ/V43tfK58MQKfKlL9IAVJ0cwlf
WK0C7RJXjF13/oAXwdE/itl6/Au4kpZEZKmdB0XBggqMb810ASe3KqKA8wRI
xcBRqzcyRx8EPGN8QVC9Zy2k9xwKsQJCBiCdsmP1Nw3N7uO7t3khiEiU4na0
KKqdtV7uZ0MG/C8YJK7v8m0F/PIXYaSHHQwzFVGvrudYEaLXRH6/OJpPcYXY
YsX7XtmB1WFBRFuYXPlnIA5K06om431ecx0oalc3vVwSnEBbLFC54sbgmas/
2D1pdj4ZTWl+fyJ8VtMdsiLwDhZieLe8OMb/I5XOuvxa0NP5dHwThScHRFzv
wU3jJcX78H+a9JEMZpq6KVnmIlNnd8H61DEBfNMUptalabZcHObojI1N5EnT
bAPpVFY8NXy+5hmigIfaB2CbxHGe30m7fpQlDtgWgbRFZ6xLbycc4xRi9NXE
FzIRB2swk8ryn5dpJgznCOifwZRsxTQR+ZUZcm+V/36oLkPP/lAownYC1cDK
MrCTPd+KtDTCRHQRhu+3SwBccCsOnHwG8DZpQmTzsSTnUhuHvdmjokYQebt1
XmVZdJ9J9p1+12Xw8IPSczuQldw1eM6t9lnJ46hh5YAUfSdXQgIeVIsgHrBw
jUfESkoG+ee+Ve37oYBXnmPvst8b2yJXVGD22kYixxuTBpcTyZQ5NuleowAH
gJozNVCvyMyGjd2NOQh3E0z8bWRGFuQuz8iAZzxrm0i548jbQt0lNvbsIaGX
R6S7mdgoTm26BfsdzwjQn5cJpEHC5YDAaulY+1MUTLCrecJti+gywab0CtWX
NWBOoTjauTrheaycXAvJ+Hwjif04tLkuz3D3Uq/E4RpVFBugRNjuXX8aAGbk
Yr8nPEpv7ORfwxOXS5fvcwFYsyEitWBLvDH0UHhDIZir96MDBMQxTmF95epE
lM4mRVwxLl1+sfJD6beSe1zu7Sq89LnXijZZQ+DQHAZEzxF5PYzBxnDuT5Uo
CFg/VAf1xK2qBYeXhhrVsVH0AirZwHLRtag40r3JvWs67grSf9fA6W9q+X0M
HMz3GVZaDjNgOvnFFLkdRyF0C3IpYH+Bp4CacdOtxzVqJ/75t/Pde4eXt3S8
MTLXINTtxNvNSE2gDsmsLOVjFFC/3cUdyE6q2x0fYQD68a6OAYHGs1sC2brt
8ncEbLrxJp3tzpcgqcB/Nj2ubuOGhUVkwdpdd1jfzfywL3Yojayi3SygfHb5
TlN2gZ4JrasmqFbI10YO0KwYUBu9xXVYK+HuKUJ3HiXSma09t9QxVfkUu53w
So/4MwM0WmEw6oqtax7eWar+UW07fUmfcTy3pba2hoN7l+RbM5GGEiHZl+WC
GFpkN2ob3VWvCgxiyJIYOnenHmWciFfZgDHmdZljR5OXQxZQjr3XFxfLhzeI
o7KHW3pFh6+XPKN68GlH6t5TLBO2+K7WyKvQcPQqtBW0EmYuvp88EB7lwqnY
AxD15OUDoNQmiv7ryhx1eLXS1ZEdBnWHBiZt11IFirxzK9D64j+UVBRfQdev
uWSvL+GXNkOdgFhYuUDkZF4B/eDaQNs5oPhoCcP9QsOPk2nruBo3dDk9t7KX
3Zowt7mEZVCaoMx3tdljn4XdC4l+Ksjm2W2S+eerPHv2Ln4IyzrUMQL93RK+
P65kEI9AQmSmtkhQkYxtASYl9CwU/9xTR9WpasXZ7ESIkGGJ/Xcd41jFePdd
6UsTkk8g9YcWd6yOnsFHxKDZyBX8OV1rfvqqXCrlQlfsVTYzJSNN6fNE5K+P
DYx+rcw8aOtNeGwvi74EW/rFYIrd8p5GAiMP58ih8nfIQSk2yUzg5g7ZFLMq
gjaJIOCFiYBC/2YxPGR37tsR3/7Bht0lEVy8VwdnckgUz12G3YdagJ3EiRpM
yTr+k1rL5/pr5FPlNLh6QhG7LGSV8JhaNcrBbyUyNngl92BHjw7nBv1tmTy/
BTHzaOvCSNcNpyEn6unXf847GA/I4BqRZOq5aQvCMHDTxukXIX6Vi3oKvBU7
c3iWz4qFWd4LuMNOPnuiOQQ1W3IuNgJZ1MuOWow+yjriyRjT87FmXywk8WVV
kqbYeWaF7W5ai6gvOxG+YbXt7tbtsuAINptZ06aMTydghK+E2tN/IGwrjpwL
InpXM3IKZLlhqfRBcCbiGEVj2Au0Bl3QThTMyMucbxSZ8gCd0wRp/mb5woKm
UJSmEOEaTC3RrporHai5cgqy0g0K6uqXLd4dORTCDpDNHSZBOgCAmrqeRIIL
Jse7cP0gYFL2923GVg4tRFr9PYhOk38qVcJZcablg+/DWyT5fdjOo3BwNOpW
pc2SWIKSBW2sMSVMOb9AvmrzoRkPgExl6gmnitRMn7QdjRmHTcItl188q5xg
r86uIWRHRkS7dYwHODi2nHSjDzQVd2Xm64Yzm51H4FKxU+hYfvlqGca/0Umk
y720WoVAn2eka3Y1Rurdw/M7YXAFHYQ9w75T+j/KXsgHB+KVERBjeyJuBvVZ
md+E6yTiUnTfov6pNbelLwQbiscdcGEhSr72YcvynRFsDd94xFhE8jbhgQC6
VxzbCjRyBSZ5JphjR3t+wG/+mZGFL81j18S3vMejaZDvNEjP+5uaQQLbigYo
XVE9BoPy4awTuu5o+CygDmNoWd8tTpmyYFctbqKKkycL7bW79sLJ5FBrCYpx
8/iR8Bs/mF5UAcfDZRAK/hq0EM8OdfVzLtLbSzmrhx27dOEtVlfwiSW1sJWc
4iFFUEjDKX2RB+sa6ZX2ablRx1k2+wV3AmZiTqo0FhItmR3rMlN26ag100pG
uufEHXk6rzKuOc1aCt6vIXzjpuc6NvYMFIHFj7HbT437FXxSxZtCqCBTA70T
wY0nd0F8ZucZ+jpRf2BVt3lyjv22zzg90ArnNxFH1kzlCHuf9ywAmsnnB97n
1ypFu22168REOBd7t3o0nQFdtuGT5K08TU8A7zo5gfI6ko5d5YvUbm6ibQ83
uUqIraZfL3VAfGRqilVxJfPj+cU2s97/4GfY5EKyYe9TUN2oF2HtcM/1e87r
jmbcXemy7XXCkdz3xwhFJ1n2kIV7SdQUW2zc6fP3tFKxTkfBD8NyeEBAMq2z
V2wBzEyY/P3277geIfgzurrmDKDVePnnFJrm6WTT+CiRntT7k/YfPRsW2vP7
UtwxjZxSq2pM9lWhRyR+OFjFj6ZN4b0AgIrJp7KwyMKYo/sznZqX4lDN308p
hzR1uSWhPS9eaVtEzMB8DeaHIwMiLRnjITllQLkRSkX2qGtu21AICwYHhwdy
kInUpRxljKbMCjunfqSA5X0TH8sROw5hhabU11S3J1eIkfOUAY/dlO5LyKff
5An9XOt3i+CzaIVweQ/ETrRAJaIDSlkrQohrbmzFmrCEfdx8DWvXDOo7P0pU
mUwJhkZSjbTK/IqqkjYyvw/pzM9WlKHvho0atQrSrqjoY2p1TzqFsTuV2VaR
7MZk3HDye6pcmslryBnXv9/kmDygnlSQyZa+Pdh6XXmvYf4T+wnD0k182ETm
8VIjvSc3sBc/ocxai3+BXth1SsulJuD+ONejoY6jPZnBBp140Nhd1RID9G/M
pgOYX5wlozp2vGQYZ1Cxn9ZXPdDkhCffG2TSMIGbHB0BHUlkKzrA6zNThgt4
AkTUaxWSDg7h9fAusbgpTHyQkB/+SNlp1IbKTPJic7+1SKwPnzLe02wo85dS
wwMcm7q5TRPIWaTDz+slXZLkuOdaI9AoAQkaj/VO6gcGZVlj6wa+FeeRksF7
jkq1jWNhVooRKTZOaJ1ddxQ11OcQfTLN/LPZG9n7jCYrNFOQhW8BKKxizUYx
bInZgWDvAzhbg1TXblikIhZtriNRCW3ab7eDevtKMmnKI98Kt/S5DzYEM1fh
dJ1xfAioR3GZK64fhrGg0hubcNQ4KQhd9pehCxwvcomuXyyEeKBOi+3nYJj5
gJtL/9GGFxWUD4qhIY3s9Du2fQl6CoPTV24pV9GyiUjVbgjYww1XJ58mtX9J
2NC69a/ITR8qqKqZerenqukJJXkoNkFp++E1EndZc92zHTXmV8Pq4XXhRz5L
11Zs5DFw+QMxrDARlv4ZzO3bTp9MmVm17FNR4yT+0JwqhFSm124p5RkOdgey
B26dUrPDZ7yKXfPD7H45/xnHdFRMw/CK7TqRvaHDZJR3nyW1kiQNQth59ri1
bZBuZoqXGNr/geVQPlLHgpavobubuGOsuBbhSgL9ZMBKGoScGkwMsXH/LhEj
w1KqXWAQC0h+Uj+bvnCjEVauBeCOZjIFr9RchBxlFdGd54BYpvcrIVxH2L3w
gG0HkrtJMH06QoXE/Mr9qgD4qV1mHk0iJxm2RgfM1Y+ljqiq9ZCzM1owKfo6
T30xgjb9cgZytyjTDSlheBLqJa5sbOrmHrJHK+6p4elOXpPRwN52w/22JGul
7dB97RLuWO07vQuuqzeQeVd2w7tAC4hVUTYmci4oeohW5bHhYMnFZyf/af4p
N9TEFr0C1m+1AVTLIeyQUcmaguvNSk7t+IlBv9e/1CrRpyKWxDI3K1K9NbIZ
y5nwHp2Hum355nx87MoGkussQSY7TRKciLXeEv7Vnuc4Q+ZrVogowb5zKO7S
9Y78H3OlZJ8XnZ6pZCMAalIqneR/WvSQlMWEerA/AbXTS9ssZSGllnrBE5Xt
YWLl/jGU2UqvOb/mdsSYZDmUyiDe8TfUCE3ImnR4xNHjINsC0PWwVA6L6nxp
E71WcPGlsDhVcfAvQcCasb9qjXa1VJ2GN6oRXRjeoNTkUwQT6uokZi/jqGPY
LmvpcGualzV3YhRRkuBwrN4HOI8N87sJkyAfzj0YaoHGgMTNzBfs18ialoGT
A4xRah59px1DCO1YqgIuP5UfyLfXDn1yHlehcasASiFiOdsxN5gpDoQrwqo7
pPJgRGp3yZUD16KL2oUQDA6W9JQp8IdUcfPvP+LdCdesqnBD9dd0AbbeXjf3
XrnrkZuZ4uY0gwLFhy3R0W9RU8t1sk2UKEOGUYPEfrY+vLBp3/GumMCAqj5a
x0KKTzcPT1l/iS9+Yq/T8hQM/omhpSbBZNNwu7tBlmT7+6fsh/TfBrKUnMO9
akCSmwFuMv4UgaTWWr3dcGAbtYJTr48xDm+sALXpjhHUjFbz6Qmi+A3klhLx
ID/45jCfXuh4e6kGg19nLhXZl/4Fdxh87WJo41dYfhGKbX0YIFaz5unD0saP
1ni23Fkl/vM5HzuVIeebf5EMPB+/WtZsIWu+backzS8I+zguXUdD4rL4C6MX
oMq3jGW+Z7aNGEBwjysWwNsPy3RFqXKNdZJgQ+9Ya31iLRyDIDUcziyM5fHt
ZYB8iK8ekmNEM1ZHBg1OKic99kYndKXjDfpcLZq8PtboP3dkKciyxdePGzPC
C7ru2TfXQ/CqEILCvtitVe5/9zOAGzF3z39IdTj0yd9Vi7heQoxfbe+chu2S
PT83cLV1KS+3Lrs9KaRhvR20uoJEt7UMDCOMeM47cXGVDQlNgmkHC6VWHbBs
BRwBpc4V8wAOif3QP25i3pIw+deopJKrQm82ZwU32+ovwjzutBaPo3sfCuw/
/6PRSiyqIeDIbvNB6Kowk5n4GgTjQjVIrVM9P5s55tAbubF6VYB8JxqyuhEo
5HLetTY63GFPhj7FP4Kvxi+TAu3hJ6ccIK/sUwxwpI+hYFwi482V1pXrJ8E+
GmOuRVsUk+ogqvj3XzOO9Fs1tk2yvMr1wODGViEuU74i83NFcDzj1fwQSqHx
FJ079V8KOs7BII8jaZ8HqTOoQKCh9qePk+2GQYm0V6uNcKDOFGDW6vERQsxT
GTuIwzDGr8/jU0qLovZLdpFOQLdO3nRVb6f13i1tQ/buu0qahgAK3UXN8UN3
e8cgegGXA3YOmSvVKYsf+jcwj8pj6dTfcdqp8BOIC9TBvmT7vljDJPBy2J3/
6zklr+w8WKtWAl8V6RzDz0bJlsnA30Pq2oQzsT0+NIyfpgtgnm+2Yc26xO21
5jF1h/6Z37yUIvrDKm2sA3r1pgKiRlP3kF3SS+ZJ2mam15kRiiMAI6rihsGP
nyJWUbZoUXzB2RB0QUK7tOhHnBy8Plx0Y5xebzNJptyOYdX2vyq42Qdbktji
9sV7Z8AqRrYuX7Bj58Wgdkw0Wz+mcU4pseCaeCqx+haPG6kFzwZD3149QhHF
cyLbLaOMwWixR9kLa34GkA+tI1/2yL0HbQ3+wdmUw3z+eSXwmbArc035XWx8
+4yxRiAm7gYnrKCTyHyDlkeyDAHosxx3DUD/zntItODvSv1k5ZsQnzQHmFcK
fhYIJRH/nyCcbyKfABz6aPlmrOHEpozdxbkg9JlPcMPNKxh5jXADRbfZZRFB
2BQBGUuE89bSx2hYBqO+AyKGRXjqN27ARP6YUSM2ygrvcPA6LLizow7hDxE9
9SYQmYwoE7ZamF7Mz/rMPOVs1lRbqjXome0kdtwwlzzdrzxGdDGIkje4umol
4mX2WzBka9YQ21jQCGFgt+3WPp5hpqAlsA0mFWw1+lg0VHDXGOLXweE7B+qL
SUCqXkr6bRaBYRLFJl8e6Ka2Qr9aJuzd6PvMO2cUuEXOZk24XPrgja8kl3Xc
bRFFniR3opjKPTXRNV/YfMabn1YAg5OJflcipoHCex3x/DztmVtkt+N92U5V
fhvCt+h8xI5WMGpuZxF4+MKeFAkxkEN8dSxkbwuOM923gHRxzDqx49R33Cnl
CfnhN8hXB9yEfnuPgD0LJXXFDg249GMsm5ODsuGFpc5xbSjo6CQYkbJWv1GA
4Q46ptqA+94tR8qrrKTIKT8I9+lUxY2d52IE/eSIfpzIvzVddxwq4gpxmBni
x+xJIwDYQoawFhwf9CK7ytFrpxoF25WtkS6aqwgQD5TZtjC95wQPoF+4FKv0
6Xp5pjtHcqesJkjo9fsBkdQCY90mS+bnZ+arks+fCxeKmRFoKtnHQdiKW4uf
JFA/VJywRsZgZ2vSOQaewKu3Ap6Zz2DA3Kd7Vb0ndKqheNCbIUVNb75PXRSq
tD0ET2B1tKkRDLtuHlcbXTD9kZDDO8r4TeO2891uVdSymlhdTZVgS+0FGc5B
AByIaMAZQ0qr3AzZvUaLyNQsLB5zmsMkQ5qbyUXu9rUVVueKKy2E3obZTA6n
SjSNwB9zkznRRfyxz2EqAy3UN2cJwwez6Rm4LyRLPQLbqwC+Oix3az89T3GU
Db3rxWBmYVVBiuTH/FHPl04LGLWbMf2ZxOc3Bx/ffrglau9j5sScHaBZa2CV
yd3Gp+3DGrpzgkftgH1ZFpHBt9OUtzV4epBLcEXBJQmE/4ULaA1s0zirq9I0
boACfXdsnBHmMJ/cHSOFl/2ajxX2rmRx9kuzzdAkxmD3AnezztcsWlwmlao6
ebEaUXdgU8n0QoU4bCBfxx8sUE8oowljTtg1WBTeeE80lb3TZ7XY4bpk3Gvn
TssdEw7ECAHfoB40Aud2UIQkRKAGxBK5Rl1ZeU46mcEW4ScpeqLn6lsS0FCM
UgtKW0M5lrtuIe0B2UFZRqAidVK8kHSfplBk06pQC98brR+wnKG8klajxYrK
hi4CiI+jq+EH8DH2EHwUWtqr3Pt4WBq8xstznOi3Un/Vdu27TeKmafUDcrH3
ODvfW2FFleANDkvsJHg4gj8NwC89wVGJ35lV5rLgf4F/WSSO5bnOvkxeH5Ys
57pOJAmOfoVCfaD+3nxHpDrg6f9JlndyOqCxQsqqmmn/ypogvo2pUwadOw7G
KBM5i68ZT7d7Fk8gmgPPeogcMBBTCerga1NSlbooTu5GALtmIwjZvBbpLVTU
cuqI+bqL23QFMdDuYdvhM6CpZuWEa29Tkm9t+UhR1Wld+2NsrnDKE8GVqeaG
ZMGWFqNrPNGnpVfp4QjbKzxsiA9lkNTb1S1t0961VPper3spQdU0dH/4Imif
cPLZ+YnBvq9ghBX8zQsjAE0Kcpvp2wuAwKfWv1FOjlFdni1qdeOZEVV9iw8P
f2gvFVzH+Uw2ABhjqeFh5qtI287myJxKG+swfmHtmfN03qjaC4TGNumP6Nqd
vuhKll1X1LjeXkTMkRz/XIG0gWLRIKuOg5mEX1SnTHJFP4QtcGfQXd+vK6eh
rg2M22Tg5kNeRzWudsh+Kzi2JaoDLgF/SEs9xtQxkIkQL1/0awGtNPrtyqMT
LmWdV4XSVNZmKOYsldvmMCAVP6a+6oo5UKvdXfp27gFSSS/rH/YyYOsbTnhV
KCMHmu3eBb3xZtVJFhjg6F7fKw82ESlQWCk8hFz34ktMNt6c4zNNIIW3GNX2
M+0tvScVTRPYa7pDC6OAaeb8ht3BhuypwkZ7yCcJCNihMiwZOPgnIcOcLsHF
EnnH1nOdFUqtsfVNXbwMEuJ685yCsznKLncM/I62GspMEdxuHHX3qSuc1NpN
lIkJ56PFUVf5aZxE5OlwiH+cyo1YZqKZFcn5bKFkPIX1N0smiNXe/iX1Opqq
lIYzmZomw7lRGFJyinc2ETh1Wt5VbHWb71GxHZRbi3U1ONqI7uCQk4fKhh2s
r7HC+/Kk6L5Y90dGVVAlaOiRg+v+tbtO+eI5plnBFQHVoFTBnV/O47lWLhmZ
GHmd+5OXYsaIXKl/t6GvVvFktyeeIvNW6L5DAv5ng/lrhDWBt87SJMyjXAfW
AZeMnLG9MSxhViNst1ClhqeLMb/whOiKsuTBVGvsaRnV3zXOP7P32Lcjatn8
XTqvcX2FAJTBZaN0cre+4EbfZorWynYWL/qPohWIOPs9Twmvl2y8qnvU4xy5
6itP2pOtLR3LT/rrsZaxIerh81A3SaTyWG5ByN20edOzP98WJ729chyNd+qi
3rYiNS0yr3C6oZ0gw+bQ/GK3G+rZtXY4RuboF6hOcwNJ0LVnxjIhYbO0QmLG
Rgw6k+DqjsCMoygZUb2qvuSqwP0I7L2ukrDqt1xIroYnmNhU9PP8fwQJpBLI
2atmsqXaYX+MD+xNHBhU3ieCK5/bYtoPZvwn9ej+oU5CgVWdjw1urdQqV6Zt
WiHYwXH6xRNe1CnN7p76Z87XA5jHmfgekBvMNo3QiC5Y3D1KqjECfApVbqJY
apvvmbYX83PllkB+pUAVU+Ix6lWELW7Vj69/Id+mdfFAXfCPtvxxHNXEUmrP
IU3GgOY+yvRLDGpE4k5LfRxECZnIF5WxEec1urGSQeQwQJvWVaXL1TqsORat
gqGV5JR/AjWEqd5CIxa1ieW1ZKNqEZGUltCoqOWw1bAQym89R4tohvjeLJQ9
IZ5Q30ozOv53yqNpmiryh8lt7oQ+Zb1scdWxfu8xyvp1NdwDMCz9Ivyau9q9
lXLO9/PpvdnfK7GerP+P+n+JGsSpCwriCAwOC5w+isG8fjWMQL1zQiexDnxt
YMA67j3dcnWv8l7IHGkx0/eKc0FUgJ/xpRxLKDwSTogWmgBni0OIJt92LTOX
BHw0vnUyF0//DixRTbaf92DKkE2LqPL6IsaNOq7FCqdDxZn4BK8BVt0N/0MO
oTjKl0ZKXRha1Eq/E/Ih/0uhzhonixz5BKSxCEDq3hBAfyd42uB4AVL5BP/q
++bpzqN4HY1BNjv8ztiTENpArusixPorrS+YDoLdEWNhafySjxASdykYkCoR
C77rMc1UE25O19TMDXCVtxzzflxoIcT2fMs+WQGiGqBfWUNlW41Col2TPJyV
Ek6TatKuwY+62YBLyMZhSdYAweqg12ma6gP0Fm6m3zAQbpeB+RKy8ZQWSMgZ
NqLTkfUvwdb3KZDwmTyLr1VUhmqgMlCNNh0ZXFxNyaxLVtmnz0ulUmhknNtz
1gG02srj4hpky5BtXEhY4hiPApkJqr+xh95V18H7LUKRwrGUZtDMyUi2d74v
v2qlDCzWrhuDNzi1w8iwDoPaUviK7KMKenmLEbAqPHzAEKGRsWh20DQu0LWu
m/a4BDCYkUNgeZjZ5HB/0KBhpiMUfxfHvA6tH8Wx7KlNJypuwVfe1RygOsNh
KHtNx+WhfSNTZADmGO0NfAdSjIqRBWBTqZQphPAxnDHBUDM1JBDVl52pzokT
X+FVRlr5h9/eJ9TE2dyphsQfsfaeaI8y6+vXyZ4Rddb/f19mxDXacRZcLHhb
rsBCRUxq2AQecsN8henn1OHZk+5wXpmT827zww/sbfAnaPKpu/A/PSVk8gSK
kdMeCf8mbi5ivxg6/9VGNm5A7sxbfHPk95IKhf6aAZaE2gFUuhEOyOqNSqKy
436UzQUchy4vqS0OmhgAU5cjLncQWx/2uJWVJTnJKYiSXJI8UZzM3aEiVgCh
JdiNFMEwR6x5q3Y5th0E0Ubx0tvYcdZbUWtwK+vU8kNesCyLKiz8CaCIRRxx
Mz9PpaNfnjTePTPFFzOESwq+FArQISYWXt9CMsW7W11WPNorn1xKsDm0cNNc
jqJ3IQUU4VXAEbmE5NgN6TnSnX1d/wz/ZFBlxUynf8meseEDWBqxLOmGyx4T
ICkV3pGmjf0wQpDli6sd+WnkewrtQ2QMzJcLo48nc6UYCSEl8RMROb1P2H2a
qdqxGod5KEgnbHiuc/jsmF3YanQBjhzfJFnxz8QS8G99qDk2mBmLQIjhaWvr
epHA9uOdwGK+yRHBmDOMiYmEtQ1Uz6kPWJnKhLxXVWUd78WEdzQ+VkduPjqK
m3o6Ug5c4h2TAKHP4oVfOSc2TJfZTuGDhZtrn0oSEI+vEW6Hf1cjeEM5RAcR
DG71rI2/CrOcXYJFm50URTVHogFMJKQ433YAuKaL/NErBwZuJkZpfoPz4qco
UuX6yGJQGAVZhB/fQ2DzvazlZ+Nk0sQib+yqz2EqfoFT4nnK5WQ8TPDTnXqv
gj78xbEQ1FkEz/wGfToS4EwQdVDrzGkDOK1eFricJCBUYACyMQm2QZBkdNZr
1IDm42PzHk3D3Kw1W8xKnqmN4LZHepQaFJN/GdJVjMsQnm1ae2rD+UT9kWRg
qoZZKa1l5DoFpp+MoKwpGwRdFvZHvaZmFfZvxwJTLlG81DiG6PAGNLlkzWEU
OfvQvHuRrT0O2t759im0wxRE/JdJuUZ68eiRdZc61H03Lw96HexELklYsYkB
G08QbEpY4h4dk6QxcZu4v94CR7guc1WJ5JVFnD/7oSmLAqJnxhUOB1puUN/g
ku7glshTZsFrsfY5dJcCJocu4jkFQxtupvQxBi1JZ2Ka9pxSO9smSOG5Wc7N
GLYMWwQMe+oT99fO4WNKyFuXmZrLHbUSCo/bfVh1HDHccXnUdbLHUKZeO9UT
Qt/bVSNJv8K6gLLMSC1M4Vmq3Z07bSc5MHDEY7H3xnNHsZ1/4mfz6Al0ntLt
MLOwphVtwUYW3grdXZ/sFRoiUq2jBzAdZIAQ267IATxgaESVKed7xjAOx1Vh
baxDcI4ZxHb5W6nCgIJXN2EXgBuY9yY7WQMs15Q52nRlwWGqDUx53DFXg1cw
EDV1QQnDp2fy2SHmfwV3MgC/IZo3UZndlLlUdSjf3hk1FlgV2bLFr0FhBPtb
YbZL9Nsqg7v0sdMyYghHl8r7yEds9pDzzxqRK0plSbhJbQajes3t76uix5s7
CyUsAALMgP02oBl3azjB8uNVYWs/GXauFYFnDZVf1e3y90uK0ajHEYSDyjKk
kKp5+Fknh+qJJXa56HJtVEyBOaIafD67Rs/tCBBPOYfLa0OReel8e7w3A5Ah
A95AX2yvVyNQa0EQYmN1gWqoVCNtrZQ536/G+nEmGPbdwuw2ksqH1ocBezdL
EbIVgH7dv8ZtiN70+S6ONnHtK2Gac2Xpsgg8dQNp4IhD1qD9K1lfWP5uJMrm
z9v6N2yDTYReJH/KU8S0Ab6R0nnr+z9VNwg2xeD2i14DiDbr21bLOj0SfVYE
bVivPiIwnE3caWf7E+b6iyH6SZe5P6obxSwn96vNWBsfo5ABVLaJNCSMF9Qt
463SiJhFaJhwCHlJGtwy5f2iinO5vKTOQZcHOr7jYlS6MXZshDa9hTfEyjUZ
rTTQqlSARXA8b7L9XvNE/s1WEBM1tx6dkxpph8SuLELanGfMrAhtD7V7WxDR
b0+0uN6eTVAYe8gqNxIEhqlVTP6MqQd1aQPc2nHQUNM/rkI6E+jnJ10VRg75
kWTBy8eCp6jBYWl3reQuz49a862t/bCuzZS+EnDVifB3TOB9dWyHvZZbG+UI
/KC3SOIw95fpMEbfBO+0K49tM8vE0nUa0WCjyMw92raYpBNHVG0pdGW4F1Nv
s1MdaVkruPbbjxqPDhPVgIrAn9xzyX0Rl2mYWqPt8S+7yVqVeGeRLuqnqLT1
OgxB4oAw1O+P6Rc79PpLv5qdAOfLZAzuLLLYzlSvLnqqBVLUh6rvAVC4YIgI
nipKQYptz6NNXlwq9uomnjWExcG/UdSud4YYkpHDm/eHT/mRuo1DzUTWoYOW
oDMUiYREgLQd7U3qS6F6V96MD9tUDYvimRODE9/Vfo6R+1soj8r/w0cD0bcm
cM+WBjKRTORdAYWMU4j8otslpp90+lHJwMrt2fA7kMU6EDadRac3Y+2bBMKt
X6dSnPxKcJlm0pE3KwQKmZsdeh2XTAReJI+rwZBHS88xrkLBDmg3i3t085o3
kjvhPW2ksFZ2QKA3RB0121+VFK/fghuQwJkRay7y/rWlWTOfP9M0YwVp8+Vq
gKSpvc1iUeNr9iR/ISn7gguUxvRqAluCqN7l1YamvJupuG3Ua1JFF28OTRpc
oQ+8g1FnrDfswmque9w06/mS+eQl5fj98hrKmQHUvMtofYTZx+D9uAuhpx1a
TBOcw0wXusJV8DVm0BVzbKpbD1QuscIIJCixkKeETPM0T+ke+e6QU3CNY5+C
QUCTcYf3LwaF/pJm6Ui1/fw/SzQdqdwNR76nb8vqxl7KO4WoYgELtVGU1+HN
567TXz6WXyoN2MIvi95If6LbsuR2lONRJoDIACY7bWuHkwK103Nrdrh5njRr
gyZjoBJVIP9rQ0h8X78VM9N8m1QstrKAYstL5G5XZJjKxVyC3S4XQyw2Kxqn
azNcqKWQr6ev1wIwBAealwbey4UHevr5COb8nFWjjE/d+i+Xf1i0UDZPomeG
q0cvAUmBUuGI0bC3neBnHnec8zPBa60RT1O01E6jtgpwf9DhAi7DN6+zwyQm
SsXqonED879Ta73qhT4OWir1AoglO110gLCaKmmwi79abvYAhaDzMEjGQE3A
mLNILmkr5x8hpJmK5OIdOKGyb/LUdWwN20bWR4pMTA/RKaG7oi1ABKw/gQix
IW7+pZIfuFz0L+qnzFjPEsjtkijIwlxl3CwciJ7qvMWXdkOSJ2J69IhN9mTE
YHrHieEOzcLT19hYS/Zsteh5BPPFDhf4WNzp1ELsLC11jVwWECmrS9/StezB
EowoQADKxq7ea+HcvT1puekHxE1qpwwTky8HxeuFScT3720nDGuyo5HueP+A
7huK2laYMbTOUNkkqQatvAh3O3RTg3gl9VV42sW8J9pkWytzVEwu5RGsHTHn
9OYzLIeOF/lIZqZZz53V4+gWpStBNtE8O9e0U5pYjS8S0gBX8nWLvtPx9DB3
89bFbaLIAHL/rHK/vjvU8gFHmrlUI6wPcDhQS3V2YSHDR5MQCEEOgEXz7Vnb
rZJxlIJvH5wUbF47Qg/d3hyNi2srCwwnuXuh1IjY+BQRsezkKPzuz15gNkYH
1//GjMHfg+XZYyTn6rFxTXTjBExrzzH7uLpBU4J2RLBXrdzl7GkXkc2aYqLb
wgTX+0UnkUe5Km2Mh06fkKdpMkmKxwYuSBOuOE1Tf5JupqV51HtwW3ildw4M
PRkbkTzCLbxDhtfj8ZYrP64DcTJygs9x33vSjvcTwsK6heHG11sz6y9nCYp/
J3NDsFhF8J06Xvk6PQoSE/LwB/FVOZs052DXj1ZpXHVsTwR1GGVpKSLg985U
MmMa/jOraQp8HpR+i1wjyjleog0bC8RLMvfM0gAGAecWKwJjY+exNjGi0Xut
ZQSWhlf6QMnDnkSpGLHREvjIuS1V6SDKe7/UX4yymzonQBaKyPZcRO6VTKh4
jp2QKskq68YLvV/CtcC7NPwbuM/A9XMcj3erweShZqxVZdJ2wZ5EhZmz/lva
k02gKSdb9JxvuulRl1q8Ngd2dYaQ73TVtiRjaMjlass/o/KGwY/c4vGQbuYQ
w1D8+cRmuhE1kbpNKLOk4zu8W4MlTpc3A2HCjgzW08rrni/ZF3UwCDGsYHe5
EZ/wTsPezLTp9dv6woTGi05X7YpHvlh/bHy1VMr7MYjFvtplWqtINARa26Yu
OMWtT++y4dLCe+7gYE75+thsX72WXLe4v9ZgMYDrPUOdvXTySLpTM4j0/3ic
+Eo5zQ83XM63SXuefMyGWSyTXGPTrPc0H1qrYHlAYdbQwj8JSpw8mqnp2c/e
DpHc4M6n6wnhf2uaM3SUchQAe7RyuOBfBQfl8mCPvHI9FpfG0ouOLZgZ60Eg
LQsQHEDtIxBjj+jKt4JxI5j1UHiKFHeEuu/IjPPA89SNAerIkkWHJgMlS7e2
SScK+D36PtJQR5yv608G4fHFxunvJJFo7cabDxkLpJK8ffcyZFj16L7CwXsi
g9ZAAi1ow45wiw8mOec2e+Vs1c/KheWG63xy97QfRmEbxn7EhzbF9SXLG8pR
0aRMWA0TXBeUX+L7LdJfI3+oVdsjJgBdvWDQzjfe/Eu+hlL+v3eB7cEqjln5
viE/+TQAzvj1y73KHYnd45w0f4QjkZZCzh0TX7twC3xDfGAsXhNaCkuOarEx
D4KO66EuK+qPa7r9+/Wv0m34MBTMGcRfYcg8uKSrJhPA7F2dICYj8OngtjRr
T20zXGcqEccdWBULc0RNffh4kPpzUIbEF/ctdxiLXvRDLbI5km0OBlhPQW0m
BujO4TgR9DSk9yHlaUEmpuiYcQkJDib7M3zZCwBoCgRJMEWY/vFi3HlP7hlj
qVTRR5Js3xXqP/RXJGkQKddgTl26fQ3WsgGU6lLDdzMRLCS+5j+hDUSd2Bn3
HP/6SBpp3sLyiqgOsPMsoGCJsckiiwNOszPzjEY8zm5UdwfjesAnwQQuY8X8
QXd8Y6klz2lJ9ipdpqfJ411yD7GodwA/OBrVs11m0dqJg3T7y1WExiZw/4Rb
pdhpbt8iiAHz4pm5xqUwvTdnwQWyUiUHMG1ejiR8B8UGt2TwLQ+7Qp2Ox+c1
DcPxRZLEinLUX482Gaa5oeKE7UK/wNRPh2Iw0lyJqc6G52ZTanlQ38AOTmEN
aLaV+SoSlHg9LsKfSL2WnVf0AUb1bP9RkvLcfxvSaOXENcvceylJDHxP2SXg
+1kSjHaNEtd/mSz9RVqOM0myqifFZfeq+PQriwc/mgyVLINjd6vOBIv7h7FM
iucq9wQhlW4Ctn6934iaSpSeiMZ9Buzrmcc2wwGy7R4WMwIXzK5tFfxK3v7n
MQA1laYHfjLwb7AIIytYviTqS5NR/WuqS/kFTpkt5OGubGUiy4nbQdgQYhtP
fluH2ElHkh7KVpWom/WN2YK9FwqmHF4QcNA/nq6bxxaI8iiEMDOGmtH29yCU
dsDttrx+DjJf7lBFAsTb0Kf9B972/7Q8IcIwO2m6C/0Oq7t92U3+BUE6hdsE
4OKL8hh3iA8VVsaW0/PQ1YzvqqsnxILEqt5U7QK10bAaGSDcCE7h2lyhLQAI
1yWthRcjLEtr3rmxwQstiquKtdBH1DnM0WFLfGeEm9mnN46OXbFqNxTffWCx
9Nnke5tk6uGGyxnbp8Z5IkGvybEqLV+CK9uoucg3Wkz5BeQbEes0jYxNq7oI
+8SIlgEObc9qKpHBHmFxJzzzflPGV8dwfDg1QPst538fstJVV/O8SUkaUwV/
dxnp3qhs7EkeIVXQDxQ2o8CciQqf0QcjT7FOr+NxmviAZ0W/q6bA9st08Zvu
z8oMJpwEItOxPM6ocyCQfNjLmAE3vooHmV+YGMsRNUWVaDXn/DNbYjwXb/UP
PLbXXY64HYbjMRMlJkF6ZMXOyk5gW27D+S9lVmJcETdYFbaLInBfLVO3HP5x
G5lq6noLNOCI3mtUFHNTy0mcb4MhjoBqpAxnC2+u3k5Vy+iJtZODOhIK29yF
SYU+3z0lm4EMBn9h7VlfwFLRTQAFNSGCYUCSqLEMMvkDV5e/49RO7WjDsi9w
9AZp/dslGpsuKJ+nKOZ9B+xNCY+Kl+U6M2924oCulzgZOC+7N3xpedHfLyfe
gAo/9OW47LJdDWlIDec3an4Ff+s0Y17Ou6U8dm0QjhTKFJ3GGq7fHyZzpEan
GYx6qauJsVRa/KfxL01rQFW73Q8OPf4IIxvnPwqS+h/3p+NjTRWB9+S4/ewn
IVJs2dmNH/XWTrFIP3YHJk3knboTArqxjIqVsCZ/S5UJnD29mUlC024lsIAC
jUKLo8FIWN+jyblva1MWWe2YfkSLNufwBw1DZqA0XUGKXgN9GlMBmZIivlwp
C+OPUDqDPhVrLFXFzsV9iXIb5ohzbY4RVNbV3O7Fus2pfURoAf6NEhXJ2GA7
3kIxqYs+nFsITQSwGRWeA8/0wga3W1iLjK+DaUGY+aqwKWR1WG/s6OV5u5IF
E1ijj6cFHOho9o260gDgIs2PBunvhBGJ1nNnf+RflKlv+6cLNQXi/E8mepmY
l6P718fNiRLx8MOXgxeXqtxYYv2/nk2lZF6RcZYt+d8xMfddI2c3DoyYwUwY
f3h0ZRZzzIdKejnD3tbSK1zJAneaRscRtDFmV16ze/fPaH1Ux2Natwi1qF93
uX2ovzKfugIxwvAREOVh1R10KT9fdD6E3jmEIq7371HxS6Lrk3X/XhjoBlc4
zrlq/5a8sRrrN+SzVx8w67xPd4pCwJZJvqiKPaxAXF4JmyHJKeeCA1ulwlFR
7ReV9/uMqM7bGCV7NwH4++URqDf55Fqo8L23vipYQb/P6ay0hAPt6w+A/m3F
KMgZNjN4sANoFinz1AZNkAfLwMI4+j6zh0Klc6Rc8uEIlfWOyKzXPgqGVvVw
xf5vqNZ0So0gE9HQVHXc7RvHcO4GOCXrBndVFMZSiQ/cozHNT1uEkDbHk4vN
mh1NH6wy7sErqihBkakLdUjF5SJ/Y+qvhnWW1B8TFsfYTqR9UDNYM3y0z4er
NEI4Z4ztnYtVrQmiDJFLHJZ0PQ89PjYcU1c+DUZI91oW1La+7nVzjShFAoa5
o8RgXebswzVAn94A9jn3s4INw6WFuqomNJXxLX6vjyeMEtY4IKsLHc9/HQ+h
Szuqq/By2iTj4sdcq17xa/8egj4smCzDJ87IwnxwEKlsU5j0ywR+DLZFXCKZ
DFlWi0I+yFHk3VEaH1kt18pvIB6kxCmlxSTwfbaWLrUt0P2r2teZHJa6brlu
TwuFEl8CIJYKIs7Nura4RIO+hY92reUbomPKmAMGasTLibS5muF9FvdtitBu
taxOd98Nq1eqkD/Nh8n0M62xBYDPt77fcbqwhywGxxftR/W8QY0zjL2YUWhm
1k6KlvcvnCrRUCFToH95hcLnSjILX8eYv0FTqKCOvJUGwGS460Ho6oDr6u5h
rnDWense4VZ/4xB5G7geJmD/FmFeDTx6yx/F59u0EXlMobWvoZJcUzhhI/s2
Hh+tkwmlg6QIMW6OV7rAqxQd1YZtPsz2fufSMqg4lzF7V2km+nr15fUZ4qB4
/ZYmEClOSrPMwjuOvyV3hLmRiUeRDGS5+Oef5jVfytNRFnDl7refoN/24755
cADlGYCuh30CNwRzYSa05TALIOjQiuJ80c2GaFlqphXKb4hfbXK2u4Kovsik
Rsnjh1M2RUCPzoZLp6mlDcVhSyb+YArWxRNYitdAGXF7Y6aAo6gTB5v9q14O
sVLrJI2ZFbtg2av2/BeSXrRbG5v+ogeQHc4xL+niN+Sti8S/AjKHjO46N0wz
fCNCrLtDbNurFsig9JcBztHC8Kvnm6T8cCUzk0tJD35TL9lEVe5eqc2lKFo5
nv+vyX5BcC/ZFNWcaBabrY9FbbumFhZGOUB3DyRp9uSXIvV/yM8cuW8RVXPI
+yc7GnGT7vEj6YSWvzc2OrPgatO6LqlLWVsFlsRLLO7ljRwwO2qMrFMw2Fm1
gU4QhDWqyWMQy4TsQGTT2C42ESMhBRkQKP1/PBjxJH6EpcGGz2GcAsVFn5Tw
OxubHeiFbzWLq9xytv5QuFSM1RgG3MEm3vUORMl/eWBErADZ4xULYx8pkI8i
GSbWErZmS/nPdr5NsXOVoFs5j9JYA8vrKIU2k5QR8/PEMxwI1rZMo3XKJYuM
nDEWBFWeSbVgHnpLi6nNSczcwb/dOe3+B3DMiF/uXhUr44KfXTiggNp8l5WH
ONCG6K2AvCYNsTOsmeWWibO7f7NUxYNjYt46CvHqVInr81utgHu5FjgC+n3Y
JjLgvVD/pvo1ATznIbtJqkwhENg7v45vdOWeVPPIBCD03Fu6bj3YHlY6bzNt
ErteFBjSSJoxJs/zkTUeS+uEREo7mWTqyVMB68DM9irA5czS8l/YycHnWb6m
Y+I7E6IwY9pmj7se7dhpGviQoEZFLN/oKEiVLsw7tB/52Un67jCefM6GLzxu
mrsftrJQS+HMhsEDMgi+Ywz3KS1HNwGF00Y1Fn9N0gSHqBUrNBqN3eINoq7n
Mo+a9Z1g3oVYpRhy5RfB7cd+76y0t6WV4I2BttnH86VweUo0SsrvpPrfLgIZ
5JSXXu5ZlclIeOGb1S6IHEj8GaxKlczk5sxGY94V+IobnmUwkMt+c93p3hdG
1+PTwpmtdu+0XJtBT8MoKqvHle5bl8FoGQBU3GpFaJz4ERDxdHTKbyXu3Lg/
s7EDs0zvtIc6mdK7xreei70bMt4f3H6fUD0hOnPexGWRQn47KtBxdQRTcRTL
IMxEgjwg1dBUFPajaC0saXAiyTplhvv2lw62lO4X7MRjhzlU9TIZQk6SQUWG
Mtq1N6JzHAWtbgupRTNDxyGOm7qMQOKV1mDpkvXV+vlWCcCD86I+sBc5ia4y
zNq0737IjDjIy8DjLHuYmm5N1VCxAzZjcK1wV2PhaSOJPCVeGxFCZ7aPk4KS
xndk+TacN5W22I5crojZgGRJ3HHMAdRnY+jcJaPybnfLgwu5fsC7tstKKk9E
8UULzeyw+TSbyZLjT9rw6dcDLASHM6BEh70mP++/TalUCsYCnaEFDPeUyfmh
J9PYkGqrieHYx6iML02PYVDiRiWRq+QJoMzZohdhcUzcSuSUjQRqZH1yJTWN
HHGsuMsNQ8hiz/IECGcoi7KIsQqRhYleHSSkuBnpvKzSBKy7HkZZg+oEhOMH
gmw5xMxhFAMKqK6qmyLf28wfAG5aJtCCEWa5p758eWC5Xdk0MG6izsKNvvP8
Cw6eMn7p0Pi6XqxjC3oSJW1uYz9M8HwdFvSKGEWmOqjSnl6yvzAD4f0zqLsM
MbXHGZC0rt1ERwuHxy6U95f9f2cAQILZl8oprWVNdAifGYEf5yxbZoCHFaPB
h6SHae0L4JBZIOQ/WXS+IwhML2DLPgLE+zzzQAP3C8zKNxM/N7pUIh2rG7Bs
MXvD/8wIBIjxuoSxYOGR2nrEH3aHr9sVk1itF8aa+ol5GUo9fmSW3s1H9vgv
yNxHiB2UJjx/8+X602qumFhCa5gcPNUOse+EVYfxx1jv7GNQpfYJnI1PzRW4
pF6TDRt/OYkShzSBbmuYzcuyN+htLLxH0EbMXqU6Yxr8P0y1Z8dq2kKnrJ+i
8j2NzPdlA5xe9o3CfJsUSLY4vIhL+FgDhNawKCut5gI9G1iq6mcu54drL0Y3
vWMec4dzsTr7nB/cff7e0jy8uo5SCCcwZCfEPNrcrzHZDhRwDWxWoJD6v/1J
IlrS+dtpqeLB8s21R0xpgsZ1ZMA14dwW+FRvwkrL4peXR6EdW1Hq76oXTJtY
Q+2JzkTNZSzM/uC8zKvZ1vGF/oesE+W79vy7wNfGgxnY1HbNfjM/6Qv1T6f7
p6fgQQqj67kb8d9uVQSsKYDR4mA15QSrWlBA1DreGDYg9wbBWCekGELoJraZ
5LI8QUvmQE9pZR/J5sudQql0x9hVOpMFxsg3GOfv+j+4fQgwXQg2pVT4StEM
HjEpMFnJveAnPlVvxiuV309K+J3iMRyD3myU1iy7uY7eAFQv+VAQ9nBFcW14
XobhRara/yWJvh9oFYKwNzLD2VpvccMb8tsSqMgknv5kPCIcWhAZCJruNTOz
aSfzyUb2G57gEc8w3o0CznfviuXqylKzPmv8AGJtst8Bap2wrSmozVzoPWds
7cMwqka8e/GbutwtkWDcrnDgJNQfokymE5CyKELCxRp/VDOX1xa6eS02aB6G
8o2T7ofMs+QFJ1CniB6EHlTS5+F052a7ynCKx5enwiZXhSnvdAjqaFo5j6CZ
S4SRXHEwHBCFbRtaq0tiT1NmOX7XtOgf3+9DleNIZn23omdIMHdtnBqCNkck
V780oDA22LfVsuFHjKrJeMkCQXoUWT4KOqb8GmhINKkk2glivPHTE8sw+fo3
NjDCYQDGZVzCHEJpWndaQf6luzD9s/Sp30RoQepRUExMpds+tf4GN+QYjprg
RGmnC9Et8vSbSymVR2A7GOvKqhuqxXGBYm11el/37GZh6tVGldIGtFfZfOlE
Kkuh9TqHkR7v2nA/EWq0G1GvGz3qFRMHcsPqQsLY4cuLbW2OQ+qZ6j6wyABU
Lg0+BKDaI5nc+TRJF6yhjuWY2yAmyKOldVWmZtMpInRPaKmjWCAOZdHERznv
RUgQHbgHnvMe/AVjmQQ7eqK575lt85Y07j9K2fxhGVFtnQNWl6Vbn3BL6Hb6
src9zLHIFAHd5erCx+tJyZ5sbrwSNc7AS9FUsY4NmGK2WquyWdCieiXKMZJN
BSvQgPY+FIPlxAFH7Wq/ogZmHXrVwjeeUsemGIRBqZCxv6J2BBHD+uGtPOiz
qHnNtKZyuq/AEbGKzCVQm17g92E9X2R0c7r7mM8zHUAFTIbmgjHLfUtL413M
1FeMYilvd9IQDAFSpkXeXaYqwszfSN2oWs0aOzJSPtquWDK8pubhIw/sybjA
I+WJ8oDvhmlPWQkQWctBJHDLELVjBqBnKenWgTTkzMqbT9DZ+dGeaJNommvq
eZTz4Tr0ikRT3cN7Un43htm/laprBdZbI+ssuWhJ7oil2c3kEPQoxTw8Larf
/svGK/VqKDQGtWECWUQp+9nrd12pGCfOzQZyjCiTcUp9dYPOh2CorjZQxkMm
A2cDDLsj9TIikPeNNokAOnpy26S1r92m980dEkAF3yAFLJVzIPCTDrEiUDX7
Kdlo+arMf19BzW5AxSN1yEJBefvQg/mdbZj9I/H0Ed8GKiMd4M/S3HnNlqlt
v0I2/DPXlJbhiblKC918AQbTcT9Xuk3Uo1pUhdRpBQaIjjsDiC3i4gHaTd5z
NBHS10i2pORDlXaflcq5wT/Kx2OehTdkwaBxsiBp6pZOw4GA/hjXlggZ2qLk
ZBj/l5bDyp7eb/x5qyEb2ZzNUEJJ/6sy+hcC66Q+Ve6/abPukcmiZ+QNYmYY
g7MbRxdQlDUyM6Gxb/wwoPEMoqoG7eexz6KdDDS9HYfyP0gfmOkbhKIBT9xi
udPQ51vkQHnUfRx7yzbqssSqCKaw8PVqRdcYEmOJfxxiTzYOiFURKnOTkVSL
yYJQv7Zsa3A5N+RDl1JFMoVIkqHtrt7vX6Sy1WPZ0CDz6VdTUiq5GBjNhlTQ
IvUuVAbZanqJU5eFcVoX1xPx3esCw4SXun6UMKNCaTGoQjh7DwCMHTZ3dEvd
XkJwn9EIHsA8f7pgwy/320aUwq5p1Nl06FFqhRGiU3u3waocf4EXobyWP2tQ
W51iHCgsCPXNPMltzuo0CF+S5gsqp+12tSgmjeeppp/yYEY0+Ij61s7z5MX5
u1mNxNsn3gZ+z93B/f5JgW0aHW9nDJP62YjeLoU1QvJ9QS+VnASApLuakrs4
Z4Hd1CsOHJKUWcszeR4nIKv5Qy0oFTnGllSdXY+5uJs5C8zgTKCm4CBI1HzC
lqkW2jHAuU+Yb5RFND02C11zuMXjBjVd9unzdEgxRlSR9ZsWpCp8ycwHKeAI
3TmIz6vy4QpcX6XgXyPuBGVY8fvKeNLr05FC3Gf43RUm6DI3MhwIo1gNp1GN
7x/1GE3SoNvv/pfp0ldtcNc2Jc6icPjE+PzYs2wmQbWX1Os4lUt6iMv5bMJB
73gUyOKBfPm7BQY2S8P1mh7xM2sDPuwmactDpUMh8LUE4u0pgCvAn/r30s+L
9gwOH8njnJoMUjrkQ8xqGmb7lyhOqFO4XZmePbMy42lhMcARVsALJk514aaM
NEBQ+odTCKF9WCoG9kkU6+Pozwl9Rkkvao+INZjldhqVzT/mTShXt3YCPxpv
f3q2e0p8YIffMy32NnCoDf3om+csmzNqFFhbSWfU13Jrta0M7YnSsPlpd1Yq
3lx7gVHVWNDYaWVr9b8fn2tt4Wl2l9U44hkSSiW1ixM5jEtFEJ/aBTKxzU4h
ui0Fajjrgd7wKLwFVh7qLtRjIzydHrX1ghujrKDa0mEo0VshGBhfyszPg3G+
V/8GLJ+wQapTUdrA3LpsEYExTk1wePGYHe1sLDqhqHGG8eHLp2yek/+3koaI
bwbJ/rv1TqyLN09me0Cf8MYU3attsy/XiRrzZLDurDK+Mr0XT3/Fnd2QAt+B
i2SwO70QkD078//W+pTFZVCq/dn1UHqMlIjB1TgEYcAaoxope0W7ZIWEt1rU
MUCnTAVzwojWpfDXMseXen+s435cnMW0SBqob3UmRwuQtpoc05YpgDZHCvxC
B+ZQu6K+Z72wh07EtDfb/dfpFO0FfeBSiS9FwYaxGQmgnPYYqVrc/pR5ntI2
V8LAhnEbQONwD3FD2CZYasaNOjvzFYcUfWLZCfM1immXyF2LNgXTKhMUqwI8
APmtMMdC2jm7S/TZAWvmvkHBPoxuwRVwPl8RTuI0kgPLky2K/6khNjlQe3wT
791fcrMaNjDgllqCP1fWT0v+QFCHAJXNxQMGWdATBVAuVDY4tsJvNB45TqVb
iMJ9QEHYHgnSNP8wPs0Kw2qMikqO1IzhHnIr3irP946j6jxURGJROEJ5H1M1
WE2E+nUF4k5sBPdfClUnHHHEYnGoBOgjI2pFPKA5rfnK3OENdROL6xk0mL/5
NYq6vMhbPwrFETAevziuqbjUUXfYOtgB+6QKK0RMn92tHv/uaDeAs8ehYZxd
TXxKlQNmAtHqMlsBiG//Czz7GQx+vLh1D5drRF9PzPW0MLjycxILn4xnqWD5
ckslcYMrtSX3PdUdF7ASR1DcrNVu7b2rQX6roqfCR7dz8Gh2cdJpv2VgD8vJ
Sr3Tjo7PdjllqopiAhIN5riSyhvq35KQlxqW18+y7p8PMNRAMDyzxOa8US5O
e9pTK3whMIn/E6ADThC3l9pb6FnAuce1hChB9FF5XJT6wioHeonMJcQGgmBk
Idh++lKEIKXfvY0IHXdVjXBe8fLQtCcTP8FM0A9WenFGemgyhGXPuMbPlHCi
izWJVbetpoY28RgsWvVqWrvaVoQz55jZdHCx62JuysJDRjkYvUOzjrc/FHU5
NHCiCbiNuLpbYofUuI+sixP1z9neBbZgGXQO/dJZBb/qDV3d/nuvQi7xtZYC
zC0/NERcjE0yTKpMNGtgl/pGTUkSPRvB70WWKLjur9FUKzrg8iIaolkT1rKD
Er4ja4NAzfAVln6j98/NEnAPzW4/vl9NQuYnEARHrb5QDWJ+rrtE7ZyG5G0M
NL7a5NjF8jy3HSYrmwX6wx93jijV6e1gN9LtoA0ppPUdZsBHpsD1CytK6aAq
X5643gDUgsU4R6CBK9r9mTNmiEbdPpz2ITMO0tXzMlpWUVQHTh+ijghVLAdV
s+AvWJaBPdUnvIpnBokx8rbC/HT0S6dsKR9lSTfEJ772tDQ5Vx3vu1+UhHPC
4NTke6aCxA1kVEvTfS0n9ojqGMo4cOjynHDXsok29r+i0ubuyRPPWNiSUPEC
BQe3OWRQ6F9RHyvD73IcKNFQtDuOFgEdeHmqUT4hcEQlCW45lb4phli5dlx2
7hh8ZSN183IGZbvIKx6BJU5lPAHcNRFwIGtHKHh6RaixC9VxQVYpv0d7HIVD
cOyUY6hQKKrAutzuUIg9KRIgpV0gOa23OBIw8fejCWad+KrQthsIIM+Q7WQP
Ysp7qUVnypUKCXb6px2njSyJ1S0s02VOB7Haqkwy09DF5w/xgjWg+xSafuFc
OVpyZX/xFJmcBd9hKPF36Vom1P3+71AJzomSzKpZaNAgTilKo+KvKa5QgQgD
jB310A64+JEFBPCiWXobee3LiOedicbviUcVJJ7RLzWYLlnfTEdEA655QDDc
lVsiD42JNFYVdK0+y16ikhm/NeX9jzyF27S78qp5mMwDVYaiUp23Ivnsw3Od
gyhD5emL/eq7/sDJxPBqBi/GhMAv9w3Y6wyWo8cNMf5xLDvT+rdHOyHzW+iW
kFCQDeCe3LTqLghBkABdpLQq/flpK94YGoMyVavLBF9dMctS+PFfBNFP55QK
Q0hhRQidAIXVRGFWPqYYPZD3yJo9WwwqWE7jOOLoRlZuuTAwc01K9XCdVBg5
hEHSYohbjmyEb8OWIlE8jX389GhTASyGaRcr9kbFuSV17/sHzpZlANKmIbrX
LztgoFH6/8nXEjJXaS3znUBAZ5FS0OXEj6mNP5srgHaE7xgvxIQoOfoIeJS0
lZ6iF5Zaxze2AzuBfBRx7Ra3JaKHZjKOWYse2KL65+z7vCqriIbu704qi0Xp
IEc3RhtGe4T5ZHeI5oFXPKE4lznIeOA8Ye0zrNLmpg1EHRJTOQKM1TM4E5zM
IuKUG9Uk/uE38BtdaXgvgz8pDZR2nRxJJqyBSx9kwIa44VfbOojAwulA/kJx
5rgUqX3tzCV0oARMNd7TuxqNWP32qLs/BGZW+M6gL7zcFB6HWDOZpIpCaXbL
zRBCoGuypEyIXgdJRuW2tGdzeY0VNs1pApia88d3R0c2k9U5YqJrqV4WVuLT
BW/ffVeHeNYLT4g2hfIACbPtvCs9IfNm+mkMC/pMijzxMo2Ct93xQXMBC+95
NNykjLg/wd4KkehZFonDyLLoHuRUJlgIAeIjaB+KTKi2Hcl+Iv6fQWrcL7iB
LJ0eHnGNPKOcPVhSGklf8oOPiob50ydwcx9wLAj+Fkh5msLEqzjV5JYRCvyb
TBmcJGedeWlp6zQjPPiaNoxx4cA+G0uuPCWhRTSDHE5MUlppSCMJaxG4nBPC
XQ1IBTVbkkeDnTvsMtE3OWRfmKKpAWmnsCey2KQTszcxenLPkxGg+KhC1Her
2kcC368n3tQc3sPjobdBBvLuRi/MZtOEs0QSbIX5An2p4Vr+185TlJwj3HNr
5sZcrV8xhzuRddyQVKG8lfXIx/dDwMxSew7CksVk4lVZ7TCurSH/Rl7hfhS7
IzW0h7MNc6zvVXViXKGFqPqEd+dLu3p2VrHebg22grCcD84OIarpiit700Rh
D29n4pRybjfj00xWghfMSEqNnuvQ8YC4gOVVeXRFhbAAdKmLlCDi68s7Ptgo
Vx1cBmKCORh9C9cea+JOmjwjD0kPS3/rl/ESXprbFA+ykjqJTdzFwVaISt7R
YjTGGPds2x0jNOtMPZw95s+J17Y5NEtoTOw+nGmu1EoxnBuShiy5zCsK1v1B
RzJHzfblHBVQrT7jzGen0THlrEUDEWntXl8MiVKFu+tomm659HtgairYKZcW
Bb+NQfLe6VwCzcQNArIDMpa9qaPC6ZKRzkSn2mjNJUCQ9+9/RsAkzB6fy/ff
ANb8PlE83rsHVBkSgcb5qgWwJAEb3TMk2Btguhi6Md8NkrZDkLPyz+BwHDTV
E4/JyVmW2mRh6aSKpXiocbRLs3hy647Ea5RMbLBiSmmKNNjiSIoFISB3PC1G
l5YYCuPnKKIWsX1XVYR8CZk+M1C+nkafEC/n0qRx6EYxrLuvsACemsHB0vhO
/tF6J3LaAaFbkMplzZlZmwX6W0S7CAcZDBUxLrPq3zEO83oWBNZFsOy0GbwL
CjHmEKK+TywY183EaFSiZqh7Cn2tU9SKfF3T3IKseuy16qt2dyi7hoc/xmnR
qeE8LeGtdoQtwJM9A7TeeAKBg/m1j9YF3kgPE70FZFbIWGqhiSj8nmK3sXJc
BxJSVMkbRrQzVSqo/xTN8gPg7fl1jXnN2R5w6aGXqlDEmYI2AcR2fBFLTcNp
VcvSesOhnn0mgx6cIPZGbAIBdj+InULQ6MH+4ELD0LsUaA9tCJ1rRq6YEWDS
5GZgqFgU4wpfkd/AOXHqNU54nuvrMrXGS3lFlQxAITYFP6mPvGAqmdX7APjd
skcPioAvfTgFjXdLvspfvNr7PilBi9pH3BMAF+6hqEmKji+X3lrhWLXSsRoZ
xet2Rv22q4ef1JWHSS2i6iBUrUSedq6JIfY5jDQ1Niw7eJqZdodyTq+fZDK1
O96prxiVXXrSWQuh87WRqxilzvgKQMAFOQB7GD+S1IaKrXx2SmfUliWzhW20
C0Upeqn5TEfzeiwduTvoeZb9MbITqSy9xYiMXOdiGX2dA+Zk0qODQRdPWoO+
cxxCYQg71jUKQVBeiOcLmdYYeZJJ/owJiTJkz3l/U3ekzPLZ+smYx+/jcdbo
iYM27nLYTMPMBGGxcuCKGbnkBbSMdypEAnEOSNaJe0pIYXLqx2Ei7Xgq2BE9
vu1+bnOIcLO+p4I10P1ynq1lmNPrh0r+5dyUoY+h3HO/hMm7sq7Aro9nJvRT
7WoMtoKL+6KGcsUpJtlLlW6M98G/coi4gsdXLV3vn7/o9nOGzfgoRtzl31Jx
KYXJXtGTfxYpxJGNlW86U9437jxvisbj7xGQOi8X2FTOCmQJxJY9cWJG1D/A
4bKadh3X8loB4ZaOIBSSA5ZOKJEkSgIe9Cz7qyLURwRx6cx2Z1da+XLIYxtN
LFkzFNDde3yxb8PfJ7Io6t+MlMmt5rxOB/KWwtx7zLiq51NUs9mIUYulGaPv
Sby5gvD+7W4JVrvtctO5PBp7m38Eivk8csoU4hvdMvLPzPZhW9dC0Bpwzgh0
f+OLMiBN9VTScbOCEK/HXMxXJ53nYDtvAr2fKFWv/cWFJzmiLaZT4nBjlPA0
RzI66yNDjbLYOXBaNrQj8Iz+PYZQhtPGmd6B1WJWxPGe1yYGGYsTDCLoS9gc
eFl0xqUeSEqWgqrb7nsuRvudoT+pzgy5tV7UQbWrVI/lV6+c87Tn6fy0vHOO
Bn6AsjRPgH5dnXTjIx73WuCIc2tbsJEPt3iCc86mGeZVndgwRPrSgIVgRzL1
8eyrUo/ANbvfwg8wfS7td55/iWV1E+j/AEKvs3GdjEaKtATVYuJU+X9h1NcO
SHGh3mezB0jU7VZRu1+mB+GkxUwrFOh+6CqyyY1L9gLPvOlucrVUEzZSwtXw
Gdao7bGkoLl5tP2i8BPlTlQDqp37mZEgfnUyHy2EpansML9HcuWcvTJqqWQj
uk7SudBPCaVKnTUos7C3z3PgK/kxOVXHUazPoTkpL8EifZRqmYFjIjiH6YI4
7kiDU5g+x/vhTbdChyZ2oMesnRxxkCGVRWioMc0TIlh5opK7bktNDV38AxKI
tZDvpf7oPhmX6RtcaywL2rSgPlnuBUhqtrQE9jxmXl4xgX2FhuoTQIPcPj3V
qeLgq6IqJnLd2X/ZQXIz+GBu+Ib1glhTognDKp8qhicFdVwhijbCCV4j5+Z9
UaqlOtusWQfzqI6GGj8M3AiBWRxfZgJ82VhqmIYfLLuKpLZo2hZQNXwMkC8R
pbkmvPdE86OVmKYnMfRkES0YJ4b6LrBhiPmQwFAbZpA4/aXxAF9d84iZv6sY
682jXdqTvQMxfBCnKdOQJTqPAJItsLUszI/va+69o4gSiUNH5tynesJsZBjH
VEOTzPhC7yRUiQtNpW0onnx6ApGO7mL7jqh6fXwVfEFKSiotLm5kfK3hQ4Cd
a6LFrBO20cVwHE5bGUBFxIDkM5nUa1QTHXD6+uBHcPSNOLVNQEhtB/oOi3hJ
bTGQb+oHEfRGMkhWaBFUPnDZY1yswhbK+XUaLdxBsJi3Yb/AYfPbIdSax7g8
1kDHY0LE4GE6+V9J8RRVTFDprrbbmKY9cLHPiCTA9vhQU4jc4I8uryr1PuGB
ygaG48MV6zKtUSiy7oBbcWVFUf97ijtg1s9P1114GHgP03WnZMbFoTJQGhzS
AxcXZyvBpeClGOXyx/9PHQfTQgsMBgaDJQMzrLU/4LaJoGT2jZ6hUjVuhxi3
uodijuneAUUBZSBWjJhKi++qtXSj+yTQPQFIghOUe/jlDXH/Raol+E+AuPYN
SzbrHR/E0TkspkFLdmn2z/M2rRkt0vPokyBeZfyyxh0jJph3o7GbygZU4lz/
89DAzFo9KT+TSDqSRwjKMQiTYh/m3h6BGtxvUuPTcLZuxGrGyteTjDPut7a6
tok9zE1efrKzBpCakUlOfUvBTEWhVkVJlW6h0eDqqC/Oo/z0C2oLQEiPGevF
Wayc8DiT9xdR+g7XrEIQEqp8cLlvgVvmNHG6qzTEXsfoY//lIZxWh9XQaURA
GHANJjYIwtiemEK9THuZb2xfYY6CZz+sLty64oZFBpIbm3t3h2gBCWz/VmU9
jEeiJHQC01Ti+NpNjCbmKnziUgEnuwosp4Y+NIV+DilRtgkd4yRm7Z45a0pu
m158mCQ4cP5qAlbprOxOZfjbrzz0xnFtS/KVbMtTdTxjxZaUzMszxCX2yKGP
lFeN1zb46+xMrg3Q3GD7+vJ35daPsuMO2swA4LdS8l1+nOnRDuTUKSZmoroW
b2uQeLjxe7iU+oyg4YQUX4RgkTzgsi5RaCtRyYIlYo9m/YIkzmdaa2ACqhLA
8hvr3Uprp1+PLrHQoIsAdAAW8flO/rXNftBIFUZLnd6xrWSZONUOWndeafvG
G2r7nQ7dkpsDdKaIxIV0PEvZx+yNl+WRXPlnPjgAUowF7VxYdy3LsseXNpl/
RyZ/OGoZBQbCSzYYkpy1KylG7Ik2FNJ6ws4g0XjLzZV+CyggXA3c7xyN9jeC
eQd8cTyWKQw4b2CpDuIX3w1wlp/moQ45KdFVHS3bG4UBQOQeT5wAAHzgERfW
xfG/5jcxSPixp3xlAXLyWfX9ZvtNr1Nd/0LF1y7jjvc5zJAMezalGADRIgiR
oo0c1x7ekml2HWt4SClG77RbCCcukX3pIEDJToYNhHntdjwMLJ4IaW4/AFl4
buj6XE/54OIYYRscErcKLtzVIR7sTDfD4zw9SotHGWEaq49rKNW1kU2qViAD
4k1H2G6ZIQSfhAd3L99P2oPJ8w+9+nwmSiHGAx0WjDyw1wiIXYHdoIsOnCy6
j7yZhqoJOKnnGcGvOwzbRYKGoYyFXo/NbNoiWOmQDwAvj/sA5MGgDU7QOJ3p
VQbLKvbo23nGIocl1Ebz4SIfHVtYKBE2QZGhnKVyD8yP7aT8INyuM37KiCYv
Vb4YScgr3J1S+5IEgsEvQsEDPdFwL+sgi2pvg8NkjGszFs1k/RJlufGAnqMW
VMiLv0YrdKU8xxkjBljP6lEW7D2mxinUZD91GU6s0uMfHGtIl6U0jjJ/Lq58
ILa0X9XSEVH4MqMXh557/yOYrmUVUWKtfYl2qfqoSQzdDRkz6RXmb5uADmHC
UvLcE4ydE3fJjAv2pzXeqNya0tcw7rjdD1yGhJHmnmWm3dTAoax+pCQW5YbO
sNNxAdA+piohWcsz9Rpeami3RxMTkK0dD5iUSpeFW/hRaXtRv4xfK158HHmZ
T6ifz2KKJ2y1KAjodVVX/a4WsEwk+K4dxz+FJc1TGN1JWhypyTGn+QPk/Cbr
CnaFfnB8h4FuZDepVSdvf8ejRe9TBCi0BMveJMGfw+QNYiKGQvjgW+FVRw40
2B0Sss2U87NCqNqqftClztnZt3H4GIdUEF2/YUbHajLOJOGFgqar3sKyQmSH
ng5EGmiKRX8BoqXvs6SDLYBf+AQLmE5iSaE2cjA4A76vYwEaVWMsq5lOUwdY
tsbCzWgRlyM1rcNA/BQu+srsYsFytgK9jNISZfUqvcDcXGfDeK8wvoXbS7Ql
CDBOmjVoB3HHt0/3ApWJ8Uk+jO69/3VBp2fee+GdE1/3w89bxTE+VwCH4ukG
DM1Di1/OKAC24y0RwVoU+xQ98fVji5MoV+HPl2iSVAEeRQMTsEu2PzxEIcTE
ufoXImWNxh8H3ne5KaOy+c55T1/77yEDK0fRhSxhQkqHJQg9yoKUtUxfkDBr
wso7Kr577+rgKFxERWrRxep3m0dsJ0WEbd71u6fNChrbJ+njSd4vdXTPv2bM
BKGROf9WbP1Ueksc0X6abdQrUQSX+Zg615YSUaE1/LcXHo68Mv9axG2SUsSq
SiZKbSik663+V+sxU91epR9e/rjAc98wHi+qR/6JPT4v+7bXVYmrHlXkA4qF
kV0XXKreDvDBz0E79k0pK1Fw2M02+GnslnOjqlYe0aFTWA06B9+7msfkGxk4
igx7Tq46LAC/eDteN8VrtdjVGMnlm9lMQy7o7k73b5c2mY0fDKVCc/0tVPTG
6RkIbZf6cUJm3tGd8xTSF0OVzivaQYU4bM4ZGHzF2Ef0CrDwUH5UJFLlFpfr
xAXpNhMMNhxBYV2lNTovmVpn2KEpyHli/nvq3BlQ22uEjBf2DCzK6CZLdTF6
RjV8VhTXU6MSp+BTcYazj/DHcR2y3SqXdP+Izb5Gp56SCpXTvHwCD/oGWal9
zYgMzCm2mpu3HsW+DnHM8gpUPPWt0HrRXJwPdlLbeZAJoO8gaHtYvvUaW9fK
np1Eomzov81Y094HTO7SUh3pWczoOh5XB5L2UBich2LoXK25coyHdR3KXiOt
GFc5y3UDAxmbXuYnGH0kygJPOVhc5dWpNRr97d4sIf25DbCGkWmRt4b8hucU
fpwYVK94oglPMiGCah6e+JommfNOXozP31oNN2gBPwOFQjW3eeWGfwdnEEho
1+RPlZlPBenNhhoXO+iChWmv335Gq3a8EVcRrtHS3SNATXVlPe/T9XqveYL1
1gTfxDHw+7WNrBMja4vvaV4WQwbNzp8NpnXgUBsPdKo6k7z781YvavRb5mNz
hulVjwUqp+1ANSWI6GDvF5T6qZhplQ2wS+wkSJJDN4OURKIIrpENX8RuXd35
7praPkSBW+rwx2wOC4S7MTrez54Ekz861ZrmMBS3NOZhgW2jU8pKMYXnzO6X
gj1Y+zZIgHOVUggokn4dnWnGVB9CRibo/v1/mCbg/HQvxDr3zfwZzknKlE8R
2w0AiwLB/SAS81JOPkdNFEQN8cyxMgKgTZrkN9JojUGge7EePMcLiWfbh6JO
benRnCuoVgxAeIvgYt3wGPddgFiVdfs4hvY0ZlKVHxmIgcoRnzYHTi2ulTx4
Gw+KZCa1/J0+5sia4yEDN7k7Py6Ikl8rq0wMJ/1FwRIIgmKRCOmrb7Y/GqRg
qC7zWQcdvrVooQSPvw6gqbtJKPvirA9ZvVKuYESLtjpOvDJzamxsfQttjov1
R11RrVInrmTuRLtXnRv7fHyd0x5pX/nly60kUPGPrOoI+2c97e1uALJnzHy3
I4sE8nwVMD7hV1mj8Rwf0z6X6swjegk8siRksdpm/vsSUqj9IgXGQYKXDfaD
rtlaqMj5SMqtxd6xTD9buD+oZ8p5ek+G3LiHrT69cgVFBYPbK85pwOhJVlPw
XgoL5GISylUoczX1F2Z5BWQQAPgSY0wSkzF8R+JbgAnl7nYFUFzu1d3Zrbny
fv+PdjdCeo1hyTn7gJqxqc8gviEhaY7nESxz1UsJ+7WOpdombunJNRsC30jI
krB5LHFVjrcET92UprUQNF7PU6M57QUyPYpjIpJhePaWP3QS71JP3pBtccWX
FKwVc89sKw8dLkukZgvvarJauhw5r2VKjnarMmDZVBX02SYZQRbPVk05v4DB
7KZ0rJwng9TOIqEII8LKFjSe0SadByTEywsktC7tFtbiq2UZIT5JlNpkaDUp
1YiC5k1USQ9yTR9sxpBTNfg585ccyyfxDDb0CDgY0HLX/w2aFVbzEOGMi9ge
Y+fSD3o70xF57xtp7bQ9j2xh5KBX1nJHHStd0B+T8jNePYGHqxlBomYmrmML
kJ1b7arCewAAFE3jgJQG8EdIpEt9uJf+JWX3jTfCPtlpxWcJEvQ49cx77AiX
FsUsWzUQAbR5Aa2a/PapTcg6V7gMLLKcwOqH+MVaNgfYkODHDGuTAmsEUW5m
fYJCSSBSV1kj3u2r3hGygspAwIn2PQH/Y9BrhXErugVs6rIU4t1XGS3ABlLm
zIcZsIV9QP0RaPcMfKgYqdpXYAMtlqNfMaAkEsxlRL6p/9qP+LRm1WO3bOgZ
79A9AeDlyU3KUxLHCuAoLgd6CGOYqWhPVy76Wc92/7UGbVTcx4ek5T3GJLE0
sjlcD8YqQKouVuirRq0QH8lIJsbhiWAMh3aU1fnQmDaSWBJrraWym/2gBQao
UwQOfDu/noHGnrWeL9ii2ps0gUkRzr/7iuCRh6bRdhSLX/muc9eOIzJSpd9S
wUm7aoaCXEifql2SDGSr3ELdL+XiKb3fhor+MBYxD3OQNv1tSW+JZx2iCVAq
diXE6JQk6M3jL/mev7pPMwCfs65LzTcAbRhsBrtzqVwJZDwdl3m1EwBWVd/z
v7OsyWx+ZPDazFoC64Zn8i4ZvbH9aQ5OKVBcsx7buFNvri2N39zKdIfBZL7h
AuhDpwfwp3nI+RPfGASb3opkRpZfXMtuYVxAXcCeQKiY5coSFw1HkX2Tj4NV
iuOYlBfAmSU9b3CYl5YZTkybUeXvOjRDxINFqwEquxPtDLFiEfg22R0krv72
/1xQpFE4/JhWhJbcQk1bfG0F/ynGkx07PgGI9ZqVmLlIazlIexPkdJJdmRqR
Lo3S9DJEkEXNDuHPslm8OiRM048JU1n7BHSmSnsXRn6q7B9ySctl5GMf5OnB
f/+ujF/mNhU2TD7D2qhqAdeoiSrD7Ybwp3wICum+iuQMN0h9HXNe/jMYvs1k
chEYk1yok0MucJbBlcKf+0+IQSgWmRIv+84X4xTBqWSdENV+BgQf9RsfbQuN
Vrzor2nGb2uW/8BXvAeTk8TF7NyUUOtQibOP0qSWp4drIUQw+UTXbK3GqjUJ
76l3RSLCt86zJsk2pArsA7Pocx8oep7bn2efqCfY/wkwkCaVa9Ln5gEVtDM2
HQ8XsYW3+KiXzoOdXCQRosV3++ETVa1HlwcL4IXr0WUPFc6qlZuBTsqxPdhA
/OJAenIbtT3JwOWYisjMrj8CwWRY/l8snzk8cjZSvaTDEIpFIXSQPx3/7sJT
LQ26kq/Sq+R/wZ6hPGUFKbS519XJ6E9SRVhq66n+7q6IaZQxJAhEm0TLYY9e
0qMYr33SllKDTAWHe+BIqqNZvpyocRxGhNqNHSrpsUL2PB3xwf6YMW25Ksb7
isCByLzj2HZmOUEwRyaXZrjpCvIOxpTeTTlh3n6wNLxqdfRtAJ/mYLwkEPyZ
Fwn4g0JmqRCKs05jqRXiEx5OzgE613KJyJ9ZcLLh36FypD3vMHuy50s9+WBU
LDNa/4brd6QHSJYlmvHmIO9//XkUufgpLA3J0aBgldoAykU17Wbp8+TNLq5A
kgnWjWeSWICI4nzd55zSQ70CTM2e73nShy6Sz+kjy0A/dG3I+k8gZAB+aFX7
hBPol0FyODRG1A6lppw4rnFDOVmIsbGI+F2IhbARp7xirI+FJw+nPQ6PtjhM
JTjdlPXYtFN5GDLc0gcxl3FSxCPM7UrXuYnj26SVY/gvAtdQPE+2hH6wrUux
+3cGYt/ME/d/bbH4EmYnvK56ZQfaLNcSTTGOgMhKE/m6AJ0+2vGCvolKH3eM
Qt1tLGio2h1GUV6HQ7welXiyY9w=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AHFS8uhOzEEv0qANUjCa5shxFe8bemKFNhQTqRGtC4pjovR6jkEwCgEM+HVx2+RETJ81jdGctIsI8rtsCu4TOBbfINYgMfPtAhYoq0pIwXzpBYW/Jwh89yYqmQ/8qwf+UZ/RCUPZ9uTW2DZjLM/8DQwcPSaWPn4uluTziVOYaXqZBjqnFFKudtGOgi9fUYcdgmgi1Cr8qg3AFyDXZaw0JPfMHv+sI1tXM9FJgZxRxGPfe4leCTFNMvsYW25Qct/kz1eFletWh2Ydd4OncEWeNwv1g90DI3nMh4hlnCk3GqyxT9z1PMHciyGxAjGVOmrmYNKQrb7p8X0q1Xm4MtWPFyG2BDtkGL0wtVE91oFu4thsQ/+Prv9xt/NJNIEUdhe+egyChRvVywp9CDJ18cvrHqoE6pVgVqqZOM5JIVpJ30Y6rWp156eY69CTNgyBMSdtf3UgN6igY3sd89XdlmEuNmrt65rJU2wEnH8rxw807hJBELzCMsDKIjnI1dRQExFm91Rggx9Iu+HY6TPT7AIdaguAtDXJ8vZ3390GKKooSi9zaKxLcAu0nJV6KB45VJ6vMJhZSuSGqefQcawi0tFBK+/3cYK6QjQ+GpuLi/YfAV2lEnSIVe5lpLOY6XED4lLFQwce/hf4uyq6fdc3QaecyaWHNFJXD1QfvEpGWGRP1PJneXMfaB+enzN323UvfMs84/8q3+5p+xjt+S0YRwYpTFNK1QomW+oolCahesKbJrIwcUr4uYTChX0b0eOrS5qBXrklYtw8DA6fAT8mqFwHVlLPlP/NBLX0ggsEOdWqd9vV6EaM1QIXJHvfz9mVeudamYGsu4XguYwkKfJLDdsIUkeT9QN/BXbQ9jjHNg3O92qDDEr06NXmAGU/zxickafAlu36QBEndQomamIdI5SU/EPyVNdKIzlUS8vSmWlXwz3/iqYpPnwesS2lTRWUPclWf3qvCghauuATAmo5RvNY68CQAk1Mg+Up/A7faVEPtHTR2aLPLvpzZp/z62HVHIjN"
`endif