// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rbksR59+SyDozUHiGZu6WwtLpngYi0RfNN0880VeJqK5h7sAxd4jDh/86ucv
H6LBRLdXxVtFlow4maWhdDuUtx66a7krV8RhsC3AbGWupxfc3JXJDWS7n74x
tuSD9Sylh4fGDValV8eZEfvuZYucDMIIZp8/6+DvzJCQINxWq2nfD+mJYQGS
65Uw3PdS+WHKHymyCQEprDUWXvLKlp2ngLGHiO3i7PTvTXiKFrb3KD+/CR90
gNyMC5/TJZtexQqhfknnVdimNg3ZD60yh707NZVT8v1g79z7qycIcVlr0kxf
J8OIG0ngsfun7nQhDFDAnquWMhHbWKRvbhyVVgi2ZA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GKPN0RGhsmGVCi6HgakL99fBtjBCNRbiMVmO3SSrqyOZmtHpC6JBUxFkmiCu
wlwwzVnfiLutKBA6Mi4ey14Z6mRUr/Pl06PjHa2l4wraBPBQB5MIe71WlT69
ZJG925MGpYqxSJQDbik3+3RJsw1tqoLR8G+dslM8fTeDVpaLDzpHRXC5v0ZE
rF7hRptBr1rVYuCw48hhCDnqRDgvHz8f2Dw9dsvGLie9mMKeDWNa80fYWtZS
M30lwZQ4cDvKuTnORI5/fsQbJH4SzCH/PqQvb7OHmWhZUtS4rY49Ex2DItGq
BuSduhBwRsPT8I6XyAmBgNm6J7w6vdpkY7kYiPoguA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
uH/0mXkDB54GpfpwQ78rnvzRJqzj5X6p64lLgMJdRVTlV/gGe585SFimj5lN
YuExeTvdRebB9cwYGiC/pZ7jA4b362PmsaNF/4H901h+r/Xd8d5J2T886iVg
MTExX9w+9xaDjCzOllVzPuybuE7qORrqg+6DLsTIaki3yTSQ2G7IQPFTJWEa
yD4OVIPbA8/PdS12dG/eYGlZcn23rOqiJJseqtdee6hacnpohAxr+0XJmYNL
AbhOX+xGaDdea1FIlA/rct90AZWMM/eQvKKwppgrAEcGM6nYi6yuMzM2BVCh
0QbaC7l8o8VkHdPH+uM/Iyv2YkX9g5LBTu8N3iuaIg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DROrmZQSUhP3elS7ehc1mF/EzRrD85wxp2til0tzM0frF/KapxCSYnRyvVjZ
GyXH28o4agEYqdt6IOJ/uu2Etw5lj8m1Np5GQWwzwPjsnVzPqF0A3H/Wm+SH
woRSfrg9Go8KsbWuHKZWA1qNG/DRVndSRY0gD8Q+DUZ8ikCIksB8yTgFktMv
CFKCEnOCpmuud8UkE0u1KmE4CT9o4qJpHX9PpeLwtwpnIW9VmYGRY3qrx4pU
TYqPKlG1GfEIXjhcZ0B/5YzSfLsJc4hGYYA2A3cMj/wwSlzA4av0bZIcbFSt
an+4zOv6PQb3jkfyGnaCjaebRTerkQIhnpjLHO44RA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UVP8Ua6KRwTrzCHhqxaJqzgtvjU6QXwiqbwiuGPJt4T9NNdu5AkbXe+HRo/E
0TuYzjhFRvZ+t4D5Ynho1cQhwJlS52U578uZ18Dwt2bZdoYoLfJGoDbDquyI
E28heqAVSFSPWVD5Ui13a1mzz8Y+vSNCA+NWczibLQJjf3Vp9Dc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Q8oHELXjzjRbRQQqdFfcU65v8AhSgwk0OD/GGhvbccnw+oKwY1gZZ/lz1Bjo
SD5cjQkvR41A7U4M9Q3GAcgSNwKi1bQCBqvVSScHOqsaFrGxNyDHK5deZEbd
rozt2lcQ1Y/DOL3DyJvi2ua1zZr8a+ZaflTLOjOkOcIvvyJdY1MTRgSWFHQU
pA4lD+6WFw9Dhfk7WxvD4C6YbGV3ibVWArqlRNsK7O42IrpZl9fMEHU+FrB1
xZx2aKFTK89tOax1/kTGDUjGHWzHjIY8Gjo5xCstgpNvwsNappc+l3jH3d+m
Pau5otbAUY62xBwPLdmPTm94MHKiKFCY/82nYI7GpI0iliwXJsfQMPyjC4WC
z0+Nm/nhMaocg2W4M9amLiPF1FWX1Q7SmkeYnPGkH1iOdPPTkLEjYwjfHqgn
ij7qpjEeO6l+7juo2IPLWCwESrl22Onib7l5zjLFsEDlPTEwVqjppu1fDxe1
vFxdjU/YTBe0lzE/3iOSgcLz4FvRPhAH


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HB++uC/eeUJ62GvFpsUBZGLdGXwjQxrsoGviKRNE2OzPCmhzdRlbIDhCisT6
sNtZlovpQfUrBPmw5+uKB5ldjZGG1M96q61fxuS8SacF4begbnXPHHVpcAnN
UhHA43DjwXbqq2aeog6ZhZmVdy9oOB+uQwCoQDC9ZVybk+Xj9Bw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
COSz9Giwgc9gxH40s3Skqvmmr8tLoT9g1ZVYBuea5rnXCBeyOQi9HhWGUSVw
3psmb1Xr1P9Pg76ZcgBtoE1YaFDFftCM04vj02aUX/ILGpN/YmpBwaoMlxvt
V5V2v8ATrYgl/5vPwgpshWfsKQ4TttRu+XBamCM0urjRyoJ3ff0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9664)
`pragma protect data_block
rx1qtkXl1M0PpFEIiVLc1YOvteiMK/Z2tRTBjhq36u0+PnUtmxuMRTjc3vMB
el0rwJTm+6N18iOANJbuvqJQhPV3qVm0zIoqzPpFlz20ezpmw2IofFnAG3pR
3NwQPyQn/qsq4QnrZmffMjB71n7nDLydwthjYFGLnQy/Vw7j7BvaNwvIRXpp
gEMdWi0joZVCw6FvYSBQQ5R19/bfqseMR6cE9WJCZO9aDIsUl0RcTNvKSNQN
PLDVHjLcDz9P95uQvfY4UsGUT2Oav7h49qNRA4SdP03/kSJ7+IwWBPgkA5Ry
pSEIjRSx2fOnxHBwIETvyVjQBBvtgD2BZ9zldFoqGYO96uQ9qAtQQj0aO1jY
gJWU/LwtVhUP45f6aCJQ4XkCWdzhLden3Yh0o80AQLM1LKaNKGyn9zP2JKhh
VpjyTg8g7PQqjtH+blI++gaKTa5xxIjjrTen8+eOjGHCEOgIpSZFgyP9wy6x
9WDQVpc16PEWnjYI9jUjuIqggAPTwYPWN/u0RvXlIGWEAiMiP4NGWS3wGPOM
PtdWRtGvziOeCS5rYjuUMDIr3O+7mJS0nDW33uc9jKalUl4Y9o0JxkkWG4kt
T04MxZ1sBFf7oLCCF8Y8Uu4UQrB+zb8rM5yfr1r+5RTkbhLxe7gRzB2W6oFR
/AhbNnrRaoniJSK+WAhv+8jlJXN5AxMGPr6QFOpQg5JibfzbPGRHhCI3ZShs
0uNDAWyVBSLdRknQDj4cSqNLaTiqD4s77XRtgDZ5s9TWPQG2hRgAwTaQ5bgY
eRfuv6N4TE1f4Srb+URX71AxzOMeLIKxivQj5oWDsHh5QfgKbIgt8oqZsriO
5NbuRIcYuP2NpSlnDOLN631+uI4rlYz1ZuVK3H192tdIW+rspmEbdqhEcuc7
15d1ducWLjI6byy5hSsYRs/abQCl57Egqxlzy8xdsj7ZXhbndk5/rQaWXAoZ
J4REvwoJ1k+Eo9GVQD6E6elIBJayNZ/+wdRv5zlZzbTtutVXFMkbKvitEJM9
0tTf2kq2iNYqJbcCaUpXEmUynQU4We8ENi2ZwJ3dVjEs0atdS0rDqyEQxjQf
yURWn/iBzpLpECNS99j7WDBTEzaPPnZdFN8cuaNypXMwT3I2WIVu6FpYtXB5
TzV2HVd+w6ANShpVDWuG49nmo4J/IGxyHHPvJGWlTuKCfuggu+bJ/gMxdVlw
d9B/4FnJX08V1FMGS/gwWTm2vzUv+WxeLEUeNTnPn3D/Mb+zSnddDmLVkAJq
zXLf9fwNJtwUudixMq3eeBLADN/VAmmqsxhY2M1Wq1HMje82Zuudiem2GeTk
LFkSekrIyG5gwyNPH13Ka0DJfErDdLZgtjACGA2poc7a3hVsEe5z8+XryjJ4
66cL0wqOVPF/Kl6ipZFzkkebvHi4ITNjoBgWZRK3sqUSbwKSKM09sgkOahF1
Kvub5OdUfrCZ2NNDbLVTSAwXOtImr7p567Xat+5j2Xb05Ss12xesGQXQzcU5
2ymSATRbTH25Hg5vOXXHg9dajMxv0FfpBwPFRJtpPFQfIBZVMvhx0Sz7nvQB
swhMskuFY0ptfelxwQjwqLAF6uyVt/siWdjLGbbiBox+ZSzJ994gOPrsH9RM
ieJ2EUGC4Y9XzuNgGtd587sNe76xQUAUGZRBIFM+2qTTuJmOHRqcnmEM2KPK
fx4+BSuClAqzMVKQJ3+ugnw5hadCgzIEL+agjub77p8y78J/w87RQ679kYGQ
Vk3XtgZispEAPVWHHQ4iiPWTzDKoyVq0uI+P5fiX72yH9+N6V3zPhkN+Glbe
o/XCbh0SuqHj7PSY6j+KLWJ2LXGR9lK3lZIdAC/l7plpj4S/Yl55WuOxWTEe
g4UGy45DTGO1BCt5Go9PAhjdnBQVF+zvpbgpBkyffHiJG0H2fp62WmPwRjt1
oTCEiWphFAqiBFd9dTfNrZdbVAJY+FHIl0NI+CkF5ocymT4pGGtZPUzbypaC
kxMGQ1JEH43vftEO+lLkCp6Y17h4dF53JH8k280IzRf/pGrUZOjTqwazreOW
WrKX9OvBVCQtNG9qQNic34T6e+egGeLfE4ZxpgJMxZfEok2XctSGhOrSYxXU
V7ISPlgt0s0tVJGX3+T0ai4A2TaJB2y+rbrWw5nIFhF+ohw5y+2l0vjgRS/l
uIPHqZEI8oWLbO2Oq/1hl/doTFedDYwA4Q078FGQG7/6le1Yk5EcUmxe0wsm
Q6URJQoCXJmU4JXeYLyUIZ0hYJkeB7aW2P1Xd0rTNYb+UGDp/ouYn2ZIWefQ
rDgFJ8MHuf74XroBV7LO9d58V9B9afSAJ+ke/W6mBJ5MSdDPomCHhDOmhzhS
I2LojGTHGyh7q5cuqjQr7vcqhFsIQiXWN4NP0EHLSL793Kl/UioWwchhMSdr
+7yKyKH9qCy5X7agskst838ZPOv8kb/IGg2tsu7ZL/RclAol2elpobm8uQvg
ZbFVaridDltBwno7Mxdn4QeVHqinh1a1UXlYr35tfPA30s1//9Vbn4+EXkd6
b6unp4gPSD9AEVXUvdA7lDNsYz7i6ow99E3RmiXZCh59I81HXBZySpWUkygg
sFpT+xkqaJ+VIFWkW7U9B9eHFdVw/M0dQKy9OfD5XrGB3fyqY/iyI0APhaKC
N/Vodpr1rJHUZB20GGzebWeYyIlgFT4YbUapaIfZ0vYu0+Nmz2BI2OwXuA8t
gWCNJOMMwTFz72VfMJaKXohVmf40hjqewrRqmVCsAbSRHGvEGyyeNjJmVPT7
wpJMzZvKIIE9mfntgCDsYIsKAB4v0bvo4yhVa8YXgJSEn19HbyEF4maIWaV6
DgfYDT8RQAJbmCD/I0gzepW5f1wBkmeOUfQ6U/tQVVQ8oCL6P3PYjR5qaMrk
zBDE990NkQyRfDfFhovaAGz6h7502ifYVcyN4f+yQVUdZX9/K7oacXbL8ZCc
xSi92AyypK3SNZ6LsnTIyyaIDS7CN9Mx9rwHZayo7wfT37qlpHG6GFJAGFCH
sntyMStr19m3mh6B5JyB6JTHCc19c4+zsLJ133VRt5ioq317FSOvpNuMVARa
Tlz7tvdyTopfpf+KdESI8o/qL+x7hf8cWW9x0efiwGGGdmSTMfhiETaxE7Qh
UDnmwYE63KvWA/TZG3sm3I8siCYOsbxCvbomKiLROCqVLWvECAGaeXBCTim/
+PZRUAXm62j8/A9geAaD0bE5v5AbZmS4QgYkUVprmV8ENCig4K5UtR2rjTOq
A4CUY/rtoFne7m+uuZIUiWDbUsCcaBp+sjoBBSL8RpJbxGohwWv7oRD3Qjo+
JfQtAQIa3jht3101JkO1L29M6osKzXLK1SQ+zDjdVByQTfB0b0pwM89hgnXE
qBImzBiQExZ8o+pmRFIPrVgPiZbCH1Qt5GOqVsWQf6p4SkSo4WPq7pVdpKee
m+o5YWQHBkn/NoR+XmQK13agfo2RhdlsCv2zai7CKcW4n6Y7BA9cjkaFnhPb
H1Wr11JsljzsF0GUNY64QqJqkhQtJtylXrPPovsb7gyzyvquyYqrsp5AD2Y3
8Md0ynwjkTAFDJw2C9+7/vpk07lD1CaMs4PTCA/LCGTBnOVYB5g/boMnG38e
SgdjIUqRKnF3Q/xdITnYA+7XIuCxVZJfKu3plSWSHL4atqBZNPa0AN/0Xucm
t2AeNia4WDUYOyVUxnBuoVf6s7AKSdwjN33ktpTGh6VH6aZPpkIBmjq3vjcS
42i+Nshk15Oi6+pQ33t2Lt/nz7zSl9RUT+ZH9aZVrchbq+T/+YoKBhOHEioe
oPsldZ9BNPN2k3k07rPP6T1uTZYQ1eQakPHGwExtdGvKI43YWqm44aCvlxkF
99eTENsCb/ZgFAq6hSg/paW8L3ronl+VPlRQDrnIUVe0f+lr1W8Ij6DF01mW
M8ejm1WOjjYYQfaMYZxJZliwZMYf7wL1k9TKLMQt2s3nBc34tKe0U4xzBIhA
2ds56d9PJUIBTRag/midwm2gs9fKO72RlF2glASXyziAZrNVdvwIC2KCwd7+
XPWZIPHllbuYUd5li7cs46YrHvFhY+Wol9hrY5kgF1EB3pCG8AYXHplWWwRJ
BlgeYUKbDoUeCejEbn69SNkZaZyiy5vtbX4qMBkvdwk7JB1NVhdtIc7WhXWT
TPuNhdg0xcTndB1G8KueXA/IQ2D69iV4gHnIzQaR7VjGWRDVqtgMSj5VIyl3
ewbAle8oL5iBCfE/Rr86BzpoLdM3gCwX9pEn4lzwHH4dgHLYujz8nnUQA5Nv
QfNgQxA2ly4E6LE2ivb3TLHjSVTSS47ABD0SjS6TGwAxI9bdB/lvR+iAByGi
ZNjEld7T8DNVmaJYdIVsh760XKpVO1mW0qaHE2dvhrbYVboPfP+BeQRY35BI
F1nkSdPT4CprKlyx70nIuQvmwKCr2oe9rclY996d7BsdU+hVFHF8GSzK4Z5k
D/t/Skrqjcvh2Jh2oD1m76iinSfHlShmlroGKNg2LWBS4FwOFpJzWg89s1Ck
hfOvydJo0Y+O44MfKaAETBBonh/ftimIjunDvSOeeBL/h3p6d0segCRXZaG+
f3dOf/TrsoEy/4hpZJ5G9aEH3ZM0fFeqUJtS0+Ld9HZOkdKAz6PZfhdrqJt4
h+CalfLmRZT/sdNccOTH7ADiW3jx9WMKaUqPwqCvTioCday3XgmGjXFGR/py
CfMPFI1ZHOJEUoWdGu9+L3aw+xCArcLuINtWgdPFuj2AeNjmUD05LuaVJoDA
n0efVJfncKl8TzNLqhJ7yCzzIQbIwF6dd6zUS6KCEilJLK+TvDApFyFvrFqY
NOP3bYVp1lepSsAHQumohDLuVJJOumlQ2il4M+/BGbd1fpceYWwQW+zKyVO9
V008sFEugLNcuj+JfCI04ys3U75sd5Wf/bMkCiFujwVUb5d6Y8cv22ByOo3b
NFDtvv0mig3sXXT6lilAos3lo3BqDhP4KkLA+piMsqxdUDXSu4lyPklejdV7
gimZVcXrsu1hymvQEYsvt9UdahtcEzTLbQgy1tQ8KrNMPg9msvld/zB5mWgY
FN50lp12vVvZC5+uRJSGVFv8gonLG3P1iMM8LMNHsEpICFOmYy8zNV8EnHoq
rRJVlxgcDZ2A/8zdZ9wj27Vw561D6k+0BTx//XhAW/B1MfWXVvMnBJxe93KC
eVpggmKI4XxYpwG1rFMSx/DkQpsBmQB6iknobvWeLlPSHdLwe3nU/07UkyQn
uqdlbboJhzRxovksOU/jOubEwIKOoq+A+d2yiQvhMht92RAFLaDg9Y3naXQy
HH/FtR4+UmdUH7sfMHQyoS0nX900XUemUN2QPpU0zHlyPiwyaYiq98d9bQpK
jVaM4Rmcxi60TJHmPkn4OKjzFYYv8QBh+QUSRIuOq+XpZeLxSgqOqOEGkalQ
eGlWKAH9OIlqzWyQvKHxDdYSG/kBfAPYYtftcrGQswrVBGQzeZL4uKI5OFYe
kSuu3LQcbgkuS7PP3dbwtvZfjzESBcTJpvGuSkBcNGoTjfxzQIzuqpCmV2oc
5rKFnWXBAh1uIh+sfH19dhCKuH0QP31TwS93YekOwVz7S0NVi+MKtSTUvQYw
YKXwIvch8NSJ1R8Q8FqYLpvMyHRg6lfNdizd8oFk7f0lGfCJt4WO51Xcxola
BCjq0qzgO0XXMHAqtjRv0nOgVs2p/DwgiOcxJ/Td8U1DruvvUDYKyx955HJC
ZIQlahkg4uYStptkdcaKvQylAzHWtXrJLCVJPYC3xVKH9eLK7UZpMzp3yX7U
+rXn3n5Qy2zja+g398KqjZpE44Ct5UAzikaQeNPIWTcJFOTBpo231GntCan3
fkfkXb+soDj6xArFuBsmvHU7rJnjUjGnCednd5zT0Twl/gZLK9Z/9ac9sJER
4ngBPqgF8xWGaOIXVjEY54IACjJQXebX5uotkbq7JFkU5mQNsC8cGZua+Oeb
YHZ68JFpjXjwBgpq5/i1yYnATQwVDWc2SfVEE1KZ8Pl8pO4H40YpjnQsF26R
yxNkVHZ1XNSaU0VInLCFGtkrwecHB2GUPflRy3/kOPp0MZ+36A8akiaHVLO9
tafX7EsN0Yf4u02HlV6JIM71InX9B0hSMcJn2hmkMtOARRxRHuWkUAAyLdGb
4Tal65M7qPyUIG/Ajzmb+dGZjH5viJ0IfjTh+wdftD4D+9caZ1snHGJxYKQi
Qr5WwcwQv+05NvDOYy81thsUiKMvup+S4PFAFU5i6raXatRfEFKe5Ryh2iP+
6uir+CUVuwC5TzctvGVCbn9Us3m4knu0SrEx90d4itzpYdhQnNw2gXzlF1oi
hquhW6+v2KJ1T5Izun6QfQHD5wH08fE68iIVagNcT949G371g/YTmViNJfpq
o5qYBdfsxUdsFbTJPN0ufO5D6EiAax2jTlL0wsGDXUnKp42Zr8Fss193zI/B
/IIhW3v1cj0z2NZu/079/CQIBK0dRhcJMUdqU9dkbFy+7qIo/l6UOEhauNoX
8dhuq8JOkbWedUAVE5x5DRVj1kF8XRsZ7VanEPyzLiuh1B2XQoIz72wt7HmC
6DQORJ12ZkIJKF8FYrIFZ1znFAih1YCF7RpLmrlwaz4gbPxvNYqEEMmEjAm2
dS78771o/mcCe0XD5Zd4vo0LGiUgcjZvM3Jde5KIa+sQzHj82+6MxSEi8MyY
BOJpX2f5g7oxOMVcVHKsUBJZkXSQDP8Xvbs9d1dLhIvl0SY633tF8OttUEhi
yJuG+Q/QhxJYSrPJTpGCtwqLQDwqeulShtEA1MjCvKjpNsKCOcUjeVtmZ3UK
WLf890sp2WtzHcyw2Z20M8gl2kIu3Axz8XS0wYeVo7fdiz93amfOSrJ14Cn7
ApTlLSmCGYf7UkZ+O05TX2X3IPMxNulLDrK2gRWjgzSpoYuAg14RWAiDv+XN
v3wL7inwPZFJ7CWFfiqt8LKc36aFLRvh4+NaNseN9a0MbrmqV5mQGCK73/Rz
EN+SFqR74gF3GEw5u7ZCG72cuhjifLuovKlreStxPqUOjVopTJqtn4eSrwjs
mLTxSSqBAJhcjGWYjAVPcyzE6KMCQ00hlf7wbsGfcPGA5Mac83zk3Ba4+coO
lse2GXzmwjlnqekWfpDKfL1Ea34f9D4XWL8KVP90tTS5MK5AG6IdAobmL572
QizUIOWI2eEvdkrGS95ztb3UyL577AqwOp24221Lu45OBN+qlUQoh17EjUmE
trwPJ2cMQxkzkuf3ooKHeO5X+sxR5ERFOf98IO6r2zf45ll6g4AZtF7OHbUV
ujPKuV2JVtQdJlTYFVsFngKdhqlWJWR0tPL+Qr0w7iWP0rNCkVEqzGfpxOnh
199rIhf1+1L66PxZq7igTKVSdA3VWUcBL+Nkn6kAkJ2FYak0KsUPKIrcHlqg
ti+BEHasoCS/1sSgIIwEZX7chsdWxl4Vi1NMq1WpHig+cW+9Z3LyujsYcZwI
bAOMlPNcQOpaqXN0vw4llq9NUbD7bUp+4FnTRvrQJIKvJRdwNz3Qh9TVNmMV
0g207MOGrC+GvyLsyezZ1SQdTg4kundXZl2iiU4Co8a/+Y6SCG+LTNXWHvN6
l4qj88kPIpwtCTwpY6vQsBodaY018HBbRBaNLgwINAStcFKTeImwjRXe5Rjc
zxUgN33cpl59OK0xS6GWSdeG8miexH5j8kZfmIhSSbT3QK0ufTxxndCqwlpe
i9A6bS9W+bsF3rOMQ9bT40SnL/QHi+DRL7J/FaGHJPV2KUA8qZDe9mm4zG30
cLCspOL9c7RVfRwYd2jpumv0EccwKnu4TsCPiuiYdOEKuJ8gwCAsE+ZJ3oQZ
v6O9hGiUxQWAZcLC8VvOI4nNIquztsAUhmoYyCKCCxMfL6uVWZw8vnb9aAbG
8f1DWLHZsGx4ipF/A1mN/QPgGvgFlz6BXkLo0byVovpqr++GgMq2ldOf5M5u
XE8QF8I7cisPb4uQAUZb6r1rJ4cwX76IN71FrSYNs3ysXWP+Diy7CPFuajjr
YS3UOFcg2lYz6vC12xXytSRwXeubBt+W+X88mpio1L4BXwnNIHP6FT6XsrxV
NVOC/tnzM3cjGfohrnxcTCD7sRC0+jvhTt97WjDs4eulFpWmrCHXwhmkX2K4
G4aLWCeV8sfhZ575yhi53n+hyJFDaCz5AU4HSYUu7qwsJNFDVn5nPey5BmHM
o6vvEdWneXSqxacnLdQDfor9/mL4hYbI52Ik0eoZQhD3YxlvE8yKpn/qfLsQ
kvEI5ax7uh9EB8jeysJaDfp3i2BclPoRLQxphrGAdo4CpkHtri3BywlJzxZp
BxGg/g4v88jkZ4TVyskiOk1pwC31DM4IiLixCGX7ZSxw9DDc5SC2+kuoowa7
fYayADnn2NnGwFfrGglFvVxiIPSdOcXzeKOBKLFsCSO1CQNT/5FLyToMfli2
08rGMw651goEC+y48r1tAVGULazx/RVaQ0t/AgS8LNRhSQG9mlbLLzSolYcw
NasTQNIQb1Xk2beL8HcEKKFrJOeJhn9oIVfAVS1x9IQo1qAmypVPnUBEXUoR
m9py0Q7vDT0sOQIfqVECfvIyfjVi/hcuj+eUXb75MwZmopj1ku5F5vvTN+Uc
bszx+phiTzhAO8cIsJmwlTkBr+ILS08jIYp1QckBISTrgV5N4Fg4eclOMNgP
RUKD577k1fp82iNbOX3QgwEzaO28Z2BFUyvxZIrgUNRCHrgnHviQrcsTHh7Q
AFV+IMwvDUYPjaNeffc/Gz1iRKehTOkcOZK5LDwymVJBVgzD3NjigglZA2RG
NW71HMV+Pb2OfXvKnAXLvnie1w8vAvddhDsfufnXdTMzBfbb1tAtvaD6J4Rc
U+G/Tx5s2KYsKlwSsvxC4Ju1W3Seh/oaHGC2UpKB+3GacOAnm0Ql9P4qMHX8
T4pqeOcQ3GcCP4ASS2vfaV+ai9YT/NRtA1Fee+pYSZITHkeKYT4onTVKv4x6
wT58bC//eOM0Fd67opjJ60p/HpjnEhKv/a+k3FvskUtv47i8ldOkwXXAW8zS
JLf7U9ylQf5b/vuK8upO1YccpYqUcQdWVgsyQvp3vawuZpaZ9gj4rRDWOCUd
IoTiDGw+M4HVMOKr+JmTR3Flf6f6ufzXAZUwNBGJvaoeCUIp2TT/SnwcoMWg
aYKRjLH6y3C2kQ4cw/VF0CXPsKGGsKkrH4OtFeEuJ/t60QNTDYTIf1S5Y1RD
a+maaDutpfe41WdGJpvqX7cFZ8XnXf7zsDwW3HtCKkS49Lv/nn3iQAnOI/kB
DpGoVuQkjDC21mbCVLXZDLYIsVyO+DGWHvQ/boYwqViL2B9Wl/agG6BRrw9Y
m9AjuqLcFy2KeYcS+kYRy0ZJjcfZE6gGNi7ob5XYT6mWAgND5no49YQNUtsx
4NqYfjEfYfKjIkIfHMi+xMbOth2w2T7bqFhy1GmG5bpRxMI07ojEn3q6Az3U
Gj7pdm0KHxlYf77N6Wbr+lL8IGp8Ki2WylAFjCJP0nbUtM1oIRj7k75OZ7ye
5eTwJ+RW3mUkPKLXEOnjNY+7DEuS3rfwYb7KNYmpTsCYmZJfsxpemrJQIT7a
E6kBM7lDebo4OyCJIAV67feDpxPecEIt3g71oGolvyOgu3qiFtL8FtV/kcG+
MlsNs8ktiz5+VGprQjoTgY6BHc/D7iw+2Ac0+mXPrRdi2OaLNyog+DtYN1Jp
TYEpDj4QhniWS5SVW05tseIT+Vw03kTj9qZmYXW0pj9AU9yRYbZcx62qKRHM
p1R+CXPRn1pnL1vEViWCS2qLh4iFaJUcz1rs7Zz4n2ZGIdKRLsvG9TSQzOit
nk7WqZ0E4fLO295ae5eMxKM5MDS9ARsDE7KeE2g4E6RlReH3ogs6PXGKi+JR
S2OcIT5tdpUum14aXCyASXn+o96aXSzPPdbPaif/evedo1bKQUCtptfuKEOx
2y39ZjR+dBK8i9zJkrx6Rygm/R8pxiisDCbZRRoBhvKJTQcukkU4CpvThAMf
AMMYc/xKEoEVEX5xInjtVZzdqOJvWdw3q3xK6NmMGvHg6HedxsDzf5QQh0rc
6fd8ypGdPiz0u/crNmwyLTjsAS0xRVoQbtFphvJwJF2tk+kqH0pv9nVt0xnr
kGo9rYHfNemAh/KLTPTUEoXb/JjE3ap1pJ3f118Yku22ol0LtzkGW9T2X1YT
uUGgpL10OF3JP9wxHG6EdXyJaxnFEnGK4ttJW6GtnAmZzHbrBysimv1kr/sP
NRDWHPbLUfWf1ZJT+Ud/sgOZJ9Zqkl1o8vCYonMlfCUhho4zYpNmZdWybdJo
pJZiJhHwsnNIJaoe6pfaU4lqhmlRzOv+FhGHySpqm5w2nMGOvSjlYLxF5WXZ
tcjkROdcc9sq+gCYOnClxsNbEteBVQqYwVmtKHL7sWa2QSBqYFnqUki9b8/B
ACZ6ibX2oJ2udb+VVcIYxIohehomootFdyy+JTpp82Fce1H5wfiPSbi81dxY
QfScOrY/0OjFZdM99LwzpM0K/sqUb1b3QjaIAOJDHV16xHI+c1WjJ2F1eG8g
Lyoe+nod2myz5+HJs2VVWIfZ1Y/WQJe2gNPMmX1+f8RcDy9dlfJFqNQYy473
A/2IF2BiCEUHs3xAP37bzWcPvZhQ6c2tEYSVsJXMic3r3E88Lmyc1lGLFOj5
8i6kQE0Zz77h2hoEDWAg3NkR+d3MD5L0/2s8w4mFb70+3U4eFQcaL33w0IRl
T9dySnDm88bGWFwD8KTI7v28sJzGiQGBHyI5ySmQOtaFAM5LkgPwi9kuGc+/
X0if1ApC4zT+LjymvYvJPsVdmKgdDVMBEB95lXHKigPezYyqRBZRzItdl+oj
/gKV8g3Q4QFKBw1iXbIN/rcdWV8yfzDncADPjM5RbsoGXsNOdeC/wwBOW6IL
woLiWhzsTQ9dTKL11hCrl3wIeIfroTAAI5yO63xMSos+/4df1eeSuFokBr7X
yKFGcL7frjiAYDqOegn01w+kVOZb14mS9CilF2+AnRz3YKsFYNW4esQfNFMA
AvF46AbQZSLWE8S33iooZeWEGR6R3adESZu4expUcnkkGYEwReGSOk8j9BbE
5cBv/8Ee2fCUl4YdrRuQUlIPvnqvtfzM4pCkgf7SGB45b88tH4Pj8VyPhOtz
8PasIVKBKh8041OdbFewK01fJ2kKzRbAbt/xElNkwzfWn/7l1vktz1MIcqw2
4y8OGRqtqkK1yjJns+QDcNrD+og2UfLHpQIg2AKriBBcngI0cevf6BwdYJnG
U53EcHZLuCkGiJ1adtVKyaHpBL3d3qytOLOqui5/2aaWdtLDkogX7vH8T+IC
5YPNuSjQoC0hjM1ATE9fD0TfpiNfv3iDffLgmJF8smrU8zIyN9lrIPfj4GRr
6XUydNSh7xVXPjZYzdW+4gBpD2ei28+z7TMZvrmyIZ2w58HFzz+UzekIcgA8
DDVaUBuJWGjRKmegLEO2Ksduhm3BZcqT9dj4kb3OA7XApDRwa54F67SJGr6E
tCVWRuGpDZGsCQSJzJixEvCokCf0/yp0VwPRkFQz838qOL2Opkj2QxriPUIH
6IFlXszf9c2JkuPvbU7t3iCUiP2rLQdbRBbtsTxBCBUyA4Ojfka+g9PbYjH5
QYzwtoD8n0+qCq98lXGN9KNZkXHKUjFPVJ6vD+XkwmEdBLcgovAlsg9uZ9ZJ
/K7p259O9xEJ8T9wvbHbNcNDhhPLGMkxBsgvdosMp5DauMf76qFBFkYrIbxV
YCf3jYute9mIuqFlf7XuhIoCPGXSBlA722PGge4xwowJFFGVZ+SiBzVjTQE6
fDlM6ux+fFKTHwqoGHCowQGtC13ITGu+8Yl4L1D+6WSE1JaR4Wx22Jwfs2Hp
HLewtrw5Q3yAs+fmWdJrKu+7WjDyncQMC4gRg+x6Kk+h9NNYk0B+dUWplo0r
O0m/EqBP58B21ORbRJNjci5btdtQUS8vW/BGvWpPF99M6deaqMap6UxakLxn
7NQvJYjhtkU/+DAR/sBhhD0QqFSXDmoS8B2EnzhKU3fxd6NnArjN6Bi93ZUl
dStiw5/cfS7ZyCvc6YmukgPc0EWeYRZ9Rl6wQAxB/DMiO7NKt6R1SvxEe2ri
y3W//MwSgXEUaCD3CF5XxZOb6Aw0QBiRVZVao5rY3ftHSzzopP9nm9ZlcLz/
j2g4xnjdEKD3l5cHvLsFXcdsDpYwRnNu+jAwmPnXONaEFHIYBmnB+GHl0R5H
lajU1GGZnEDR0GE+IZ4ndnN2RQhcyEsyUvCLQPwZW/O4R5YJ3dGFJbz3QxS1
4SdDQhgoU5GCiC93s1nmXAhD2E133C0bASVed9Tie08sEAXlJpamwm1ElzS8
8UguWl0qnPIuBvk6PW0AG/b6HRBvLQ1bVVEAtgn5LdL9SOG4w5vaLy20CwPA
zLjt2MKOPOIW6yy5iYQqssEhhYXdGz6dXgFwNaqxGbDjTCd9QY3Mj3F7kwjT
9UvTDMn9m3+EnLBX5TjRmUr6iskoZ7TGWnpXWBrXDtbzz3yVICmkUcyFzkub
Gk28ka+8YnGxXVBr+YqvYn/2pchGb/ZIEdA8dZodKZlM43faJDzrAs0oWc4m
Qz9CqtCIdjUCQS/Q35LD7KUPVHHMDKTI/8fn6YPLikmPYfbxAFnFa40Da99s
hfxiMYUUKPrCIKP1Kus6w6V/5jjzuHETc+1+GisHR7HMUjAnT9gBC/z2/4g7
fL/EHM1rzEixjPWIiEXTozQ9iAb6fW+xQ6QkaASY1NA1H77XUkqtghMsp8fU
jJnj74Zi7FEwhcbRpFjrQ0RA+SzLj2yZdBW430XU46m64T7Tensoa84llW7s
pd0MxQKTTUXNd7uSl0vPQRiRehFPOxomX7p7Nkz/HtI4dRp7Aqls+mABA2Uh
GEwN1E5gpgMEdtazfZAMfdhnIDvvmb8xmjDPCHTfSOTQCA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AHFS8uhOzEEv0qANUjCa5shxFe8bemKFNhQTqRGtC4pjovR6jkEwCgEM+HVx2+RETJ81jdGctIsI8rtsCu4TOBbfINYgMfPtAhYoq0pIwXzpBYW/Jwh89yYqmQ/8qwf+UZ/RCUPZ9uTW2DZjLM/8DQwcPSaWPn4uluTziVOYaXqZBjqnFFKudtGOgi9fUYcdgmgi1Cr8qg3AFyDXZaw0JPfMHv+sI1tXM9FJgZxRxGPk4XF2UdbYhvlmO+NvkAHydQypTXKFVynjlFLskwMPoQMq23bVGFmxQqRUKSGYY0vsJ3YDO56JOSvZzXBbLY9utoglCDlhz5VusnWjWu2vn365qatA6xqZXLREoeo4fK04hoGg6ppFEbz3Mym+1UkDTqHYTUH1MuMg1pyE6D2/JmpT1yGxfj9t7KVXJnjJazVVxX0bIm0AivQrzui68/ZBAtrKcSs9GnAFIujIySv0B7cXRNfdg80cHjd4llYwEt9/gWKoRB8uF1xZ0pSW+Zm4Lum32CxieREUuB/g7BCVMI91EzPYUWF3oFPYTtS5w1tENhwRREn0TXisyMJPPj5JNFSHR8LEtw4Xba8HpCM03467Zn4WYMXIPhURrDqBQtIHPAhc64kIZHCXm94HQOu/eqEWAzg3h0ic7Dlnjlq349RoSnSpcnkAKXuj/c8IpFVEkzB4jodlAPvp3rsIfi3XnJCIG0At5nKtQsNAQ5QPAD8n6p10WVFOeCYdwIAVqsOo1yiBT6CCmEH87tcz3ila5BWwsUnTkA2UV+ezMMbOkjLrwdbRymJny4wAdXi0tuf1/sPUJ1btlaSxCGiGsEdwkDGLC8KN4Ze0CJfEvAEabdd7s1bcJeaUbd+MZyLGxdKi6CE83AXDQgjcb4ycPMQwg4nHXXfQz4zp+zsgWKawUxcPAWGFfG0t+HNdf/pQbIjtK57/RRZwSws6maPu4nCl25KhUDFaFXKgsZ6zbT7+N1L3K7K552itq6Cl1h568HfoBpEO/QT8Zs0VRJhMjEMN"
`endif