// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
i2cezSjNGDOofLfZ3lIjFkWWqWIrwByRrU0danSS5TM9JUqb1wqkGeQjXvDN
d7u+715pBXWUNEg6jBPklRikU83i1dRhJu+tSuvH2iYG5VuMv0I32bW/Sf/r
9KvSFFgEnf5Yul30ygSuZC5rfnpg6oAMXpH8bjexvjPTAWSh6TW4NPLteOZ4
GKdYIQPcWyCMGH9WUIef1SKDde+2htfGirLE+3DBvlMEfvAS9D1tig7l3LYZ
RARwusKAKElRX/cHavKvo/WtAcTzNpkzwgRn80kFTukBB2+gG6coT7USWd5N
BvOJzSb9e7VMVmqwTrjXHGpzh9cbffi0tJ97gJzeOw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DXZhtFP2gqgkDaIQ0UMGDbHD2G9N7tAbk0yf2qgVbQLW/On4TLcefnqTHPV0
ncI7XCtQWpVll68m2Z4gAlkJKZ5lDGCp7X2Nj9T8PPwFsSssUe8QmGT0a8t4
KAXmR5CZKQwP+/uyOQ+GQlozaGm1eDk7LeoGo0Qj+la/d2ec8hHusWGJm15u
tRu+j2swgpH4eUGJfD5r5Ek5ObnFy4egV5v6RaguyRbM4v/r9SCIQFqTktlu
XxF0QQPqLUNMUIIxDTrbEXzSMXRw5bkiX70mYjUrmTfajxhY56CAzfdo8O92
xYtV/B1vwQrFtywxoyMA4tG3OaMfWXF5EeqEWl3GRA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Mn+YjOv9axaIOESn08iFLWWCyHxA9PDfLU3S4qAsyoHfPd6JkvcJqcRp2mM0
o988jCn7jP34YlDXr5yFl4CTZxcowYfG7aHrsDPMvLFU/NUatjOhgPBXMNXN
rdViOcd8cZW3b0rqaxRQsHLOqL0BXbeEbyElBZ1fms69wRVIGqUAAdkgcXA3
PZS9OiCzNhROVuqkTZ2lIaRBj2NC/evDMb/LEoG9Ln3yTMME+mBbUQe16zR/
+VZAhjTnrpJ2C7D3jRdQP7z5knee9873/HcL7F76wsspPAqOO+aEoFoaADpz
sIAHwih4S/xBjd2s+4PfQUDPTp6V5pW9HAJQ8gciYA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
C5+TlPBQV8gS+tdFRZvnFBPrJ8vbIJCqLlMxKfAWuV8TsBU8YmE9L2NswjEr
VwX6wX7oFjl5hf5hZFz0OxydjOueARvBjm2aw0DN3JYrwxf3eU+iu0LiETc8
BEIlqRddVjO0/MBKIsKKbHs4fjPi6SNeL3ytGwPc8+rBU3fqhfPkWlWjlUI0
cti5GLUo7JooyDy+eGLfpCX7esijuzQqMWcyliqbdgX0V5En+OpE+u3oFS4m
bS4SlE7TIlUcQc02/jH6isMibWOgVuEZYy2+rfsxGe+8aju6YhdC+OrONhJH
W2usRtxu8/NFsSglOpBSfeZpJvZO5GWgl/VGfYOArg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Mcauc/L68oyffz73vsdi8kuHb8uhEM3azXGIZ1q5JS6sPITEAyBcNIten775
ldCiEIWagtKZXN9scZ3io3qgC+NF8TTp9ZLB7gC7VF9HfIS27hT2GSweGwuc
yrDfim3qxoupEf7IX8cSkZrrxrdRIJEGIYmuIYatTkhXx0vnW44=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Sf2zJ1qsZuRCXYn97Gd4dHT2B6JLddjG6sJDqlo3vzOQnG9GglpV3bi3Rnlq
BYF/S2Ddp2brHA2P6FBdeCzIaNLx7OiGeXDOMDd2e0uXmrzR7Nc9kTttzw3Q
VZb4v6ujRYBEOptWM8ftCZTdMirfaZbHpscRF3t1zzYi9N47Vb0dvqx4qiKn
oNSk/+x4ocN11he17diZsYt7AhI82Cp3JGRA/45OVe+e32CzMR9eVx671D4i
jTULncVZuzNOdeXsOA0UM13pXna/Rpaa7D9jd/VvwLQpSEYLu7QPqkwCgNiN
NtysQ0vFkosgOD2z7CAkcQQjzURDUtmPGd1H5cd3LdvA+7O4JOU3rOFjdFJM
dcwzlCRgjRzKejvU8QISOjNoO/PjsXJJzyBcv2jHKCGNBvrLhRG3NvYof1ys
6qluNxKeTPqpea166nennYQDYhZu2tGgCFi/dDuAhD7X3vXJaDskUVqZ3vBd
ILQQD81aFHbsNFyMVdIFVlBZiiHu5mbe


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Uyepg/YfjzJB0+lgY6bA/zV2cz4TVJBLjk9z+IHsKsQKMke1+6IKvcasywL6
eJIAQIhVP3b/Z6XPjmSgjHlsa5ASMqVe3wMGBQ7rPIWXdcG+NJwo4kvubyZj
bzP+vPE8k+BTaGnR5z7VYe2/S8pAiiBglQtTHveEvl6O2FXKU0g=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qBURNAXuyOYFmoAZJg1CsSKJOL0oamHLXH/tNocZz219bXWj5t4hBrplAg+1
BtIVVGbMm2dYm6CO87NnOqlPqszLAYrLG+0Hd0DF+pNkMwADjas+SAXP/L2a
olLCs1cTNx4J+/3RpjE0v7SUUVIK1F+xkagzBtltQXDO6fZ81bo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8512)
`pragma protect data_block
dhXTYr7H9QAYjfQSB7bUQ8Oo8UgRRJytTRwuBJenBSH/pORm/0IBUcJMUHQA
GZUAUFJc+ILV1tNoKK93Rcz/T8ysrxr9RpLXvna/dNWwlCI6nr+6mq06P6dD
TGF1hCtBBfK3FSHaD6PMgXApZEx8Ppalb4VFDjKKz8EWkKFIU2CQDazndbrD
nZN6CO3Nf9gqz1QE4ImgQl/eFgQSR9/Jl3KcpHRGKOCS7GDKBYXPQtjMaspY
RHTMlMU7WgbJXSW2CQngWn4C4t3VoHxQKRlKsBiQtNhDssOM/pgAZCO9Tqt2
RKPsil0H9fAOMWEPzEuGovqJJFdLr8JBm8pFrufFgCUDZ1rSMAgTSRnPa4sV
f6Es2rHCFSvhOU1csKnoFx6i50qows1qcKwZft92FZM/RgAGVUKLBkUk+iRL
7f7DeC71Vjzw23Xn0SrEllUlvplgqcGpjRQ7bpk6gEWnDZGtMu+J5BUo/hsU
xk2bYquzHEm2i+gkQhVnuq8e+fV3SwMYo3iqQZcVvwno5e9hqvf/TfjyjTux
9IxYgQ76mdne4NOGhkAkSp8Kk6/hqjw9yHBFtI6szEcA3NeSSIFjRooeDyo2
PfLO/uu56HyHY2X7cNBu6MP8UkW5uWZlj2iTNSc/u1/5CJgI9p8yxV/Q675/
VQzaIpYBtolpqiG+RFOkjUXMKQnDPwSQBGer/RurIfF5WWfMVnCDSrkJhgRe
43yJKQ74qFewozxXyDLEU73Rvm8c/cCepll5ZXv/yoZmilbZMxyXfziIjCf6
AAq2zI4V9Qxu++V7nH1DgYSPtCubz2Ms3MAvDTYMuuj7M+bpXlc8/1acZT4v
2McG/lXntH4rijbUpfnY4U/SMWcODpKXpGiCVeNxoaUKDBuCZIrn6AwCK2Bt
VSEyl1JwsH9CwWcy+e2i9KGa3fxNHCFyf0Ox/TCIDQSjp0O8Phbs4bcDoZ+A
b5nt8d/K9Ixrbwv+BR1fbxGGZT1uLybHpoAnJy4aX5g1MWDnWhXvaDDAJZRs
L11LuZwGokXx+CVksFbhj86z1Ia9NX1bLTJcEYtflTega0ayuKbABYjNiTOj
M2LUoF4WUB+fiuAcPSnaSweKv4RcfuC3XpFgGmkY3ijGH1yDQH66nfB9qcwS
EhGVhId0OpZz89FcPOtdKFnCoi8Nj9+adaWxayyps3JPJGdkc8/5V3q4SXoT
5iBn/4ni1XkIwoqw3cKyMGTiFu4pLA7rI5kxPRMlhq+C0aqcrO9/MRVhKCjV
kqC81alQy7qiOuUPbgBeKH6jElSEWSYhT8mc6o3je/12y/xXdvWDPdDb4duq
PXQ9/xd5u8XIrYC44fXaSIJiAp+mDBt7/d054cs2YyPtG5XLBu3HLPCXLAuZ
di9c5YVpICz+jJ4UfDcLv0ZWwFgcfejORBIeTMKpQoi8nkjH2sVQUAjbHRqe
fe/sAc+cx+yac+SMPZjkKiipN1MiQa5dzDhXnTIRgfE60ul3A+/K2ci0XG+y
Ggo+9L5iuJ9FpelFZAYiNARwvXcGp47IFcjTO287zQvQsaL1SQUCmlcvcq04
mIhH69Trv6968NgELH7ZHpiJvpdvGeBTfdSxIr+jTq+FYk7PgklL7MlCgQMx
+WBz4qF4i9aPb54Yws0xm+pwDsyPZytsmYxqKfCG17c75ZpAaNl9QIHUMGBs
N+7OOedXlalez+D8I4it8NF8dga1n1JROztgtYesK0JA5ldQ4tiHFbXn9yAY
rcAvdAV5HV0gkhqfxgo26rHS6RECqxFrCBZDTv/GyCf0cnHMsk8vvxR6kUC2
c371JRdzh4A38I9eWXYGHs1b9hvtqreCON9ilSs4XJ6MpcBSrnTwBt1+VIzX
+kv9M78ExPgBDh3X47ZC2GJbq4swEKiM4wZ/F4ag8gAGLJOxQcNI+RnVPyfG
EB+m5vwb4yQZ4ZRA9Wk2aBgoOgVXKlN5R+kj8H/nNQ8LjKWWQ5qAnoA85xHH
j4Vgmi3Z4isAN3zYIvFLt0G2x3n74h8hY8WQrYLAOQgniqtIWUAvabj+KNb7
Cp5PM26Q6lOftWAf1IV1eJDmZvnvGA3g4k8c2gpWJRa94Jj+rbSRn2/cg4Iy
QQbeDxX8BsjkAvVgM/wTrH8JQJQ12VN91YFppOABdVFRoPZjRryC9l8y97Hu
oPMse7m95lrNEd0MR8Y9b8OQRBzvtUqalGzHtsDnfx0ZAisjqaBy5I3lH98y
qTVHkM6aUL1/7r43P8QV4nbP/zLl/PGvOqiR+xjomQZRAseSxtXfbFekR7vP
Pv4QvcoGJhIz95DTv8cwjcxL2KGCHY3DCRDX+zxAoyxB+n5EKZ2hXABBl/Fo
zgc++P/csiog0s4a6UYvJwvH/AG8zR7mBGAQmkDo6uOzJCmuvOkg54IAGFkd
jcxTIZulSI/5KM5VgKI7dG3lEoU4cEtKQOqMYte7JpFL1iaszMR8+dKM67x1
ADxywr0h+EOxqcdCTdtPYM61nI46SMUTw6j4Jiz5LI/ltF4E1FeN/X5PDSbF
HboVPOh/9IpaKhk+Z6YJwYSeU9IcjW4n37FDE5x6Gp9qt6jFFaUZ75GzW1Jw
ZLJstPqbXno0Nt4kRNtVt+DjuQ9XvwiQUEDm4hZv9T9/8rZbS2VfJPTGyf3p
n1k1YY+8CQ0VnjwbXam+DYXz4KaaeXTedGGwMlsUrV6iD8aeNOzy8eW09Osv
4tqJ9ioEkxZNFz8l9QTNL1cb2D00R3lPBs06qySJimYbljPg5/RxgM72gOM+
garGGyL3P348bK1GKboeWV0ogJadojTSaBS60OP3tkjWZcByJD+4ttcy4Zcw
IraBZVgCEMjzk2+s9ODG04vwaXgSwwNGZG/OE4qTCtYU3PhmMVpH9PZofpwt
LDsF00SnjhxuX6xGwGgYRi+uBQMgFUBy15YFygEyXRPoD8vY/uDCh7SSMGyb
hMy6IfOUub7zkLWxAzvhH3F720Rxz0kJ0wl8+2N/AkH05vM8FKOoO8KWtU0T
Pv2RkigwxQvzRCXByOPOu7XH9pWMNjk+VKRp2oZKr0uSQrNq0GPTICAlc30K
QIAEMs67jPaUs5Bi9/+ta0BJKl3Tor+Wyha07/ziBXLDKxx4xeADackcL5P/
XE+Miq9UMcwop0ZTkUqFSic/ePewHVTqe5caM0NxrzU6zf3QEkiEM7Hyd/Jy
YBv+gO+fu9PtthRX6QEksEuQUZnv4sZbc6+Ae5rBZbMnU5QNZgNzzz41PTUr
VKofYE0DdngAHRFMAMehqzvZcjbfY+MHnYPw4UekvWZriBTw00Rw7Nw2eft2
jSjFXmCwqubvqUKZlgen2C/3gyNi013FGLehlFKlnbgcJyk1CdPeUDhAYT2V
xwre4rhFdF6fBHSg2Oz5qkHrfCn3RrXlMGYksHreKQXAKJ1vXVqKHWYcTNu4
L34xN6uBH4H9BDWmATWsfRfGLcJ4Ye0kOlYSHUOnF02aiZjAt2u26e0oh8/O
ckvkMtWzTZhPb9VPIFsb9cjGhICIAQ3cIfBIBN3xcG/RLlF8QunSHHDD++Ii
5MzqbuvZeHzbeRWLk+xc7VIdFnjQ/lB0YWJt86n61bk+WSP0hFCvXPY0TjYW
bF+JvDDrkhmAW9rm0oqepEGPq3STutrVgQaKyfW5oK8aPCjesumqqepEmsTO
pHEYGQ2rpt2n1fB2Q0ZKO0unkAKOl15CEc4cbHTeHdUTCc8jOrtQIRnG7t9e
4ZcQ5vAF45wKEmQE2TY+CvYr6FngSmDUr9rtOGceAlOLjnfZ6GOy01Y7jkEF
brv3xKNXiYPfRa+tUSgO+FexuTOQcXba0fl1s7rGPe21SfPdVAxu83dqLL++
SsIc2WX5s42Cu9G7MzCdwqxuIoLL1PP4oQj7bLGnwVcVn0LWgvTKlj51rRmd
g9+862MNxuT7G6eTTRMaAXLW3QtxkSYqIA8cYdNVqo4m/oOmRRvs4uyOywn9
SaWVsMObswqyg8QA0GJpxWWDVV/BX1OmZYW/ELyvYYQpWBn9xD5EN+q6PEu3
06mcb7dI0TAjB615tBnLd/S4u/zgfRFEYnMh922vILCqb4r0oRt+YpW1QD4O
jKWcqrsY1SAex9T/Jq3ht0ZCSvtDfoVIpwlYlyFeAIftpC86p1tG5/5lQSI+
4CyOB1H/OxcZgSDtLVfpuPUrSc4M1+gW1vAneJa9jU2mqjA1U7RHJcDiqv+M
8wOcjWU+6nKwUnWa3gzrg5PtHz4SbDNY/g9QYCuntW1iPlQXDZoz+DIF2CVx
BbjjBjf4dcubtlFZxnYMJ47jQfFvawgAF2EAxJifDSnHgz2QrD+xQhNAUOhL
u8luhhbUnWdvwVeXNMmE4vUuqkWkQZzShnyyBEOR6fshJfy7EbEBEM9RSKl1
TMv8+o0h1EP82xqcg8NZ0GH8o3ujBwQSb8UGQB5dHYeARbfSIx2gSh3WlhUp
zrvSN/OoajdzvnVS0MNaVJzQlsFlZz40Lol+DxFNBs4MEGCeX1dgoFLDoNgn
SxY9CwkLae6bNeoOg5npbyVsBi7gJUssbPKp9oCwOudKXHto8V2YCGV0etCw
S7LelPy4TFjAFn9KaDfGQHanB0ftEOiWRfxjLU3kHAs8LWyuCaCWZ3hu+eqC
X3gO3QUiZRRmLcECHuzjQtj6cyxkb8l6+8mHl3MQJ2JGR04KEFqN1n1pDTmr
rkXFF3cp1T8RfWW0MlOMynK3q8LsePq5e9ItZSQCs9rTj675+HDNdILF7iAi
8IyQ4mCA1lg4ZD+KANrlU+it4s4xxPwLSdobGnQy8LhEHwSHXx8V/STOcmHN
F7vfKKb8SCDYtJgD+lCBr/1oLMbMEC6kiC6E5bGinTbn3gUIL5OgD38J+6JK
kxogBbwK+9kncmJDgq7f0lkPSKcLTTbH6EjfTp0r7VmQHKUSl0xgpP9JFekA
BVOqj1Hxh1phq8bQKoFg3P4CuQhwuW3ORwHgN2hWYeTOpYFeKXqyVBTBzXp2
6mkdV+ECynDn124iQrRG3O7pu4vVfoowElr0WOsL6lVjfb1nvzGB9XWzzCjq
3C0JbLmtTe5IMiX7/xgDRxuySGR4Rbgmy+WdN1ZQlLlRp7qNXc8h98eBtcwL
I60xB0/Q5HY/wiJTb6d++ktyMFPXSd71U2qsyCWa/E0Cwv/1sU6IY9UAH9zc
TxiJVLpnGlpxtyu1ciB+/hC+dxQgP+IizM6heZU9RmgzoUol6viThM88UlwA
Wwdn6RN29LfKJF27Qo8uC3C4ZNDrXLciTWrWJiwsrgrIUOpeB8w+b2KmXWB1
6pyXOCoH986olGcgY71F1zRLe+HunFQfnsvcVhonhvFPpYaRTQoHyNoVm+5u
GqTOe+wrW4l2623I8BLMKcWwCWRPxjBXwUSg3/pvw3gRNVTHDjC/fiDhArB8
SUuJQZNtwFBYTZR/S+GsZ5HS5tO2p6txF2oZH74WYHI1uaV5nIegqffMJa5z
F6kLOaJugz+ECyzOuEeFbJDOQkKBp1vRAxtNF2CiUcHT2yz3oD38Vnn23Ejg
Z/8BnUEn8vIc6zb8ZVGks8RRE79uGAYNaBACRPMwbMZTFZyptNOpXc44KNRs
+CFq24OmSxk5yOSRTilDi9WY+TYRH6bfPtHJGJJlrEi5a4+ehPMFCPhLyfyY
qoC92jWX3Hq5xCf3aiIznQYwYj1LsdQRiIZfZca0fFKhafEc32mzpxrtWTyS
tSyzRiJXvstMN7HywXiQJy5ehRR2u2VofoPkDoUh4d56gcE8IaVCuzRP02I8
UHJr5uirO8MOd2xhc59zPtYHC4OOxbFEAUKIKH/BpZPG11HJ+OdW6ZvaLf/Q
MEdjUPwrmUq80TaythcZWSv7L97m0gssWGC2V0Uffpiwv9HcHT2srXaFqG+A
Jg4rIuBgfuzPseOHBHDiQJdkUuplYk3vEjCevNVJDJJSVlUYbLA1Y9pNAj46
FSuqNnjKNAtGe1dRCmL/7tNKcuxLfWJh2LuGUfv91P+9kaLD+0+0Th5Jr3p8
zEvPOkBKuehBMYzuaR1jQN+NOQgkpt9afJLoUCey4bq7tkdL0bATMmWtSCCq
zH2BI4jK6pj+uXnSmnTTMPoDgSEsOHwu6S2mBoiwY7V3Ok1N3FQqzzPeefLM
I787Xy8HQl5oX4TZWHeKpr1bxIKxQilR8h9Xw2VxvQeY516vgnKTaYvITdIK
rB3cb6kxueo9FzrIXm9zbhjVYZFrkGbCmoBpfl3Pu8pDhHjeH6a+R4L4+jHK
2wYbv/VF8ueCk62L07w+jQVvhZbefLu0Mms+ja7Z/SYBPxlyc+/RrGRwxqML
SHDzISWDVlePZbCimS1Q6HV+Kdb6WU21j2Yv8Ns/0yXO7zyj4Ghc6f6N5jR8
4EzIWcaP9QdI6Fl5w1zeibcQTVVFKfILcUgcD2D+Rq9AwxwBtzt/1dVCA/Zw
RymlSq7SWYsCALHsD1zuDOTOwuEwwk10MUvL04icrm5WNr3kHBE2lOfJ0GXN
oqQthk7UnGgcsmS+iUrIydeZVUiVXqXq7GFuhAt6uYp83vddg7I7ZLC2nhgX
0eYQvAHeNq7WjKCGF8yrbRbqh8mo3V4p1eNx6NABotgdmmnuTiYDJrtRgXi+
7+ytI597hDIYaOTBWvwQfwwXa6ko+ktu5+PsglYX4gqYOlxOCiBwCcfEtPfL
a32ZnkNEllBVmXDvSWv/bcmv2F4s9rUk3pY88hvjVUCY3jBep2JFFCxv2pei
S9DC54EbFEDAolOv0mqjtqDZoNB1tgKx0Lo5NESugawK16Oc231n5sMttFEv
hV89y7HNyAVNLI+gAjn05Lqk0zhV3upZhrFMFmuF5dYiHj78aUke7mowaaXO
Lz18Q3zRphtDoFW54KWGDFPe3tnOHYXPulDNzcyvE2ePdKXUJ5iQQQJaU6if
IRDgvAYujf5DujJxNh/zEzUyM0WrUjSjAsryIJyRhFQqSx9JnjpiA/I3KVPG
hXp4HSdzZcfsYfvNzLRS1G0Yt9m/3zQpSZpCaclgxtJEgZx7/q0k13rrsAJ2
5f0VUSFDQ1f7YZJK5Zy8EHPdyzmUbQemyPAfFOhoIU5nJiOBAG0nBOBv+9T8
LsR8d27kyziNG5IDylxLNMRRUogHBLiJY9Ra8X1kKhSvcMyBOsZ5BAb5NWlI
OLQk9uJ9I7EG1cxjmYn+xicZ2lCJ0rmqbMd4EEZDRUx+TcVnXzXV4MKv5Y4O
DqELZg+xo0TZYnhhgX0OV180nS5rpQeNIxetwgPkns4XM6PrX54q05L//5B+
hBg36/1EYOwEX5IYoekmfakxBjlyCudZTgqr/4YnW+WwbF2ZbmzLvDNyfANd
/RI6Fl3ohBFkHT0lVy/kBXS0x+gOBMPdv+TR8xWHzIppMLakIa/UnkxjVY08
952mHbjIuIuQsonFMU4AvawZIteB4Xl3eUvJWMoKN5c4uHB49FHCylkNKySn
THWhWDdwyvUCN8e/9DnFnFVq26Ml5JVxWv1uOZYNhrqV3AWPaQafW04c7b7j
1vGhy+Zyr0W0KFwpmfWJZthmNRc0KmOSnLJ8u338GEhUyNEpaXZdhZeIubI/
CRDIXjrb6MlCe34aifLD32+5+1rlfn7/BtOp3PgztyhXHn/RkkSJBRN0SKR1
VxzQj52nklJWaVpVWWUbKHkXZCBqt/lBNurXxP4rTML6NJyk/Bfc0sGNsPWK
8IYtRcqPxBAMlvf9rtMas1JQsR0htpetExYCAymiZD2nJy3M2dAc3jwzWLBk
3kiWwENDbU5YzIqvNKs7YXfjj4o5x0SuenvdR7zEdpBZL413z8DAONKcTOs2
Zs4aO6oJjcK32Ocqr822hVVt67jxxOmuUe26SyU8QHBzKycyK+lADksat9IP
LHaSwUxnoBqJcEqfJ/d48zCVBE1E7/ziqAZHosqFUqo0DKXmNixVWb+VDMZ3
XtIF+2bjvwjsym3ikp3pViFa+3MPCT13YRCS7SLGdY7Kfuceg7utlrFqABtJ
ZSGI49QAfzQo+BVYmpz6Fa7Q2G7xm39NxxNGjZ5kA5K5ph0JSDpNUfrWjNHZ
9XugaApRSytTAwSvHL9QQyTIJ3gEHt7CULm/YgtxVwShcB1Np4B/MrHeJQc9
OTzOvmZPTM5b9qmSKo3cJPqc9e0fiyk3WIkLG3MsL1MsQaVdhdz3ZzjELUIN
S+MNZsvf+ZdlF5h8daYY2xqqN0Jcc6km8GDOT8GGZC3pbgJDwACIL91YZnJ4
Fa549l04FYpVm1/9npmNEK06brXIY/4rzZIQw9OCYTNq45wWpXaUK7dLwWjR
29B4HvgkO5q0kRRBG34Hql7a//maFcqARyBIBoo8OvUl2ZCJIaNM9SFBNR9U
ZdmXBuyTXDe0i/U1AZuTCrzvaY4GW5t8dzIrkHVfNxBRdKLBkkIMHpmy3M66
TEo5l0MZ5C/dZmHYyWyT2g0KHo+Xf1kMd/Ngfb9nMXgSwR29Py4K6nx0f5R2
IyjqUoIhNA+jmY30ZO6FyrH/BME8h/SoDIFpldIB0XU5itpSjfnhyHP3xY3w
L+95R3Zlt9s/6bH9+8k3mx+AWD99H67+KuqoF9xDkPBvOnKfFRezSsnQbJ2v
PfYHfzCHom/f2QJqFznsl30n+UOx9+TQbdDl/YvvVheewq3lq5QESuUidqZC
7iqrQGFMY60jpNHgDIXfR+F7E6UjzHZb96EVF9nPhhVuuBj/3W1VDKTrVhs9
2xHsgSg/tS5FDM5al2EgmpMfzTWScpgLd3xKabQwguyTGDuAXbBxhUdH/aRJ
iZW8/CK7AfY/ZBPnopBuepiXssY22yP9hzh3Bp63mRwLq1EjR47t42EQ1aev
LP5HQCyxHAH2DwYln+vuY5K1/798a1J2wMooHxVfUHQltMCQ/bFo7nVmeX2b
1G8Cat3qFxKB1SqWz8ksHBxHoQuOjbkJaq/YdswnHJ6noomYyB4EmkLzbs0D
RoyM63MQohlU1dl27D4W3FuPLjI+4xfhbUEICJsKjVAGlADncM2ioqz7HJVi
9uq4IEz+uc6899pJPHaDgMzr0fJh6+wUapu7ypx8NOXMHsdRqevi5WuK9dQA
eftD7xJQqFLvUyb9CvSeCtPZpPdgh5KPag6OoK5Ll1pZP8rxcumUC1F4EMDn
QK80/lzt91uRGEDzTOts7U3KNhNoDl+WKyVhijr9993T/5ytIWFPAqZx0wj7
XihViE41dCsZ1SVsFWJUrqEvJ2KeOZgXmyUj6l5WbFY863c7i1A951cosRsh
o1hhX3HLJ2mpqkQ7V7Up/X7dttk/tv5//Oz/jmY3ATnmunI6AfpcSBKL+mzr
TZBaWjCoawnMUGfPgzU5oExV+d0YV1/n6GYwVYasYCfN4esR/0Sk9197nxuJ
OGwtFBH8+ttYTXt8DXvF0x7wOTBoe5zwLCRgTjG2WGFBm+Cw+Rm8rZUbQ6Gi
FqRSBgQcddJHZk29eWIQwwRiTqIOYHBhUEECsZLQiFY/nyAS1kki6Km35TpV
2JGskAcdzOcCe4IYCzXKQhepN01IW/IbN0nOWyMYrbjezqYkqmLXvMWcefHB
TquVDgCXpUSXSr39oIz3r3Y9YCHUOQbNb6TpauNX9hD5TwdPDiFCQ9uJmcW4
sJBP4o1L/ufwdWmDx6rYEtgMcF4XOglbowyNRsd78Xvw3XovD26u62erBf0U
gXddog3tvbr7lhRpJCKEhuE8X1nEHNdRHef53NKpCoo2A1MGIjoRA0STyb22
Dn7XMDsb8fQbNO9m3byXXXf/b4ZqNvjYsqJCmOQNm5fF6oS9has081gReQ0M
c39w5Ev5ptCpcuItkkIGlQNIYQv1otPFHeMBTM3bEleShINfj0hxek6fcLVk
yOimipltyeR0P2RcWALMvTQh/Hk3yx4B3S0ZBCHQhYLK+tbPnXB9A7hvTL7w
4MJa882ARefI+QLgRo2s535OGfScyRTTxqDqWBU7JQKMdtUzy1xQ25vW/zXN
1/AEJzuIafkuK6dy0rvbND9IEWxNMNRJh0LK1ckf+qdXbthYRVfYds98Z1GL
Ldo+BzD6f1BLgp59ARJjGhAPVhahlW/xhodV7DBLT3cMFIxSsqww8aD/fM26
R/3odk7EC0jGVnHEDMSqrHE6Tbrn33SMvoFQnRfzhMeoCvF+AKVS9UTTgLWo
wJqXgn+wx3BsrGOSrrjdSSc/Oy3rXaP8B72+OgFfxVhXgKpYgdXtp49Oa4Cm
xN6Sr5n6z/PNXSrQLLJvZSenxbcDwQOElpOg9+63IBrA/JqWqj+mDc9sbNiF
pyA2x6OL4EXTgnqOCEFZT7cDS4NRq0DXHNKExNQVUT6+eS5XS3MieRii2oio
D2hMM5g6zqodO9h7ntHMZQyRSpMzgVYLV4/Uvy72cItgvMPhaulcQCZXRPmS
vLZFDz3kK8+Jased85lFQ7VOCSQyv1k5JAQu4a34eaT3HZHrOde0h8n3T1bS
httk4MO1IkvJaFaqs7eTvARtQrYr5mARi1+ITOVmWjCzb3C/Y8OM7j4UkJIA
1uxa8kmNiUJjgqaKRTxfpoYZWCOgany8eKHUlyIyyGwqgZMRzJr/snlc5ISX
uOVijC9vwnkFO8RyhGFIMWP6L9jQDwW6p8ypiBtcEXSRqsVMwfdOuHox9iEa
KEzXgUD0EUoVnLUF8qc6fcmLDssWObOcpZQhAdHqQFcL+StMLyvNAU2JlXS7
jx8bLN3cc+7KTNa7do6ShWnvC8s2T54aAd6shsvV3R0nZ4fYrSEElttAyK3J
8SwRKCneX1Gj9XUoG20Bo02xk3J1KqAvckdkPkv7be6uQLPSygDMUX6iF4QV
1vI30EO1wY8HwIusn2HeCT3mjwevBZuYOmeNG2YTclt88lgL3qprUuAA+Fbb
7T5rq315ssGRww9Bi2a3rcPgxHaQmE7kZ7BhMrrBJi5r5CxQTGjijtsAErqE
/190DlSn9EtHvacOTovApYGd3S9zIVQdNYGBsM5QyS1GmLX8djRI2cV/M8Fp
mOWmLLv3mzGyw262BqA7tARltKzdHm18BwNUkuC/SIdmgmQSfZd9/CW75GC0
0vuB2h9dxYZfTTVj2axxAjWGLI86aFihhxWIUgeqF7FqhBDdadxLnWCXAIBW
Ioalb/c4i463I4G71RvhpcNTqBw6D2pIjGAIQ4L4O5vwePLW6OZcnUpB89OU
r0r7ESu+NzGML/ZnOKVw4w+WgL3KxlTZVnKFXemUxrVTJTOarWgOMqroGOUG
1iPatwRw6jgydwxnta7cuvpscnzhmUUfRqtP9P8Aq5ATbAHb9oile5ZEorm9
pNTLFIcyz8Lzfmn6vz7xKCmrJUO3faHdrzHSuOfI9CgpuD+Jd02mv0yvjack
QAhQtWmyQQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzdDRn8pNKRF2MrNyBOWhO0eMi5PMFtSmkR34QP+ht2XhMuNFmcea9M7A/SV2eudVAp2XazJzYtXGch3voGNhPMlQn67i9GaXNteoVJG1D9ecKFVikFaZhF+VvBWz6HLKmhP2ZLgvEsltCJ1z5RFU5qqggm0Ut7GWkyKuEE94+YdNCpVvFYuuYtsyhJ10yYtSpfDsaMmB7U3gGMknW4OG4x+bSeWCvzSCOScTmDHQNa/P9hd3i++GYjTsRxRuyp4+XTg0GjCpI2hiQs6CEH9SUI2ObWJipsMRQp5uUwDeq12fZqFoRFmSbZEFPjjkQpMkHuD5Wxjs73umMSvCevmOagSM1qfP0Dqqg1sCJt+p7o1oivpeCgob/f4TgaTClrtTTN0j/T+zUQ7Vzol9ChKUuEHDZrysxVD2hW001WdOhmIhLbf8aQtk2kvvPsQPCV1GV8sg9hetzJNL6Irfi+W80J+fvB4KE67TLWW/qixIkgJzZPu16WC7FBoVXjiak7HBnhi8WZiFQLFeuvYcis2I3SFCyjyx9+/ZeNXhiysgmHvDBm47XmL18a3dxhhtFlziN9FP7PoIvfKqUQOypt9SXc1kbIg64LicGvv1AoIQvBMbvb2msWPhKAz5SgXq5Gux7rK6d1S/s7vHsXgFhUBJtNJsZ2xBs6vr7l71RuprxALpRIBQ3CmEh8MIi6Smbqy0PZHTFaoHXIwyuDByfecV+d+1Vtc9PC3i7WeAjGBDmyAzRIdrpHDWYOpa/Nca8IvFdH0yzxCoOBqzc6Li4nzUD+i"
`endif