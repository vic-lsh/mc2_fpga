// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZtYP2RO2g1oO+8+Qe4tNHQRdjXcpZ+jlrBUq2mScamy7Yc8p8lcqN7SoCUP3
OhjPGIwIoH4jJh9IM9K/4YUmD8psemd2nsZxOxmX/baD0DPzw/cLOb2u6hCh
ZJt3VV8m8JRRn25bYMPlGoiwSl+AyRez3HhkUVy/NSnpFfAXFYSe9Fg4IYU2
DxCNQMlBnoShwizCe23cey1irGsZoSrkaBVMV9yrY5Hc+LtZvuNII01t7ftH
eQo528t9VaeJCQHfVmf7o7D/B9unF3INNtY2CMXZreLpYfE51Pz+xSZKgRhF
ytFITjx/VT7NYnHx3x4oZ66mi1p/kQX3+LJFxJ3gaA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OUhcFRcfYgXEGKWVUiDLRIQVHekhO7lgiVQnKZyRSXS3VMaqyJU7RPT9NpZW
3l8H+b86yZs7DrjBLTzxNVCmjWHHitTVsDLY14n1mfAZyL6+apf3DWKqS0VL
Wj9wu3xKXd3zl7NYwXsZk03HEIkV+SNwP9rikgkelQLO0yWEz7O8jxrz9Hwq
CeeSfrME3z+ceWcuwqhJeeqVKUFhzEfnvGiU7K5Ru+Huo91YQOPCq9hKuFhJ
Ax/2WK5Bmak0Z1Udii6txkrWchuEUqGzoz20h2+aqW7u5xfAK8/Q78YU5FcA
6rdMVhn6LC9nAG+vx+vtfyNyP+H8ZmqeF6wG/+E4Aw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PLr/s1sAnUvx0ntFL5/w1X+m3Fr98XayrMMcM+i6pbfee/tI0PkUUtb84W4D
jHQxOiDwWoJ00KYhQtGLv1y03OnsrfpLCGuLr3077ocK2muuqvZQ9zw/Wtog
vFpbbK506msTld0pifFxM0F1XxuliLOux75jKrCSA4wAEIeTa9Z3ce38pmr3
SoYHJQSmBq1QkWvfe5oTNHOFvpscNX8TGdrzI3AQFvokPION667kZ6fVROnV
8Oz0GRq+IjpigfY7qntkIapiT8E+CUshm4g6dSo+SknPmMYmOieKNbxEv9g7
PT0zZtaUAhAe6Q0k1w+LcqXS+j1SRTqJZ9XRM21spg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mYSK7TLEF1FvINnhbidZHQnCMWCg+A1frhktXmCW11EfWhnkyWEUxRsS2TEO
yRrCy5Rp2B/muk6PlYtfA1ruP+clkpn9bkyRx+bFMzWdcl8s3t9urQSnyPw0
W9gV4v0QlPoAq7rfLjcEh82e0MpmaA9wz7MYEcdTHOpnQzccVkcwjhyVzytH
FhtxHp2q27SZj0ZaCzD5XKVRDy7y+hUuWQv2yZD2kA83R4QFJwtkUCSJ12gu
pthA3EqW5Lstb6oIVEhlH0H1VQw236lrIoylBtf/YnGVnFmwBOqMueCg2A7z
nG8CxeUnDs7i2LvI2zvfHd23OkMD5SB31BQXRt3ORA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
d5hgr75aCWJEyJPgcVI4Ji+772pI200tOWYEYxf61IVTVEoTgLiM3O//kphA
gjYis5w3v2BKryKLWjn4vJRQwWl4PS/lvo9CPe5iNgEF/ABRd+mZV8aoNSTl
28PoGHkHq9fNCCT1r3qBDEn0/YvwGNX3aeo2YXAbMeV1GuaP8jM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
rYRLpsso1TOqpm6qwI0+bH7uZv6nERoE1nbSlRr7wgdTIaloshlp6g8xZ26l
B+G7dHLpoZe8v9kKQAj3m0QyTlmk/erqXBPwY0snctiPYXoL8vy9Kb9sKM28
8MUX8/08TmCfENykS16+X11EerObb5abzwgv9J9ZDxIXCrYO7Fr4xJSFvFNh
KdI56fe38ifPCwMwKfcH+6MBHn5G5eINFzew83YTXJFqMuJ+l3u7gefRwg5M
awsmXnZMAWmstdWBJ+Gh3JvBv4CpwPCMWVHf/UrhjEU9MTYqrX4eNqrfnCKY
Q9fOW8JvKs298LkY8WSZaqwXeDa1s/Slvaf6Y+i9HM6A/h7BMjj1P9saVhgo
kUcUMu/wMhEPB1v37NiQIoZZNkXJYyKKshkkoDAcuUmHFwJtosAAPPR83OU9
6xil2rqT2y+LVWC39LXwzj754GMpyxE/CHCIVLbxnztgl7vsN0Jt1tQ2loAi
dcO/SjjdpxfBPI9zKlP21ztL2iF1W89U


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
S0P2DV6HuUXTRc+1XRVgmnfL4/v2f8eiTC1od7bVSVtBOkga/OgOqXeMrfXf
rpJnkDQJPzAUVEJnzWhYbj5ss+6q9jO0qhM9kji207wwGjTxjXi/+hWeoN63
ZoBHmiNM9yUi3txf5qWVHkNtkvVNugq7e9NDWWgiYYDAU+4OjY0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Zh371G5ny6n4dL5TllKa8Jz+cNM2J7moJzcoMwyO/tCtLGRzzhFGkb1dX/AI
MjcNXlbFk9Jwh6fJmoFy9+lKetuQ43gIpEUnPb5g17NCMPVb/splbS0NqDaF
TduHcdPzUHn5XRajVq7cfhcOXCGiqyj6L5iV35jBBrxd2oo3/h0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1376)
`pragma protect data_block
HsQ97yHVWoYxC3lBiFBoZ2B/rj1Ir9+8v/05PlEhQhSEgcdg2V8zpI4MHLkS
pAHOxH+WaS/uqgAyvUNCYU+nCY7uBljaO8L5usaJCXGAbW4kqF/5yvT+uBLd
qF9PFpDsP6dFDi290wyk7ankldS8SAKmbi/t7fPNnwaFnisA7E1yH1WWwxGq
5ybPNB98MyNmBvfpNsiC/iOBywOleXDizgEzuEZDQj15ZoZEi1qKiHL437Sq
7n2Cg0pA6lkA0TpO1aEm6HtZr+fwf2dzVmh7waRHVMFmBj3dVj05kxWfzcGf
uELibNtHhryqz4YgTgKLCUF4FXPCDJyF7r5/aQLtiAiMcqXx/GIVM0RTYv4d
RdSXTJSuaZ9lAfvEaxGMTvuoOoC7WkQy1JqilRGEMHhMnFosYeZKj2itpoSa
qbQ/fqNQ5ul0Ipu/Qyy7fMxLnKlfnWS6RjJsYG5Oto+1m5VnY3DWg99ocsOf
4gzh2QhpYwWi9UyB/9j7PMtE7XTe18qmqKs5hDGf4HUZGw+Zxfe5xqzRXwE2
5PAGoXMVgsDAzfHxiVmmEUfD/sD2QuAzo+dKMLR6BeuGiphnc0A4Hy+b3YrH
Q+KiIuiv3Oj42BE2u/KGqvOMC3z7RuilXhyAwz9KPvcNdT+aVYODE7Q0Kexc
XFHLJzV0DtSN2uoLvdU+R9CPDf6sfYmkFZhBjgVN5m9bVrp52lvXKPZAao31
FZOz/5WeAHGB2VHQGMeC/GkIrGBaBexZe6HQ5/jFxW4vJNJom62hABSYRH9u
qlhadEDU3G7gd2Dr0w+FM7NLVeXPiVk6vPPX6Ro4jgn0Nj/hrslK2HUIY3iW
h75JQGRr3o1NTOsZ/6clR/2epSoCQ/Xn8HGLjiHh4ujTtlBsbvlu3RzAeWJV
y4IExPK3I1ouVJzkzzkyBJ2SDatJ9XXo5tSlzlCj+kNlwn/abu+ZeugwIIk3
OnY985LWFh28WGgriMw8ncNQcqkYd0FjfDxUiNOCj4YTB5ybESu30pIgr9BU
FqmreLsOn93TUJaEOUN8yUJ7MV/xLpY85zCb/oUeSsVHx6tMI/JZpLbFg+rN
HgvPCRvGeWsEZN4CfvZyShkCqkuCnWlpkOlZTs93JxOej3BMb3pWt5kz8JmP
8mMEUEdH6XOQl80191kLZwTkjDXGlxU8dpe11O3ajvaxjoO5FMgNQYxPM+n5
aYXEeXjUMdxPEOONu1sEkKiRKKGfaF15YyO9G1pUSUrZNM/+q2/Ly70FBLsq
gHpY0BF0/xuOy6S5wgqoATKwthGGCKZsJSEwz8T5zPOrpbQLktCvu1BDKuGj
EE0+vgG9IzLRcdg4jZDJJQR648WBuffono7q46pjzgt4dO1zjsi3SMtVtSks
xzms8dI7ROHW8lhr9boLSXGEj7OQ/A4L4h4fFtUXwlZdpxN/npt5JTj3d0Qx
F4I4z4objhRNxyczXLnEYdcWMGpJDx5EFaRq7voT801aSnJ9AX+6wrtC6qmO
VBDRvSM+TFa1jOj3nmctB3Z1rm0MM1E1zSdx9CiPMDjdsb/2gGcNqEBL5dAZ
m4xG1LczfFn2bhybNuek6cdjJke7U7rblUhJhga9QlzjXvbTDMu+WUsA3BLJ
c1nDnxWZISsSZmlWiP6Gf6qfveWXUiS6rJT1yoBvSty5ENq8I5brwi0rMqNl
aTtTFqSMfydgaziVzIhtaGmujn/QpuyJGGI6VQfhMtbPObd9jrOO4Nizzkye
dL0ma3UEsR97VzLiI9k79+6EGHFzcVfcZtlnBmv5XGf7HFs+1z312EYceTA+
v1z1fdn6/FYPlQnkKz96jgiKm9ndYZlrkak=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qTf28Y+2FKN5dDsjFP+HTawQQhrhZlBf/1KlAcZs1wEeNX+mdVhOOtBtX9NSmNpqPbSngFKy9C8icW+p1xKAbDMobs7hwDrwyBTfLpMHKigH3y4BZBpzWDZ/tF3WMK5Dmp3Rd1ZdBP09RqrK/3YMjTrsDggPRRhEoTz+a/ghNk66zuwVYF1VplJK3vkgXvgfG9mPMnvBPRVVo78zEDTKhOcuk7SL+QVbxnvvZeXKRamOIpnJWn+Izo0V/7vbkczhDvHG/sWj/y0yHWEJlHxyzV1B2w9HwVKc5cGZtJ7UqPfhmJxHfllI5T37Dd8N1WXRK5Vq203NJUHwoH/kvIaWYE0Emj+LMVKYnG4pr0Fal9kDo00Ppwg5I4AsYnUaRJXE6kLpJs4Ek6F4Zt3N0NNA/bTWMcFUvr2nQvpfa+joNLneja5/lsEaALHpd2CdhEcTMWDIXL34kMBeRYz9UItV29Zpjel+Bht7dRTonb5Pm5cQBnOwX/Pm+eMS815eTp5fIeKZggBRprFwHNl6pliEA6saF3VkrBemlgguG0jMfjpIpnpjw+T47FVd7FGQ3heuvXGypKGQlztzknq1Pe7242n9qUVqkay3NVOXgSdYdyD65A3yMNVyRN+USj0FAxrtH5De3tuGhkL7aWldsP9pb6Rlf4XuwD9M3Xzb+7rV3VGRZ58b6VlNSBl7W/nNwMBT7UsltQrf5CH9aDOASl+ZQJV1MTK6JwGGFPmdLe+5kBCoRKTflg1PbEl0oiwT96BtVjvrNexPceqsIq/5m64iFvg"
`endif