// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pcft0kWiXq06Xl2+7CtOcXSge9NZ/EokorgXLMx8VMYJN6apkN/cjiS0wt7J
rVlFKsFZG1r56Wj43Eq1LnsZwDOL25MUf+bTpENX6H4abjN9Ncagc9f2NNiH
LUiYSk1BwroR+AgkhQ+z69TNH3TQzcqLjIXEvl9i5DAsISjRsvchDg/aULXx
fGef+vBIr66ZsveRALOLp3bYtA/7SbYP2uyRKgaJUGPpiAd941XhKk3/LI2B
GVd38Hct7fvZXu/DnxyaNUYJKEanzYhW62aGi2iHfESXWVEJvz/ypeJPF7x8
x6DUz8j6uXo1KkR5kQ+TBq1BaP5iUDgMGoD+MpwWcQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PHVWl2pjNdZyV1jCAcotYQfCvsLMqKiflorAB1CcKPskhmBGAsIVsZrmL2V6
bxcL3QcPLsX5xy7v9/xNSioUTXInSK3Q2O7XhS//OqYh4mNuwV/FEqqMXKkn
s80Tt8fYqFLrICXVkeeFb3sqm4ZJip8rqe1984ZiPEYRbD7uFpOxT39guQ+n
4ep3AghrMIofGpstElT+EF4U4SGXbVWVlRV20sDnkB4AnZ/Tr/8ohEPmdFcf
YSSbglo0lG/Ej7ePRidb+ogIqfARfgKUSZFAidkq2chZz6zpZJab/kVwgVmg
EK+EiERnyL7WesdhiD6Shn4W9UCghBpAK4E+H2GFwQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JoXFlNiqyIeek1+t5Yl8Yv8Fx4kjse4QlKnE4hNWO2xlIcoj9Xzh1gP4rMtN
Hi0y5Gxa552O4JAHFdyW0jc35qggX+cKuZyC7V1GXJhSlXn7yNpWSX1GKzV7
o4YKO6o2GXzN86zSBnyrBFJWQg8yWeKvApTU02tezymEql28MaRssYzr3GZK
uvq1uMZzR9m97NZ0B82S+UqjvEflU6OaxM6klhlw/gcOOuMoxn6a50DGFdik
aBOPYPkwFq9tl3wI9RPrOMb/OqyxxILKETHrqWwNBmaNudF/pzaFsfbobIJb
DUE/kOz8E5oK+6vC0xDMBr7ICmUDjga6Glgr4IOKEA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dy4EOR4o16veCqMFfDYioXq/ueELfM8rvC4WYVPSWFlPLOc+zg1fP1Rs3rh0
M4EBBh6AsZd3a/xDZ+kOo35C0PMBS5SSYZzmEOx31r+cCKpHGNV+TiOK41q0
CiksckIrp/ZY7CWXZosZA+p9muGtUHU2NUrlWCpsSjMqLH6agaYRipd4wcL4
xo33T3Tff5l21pH6mQLu/lT9N1T8zXruAtvfY0B+tqxgCJFiS9ExkOWV5h8b
d4Q2M8FZi5+illdnCtPZ7UBMW0oJznKcoaKQrAYdqcayyD92PBE7pxTtbdq+
Eq9xvAfHoOjIlehZiUaO3fCXb3CJpkD9rovo2bSnwg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jdEgDEsI62bXJxLgVKqZ0xuUdJmb6i+3N6KA68lbbEQjfIo5ydHA84w8cDiO
t8aOTJXp7GHSs8K0CUI+IBu2pM529mqBV+CLctR2BQnL3gsVX+ezmEitmxIp
92hkEL2rBtRY5KkLyrBlL7BqHuSlaxwQaCzAxpp6OLTpJwjy050=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
uD9oJfAGQm2KwQGY6Jgf/6SUHlWXSSU6TV0lTcWlvvTCto8znPlUnqfHVPRX
WqWpmgiEG5poSCHZVYirGTe75V4LQ/gouSWK+2M84CZ/+oHhQi9y68xB4qKr
q1jfW03hxkffwHdkiSwk2WsNR8VnPTQBTVDlC0sIdCnbbFpJng+TzcA8Og98
Nki/dOHpZqQwBYoeba1DcfjZEQhycg422mIDX/9vJEtPvzTSKzSiUkgU4/E7
EsK4eWSRwj3Y4L1qC31Bg2/Xa7Cn8Jzh8Nv0kcXNAeTIa7lPLIpqcko4UoW2
kW+wGmqu3THZccXaBkT+sz6rmGT0Kz130VQ9GqdDPIhxkqs7uANYcUzLG0Fx
fD7i6dj30PN32wIsVz1TnOVrgvTKRqCnNnhYaIFd0DVTaufFR6eXSIwaKtVi
Hrs0Vyqfq4xnEYtThO15xL9Eod8wCKiuwc9EUqkjAg8EIFH/iMAzkdTkMPtQ
MxokQbmWQLEj1uL8FqOQVWX85gBjP0lt


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IzmuUNMqVWdXcKZZ2iR6HOvVHCYuHwxrPxNsIcHugzINYshnmbspkhy2t5M1
iFUzXTS21yy2HFa0Upkg7MGvmhptfsFTl6Vynes0YIolKPOHNYivCvUxv9Su
6d2Uofe4qoUoXf0Ut2six9fw42W7liwj0s7cWFkAcPsZUtZbIpE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RIvFaBzmQF6rjXC5EgWfrTDikVtD3BS/2dt805bIP6sTKWXErXlzixYud1uL
9rLHpBc+832uOqQQRTPlSOegOazggcLAz4Q6jU0Iljxf56Omi+0i/wJ+SUqC
6eV2CylCjToNYdBi+kAs+/E35mWlXirdau23TTdLScuhiBZq85E=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1008)
`pragma protect data_block
Jm70f9hnIIoTSu3wruKxriiFx+9A/q76KFnIEsW2T3uBfDgX9eqhf1l5ZIec
SMl+5uQ3gcronuQFM03OoI+UMz4ceRhY8s0vGPM8zF1NdF9Uk6wGvcpT2nU3
aqAAfJEoVUKQMS3MidryXZ4PTLhmF6lm2hT16e/sDn/H3Cz5Qj+FzPadH8KH
wzVpKsq389nJRuTLPqHdAvuP3cHKpFEvq5sokKKcjk26aWw79nPsIbbezkVy
SZ5v1f/N3DKKnokRo6qqgK3fyEOcR+1fQTXKqAPF3Y9QO0CK1rE+pUfLsF84
NYYV6sZepr+lhcWn5XEHuXLASOXTYEVLT8Edo77VHgw+BrAv1dMqiMQYBOwv
QTegweDsPXiTv0Cm+WCXrELpOUDzGK+z26/tim6jGrcp9WaqHAOTcJTY1dtg
dbLC3qXC+MrUW37GIAvCFZKe9DRWTJD0FhbufWNKxQq0Rq7BK5/5qlr4ZY4B
5cPiBnoSS/PLZw+TYJUrVvTBEyBOgHhaHy99pXRLZy2chMVXb/FClOFpD1eU
pqQtxdf0jwsz731Z3A0XsSZQksZKe1LDsA0Z++3XgSb++rMxSgjX9XbDod8C
qrEVfO8ix5IB8iTkvcGP336rvVVmVCG33NdSPeFasFD1D30R1YiyhJPmLc6P
bjOjj51h/wfmuTQKMcqGeRuxWDlZg5tSS+MvhDiAagF4IyYwRNRKCHdheN4S
Im5xmlzjpvWwiIKGK9XhV7w7ol0idyeugMYqt2dpPE4Njp3eSLppgoNdycAG
wcSmoKr97gLLL7E0m8zIKPfqC4vUfmYmZEtuEj+x/4e0sap7Dnj+VVaEGve7
L9q0inAvbwoaNt7Uiy7nA7MDyA6fbuy08U2Ik30tw/m9Jy1Aui6RQnGquebU
SoHcE912rg/S928/5GTriQ9EcVCVkYPAxCcH96706LFkUmmQCEeqk9DgKYxp
3OjjTF9C6pB4XNzKVK9cQAnpE6SmM2QnczfL5ZcR4q3ZAxIP0pkS75EcJEhT
EYCL4EX9BDxsQj2nzBbC32p0/a1oQjYLECm8kCkPVfiZvZqKXuUBjawsJ2+M
1hcYH9kuQ7cmza1i/ce9tRQh936FvrNNVvZDFCNZfCRfT3KXXDwMCKUBvxQI
q9ray1pkVPjVKZBYWwJdSZWEIh+aqn9RLVy7SRiV2u3Kd0BOD1smZD+/wNjI
80jpW4BD/zH4nrtWdiep9p8xnN0hNTtUmJxkxsVrxnWwmFoGByHcT+vYdJpi
aMEKRQZAYLuTvvmKLUlqwzl9BT4EvQo7j7KDO+eH+dq+/gYd0Ikf732DY7fn
Q0JY7gzyN1osZwDDXPSHB/gA

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqc2e729KDVzZz5LSiX2qLZaS3UV+B/x2R1w3m25k9rBjUL7qc9IauDo249dXyeExnfmqtlWzvmd9pWiwP/1I1Oaxdbj/BF071ny3NnB8TDrGe7wXUQG5sdCzKTxpcbKe+Bk7Anrdk4SlwqVzqV2qeNIKlPCwW35ulldCkWDTTGuI6JxlZijgQCFDvgltOss0RCSt16PhV75Q4B4hP3IIhi794/wdHOpu/tEbtnIYEjiW8699el0lqo90pePoc6+0g6CyVuaA8NAPUiHBSgFeybOCCSOa0PgFTUuhchvYk++4O6HGOA0qAKpC1pCvizfyNOoiBiAOXEoORNzeLEIckhSjW/BdWQZ4j1Vx/H9EHsGRk5qXPFmJoeDLX8y/Ea1KNArt62ZBCcbpztc9fE2gdPgh3Wvv+jQPP2THAJFXIqqiXqnNT76Sd1QbBcrZoQo+buQYB03YJvzWIQMTW4FwtaOCjkIeRVF3Ieow7kWJAqchyWH0umTB8l1umit2KNGU29/ZspbOvlORaxMNxLCgc8jIP41AddT12+v52EcFjciNSSop89bGziM1NvUBI6ygDAVyvQe9bwc5JibVWrahgjCe77mmnWsoXUQMkH0pLZQmFDl+VbJjWK+S9wrqkdgvwxJtZI7qU+2gyd1mPfocujZTqoE+7jpWvEB4btFGjBFZCLGsyb+O0Akas8Gmp3vQx39GLiv6D68z2OYvoDUoAO4zvxRAyLq/UtxvBBx69hSUbmlxG3CHlDTgKlh8RoZRWFhQ1QSRTL2c+KvKYvw8czV"
`endif