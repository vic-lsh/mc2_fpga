// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
1UAJEL/LZtE8l8arRALDzmCOvBwRBIgN7NZwZ1X28ZBCDMFLUsPTeQx477dp
PWkhWsKdHswpHYmPN2psau3Uts8YpvsGunFK8U0MrWyyNPXdvgZwpnQf5dEO
wdM3Hc6dXPjBu+W7s3En15nmEoMP+1oXnXxjFzyd3oV+u7NP2IQykchVvdJB
m4+rkvcz+tpp7H/eCvdn4couwmrh3reEnlWcfJNLg7zCAm8KYc3CnJ7TJDVX
AHZ7HQEYpeV0x2j35NstYhEFK2qAxowyBGaRQ+y4T/n93D+qWuaeGBkhfZFi
mPUfa/molMzX046Ckgdz2hBNsLJ9ksMzA5hz2ZCJBA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jO80M+IQi9Br5JiQUzoCFzoDWIZ5Wl1A3Lusl6zKq0E8fDe0OYVnIuRPx7/c
bW8fl2U7u3onGAlzDqRWu/PK4kHYJYpSluxHQ4wNK2SqxGAdsbIiF+vD8lzT
gLNantw+MbLpEEfqmApszh6wwDh7x2jPCH5eZlJHgqHOorkYmd6GKBQhZtkC
RFXWDO2bx6TvnSS3EFWuF9+Mwfrws5vNs9nNQElbqtqdEB996zU8OuKRgbUo
EjziJWiOPS7y5IbaGCB649oRjc0GHCI7Tbvw2+MvlZTnh3foyQ1/AyxoMkoy
JLsSn9SV9Upk7u6v/O5s50i7NWSFNhN68wik2R30wg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ti3nEqze0f6N4iMJuwJurJrumWrZyuowrXf3zotcVRS5e5PInGhaHESZIUyI
BkeBnQhloDFtP/sFnPQKVKLt8zdk8VbHlZ/1Dax0PNCpG++zk9AI7jKqFZ4/
uaNOCeix7ezUz9M4cO8hHw7g+1yxV2Pqr1OjZZtD8canj3Eb8p2UVzkIFuw3
pANxnzRIqD3aCpxo5c8Rsowr0je9G0tY1HPNkC+Ky5lfTiTUob/ICPr+tNwS
NrtqCOengHicjMQT6emK1287idgujSB4I2emkPe/3UUT1oub3ukSCLexh8PA
RmCR+bd9VRIfAvJnuEH2PlMdeP4OyXMUSAv7G2Xkxw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jQJXiHz6dD9wbyP5jd8Cj4e0U/Yt+UPsvrnVuf+0paYCK5GLDZX9G0PW/BfA
LSy1oAiEjNj/onNyF57cVLP2Vy7MXe6ltwi9MaY61rOIaJ+j6KtfIpzBc1Qm
ezClIrylZK1YNJn0y92c+CBGeJufewsqiIPqiU55US5BJgb5EulmWJIm/sVR
s3n+bbxA7fxiQRMtcSBF8dfEN7ET3IJ8di5vMkWSMNcuMGafHFds+BnL1umy
1CbTPAJtUl+cZ0Q54+tkEcE4lAhH4lpi30nKSOP71iEwSWKQJD0yq7X69haY
kebI30RVHiR2j+2FvfTa/LrPTOB/wPoQG/Z0AMfMwA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
raPpJNZ+SgcOkc7KCHoQbJHg7zVAHeVL5JITTQRCOE0wJFtypICMgu2soOcS
yQaNa4Hm1YSlawMjcwaNE5fAPRTXgk8/t2m1RLzTEhOa0NlQIJyJkvzZ60zF
s76x+YsjYjuziG8Q68HmvKHRcHKDZqaF61gWU5KOwyeJzzJKKr8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
YjvjQEEstJ5kruMXhr8EYc0Q/apR8+pMInuI1bfONrTej/GL2Qh+CIEMVqgC
JCtm79EjHFnGgmtKRNiv3lwX+KBKKGiWLFP5AASKLemcOWbiD30j8T9kqZHX
TV1KOcdZYfK99lXeIZHUvefyMDFYXy8kyVg0zolfA8Koy+PLfAflzSIs1Op3
eP1FmuPdTcUm5uLVJ38wHTvWW68ZM7g6KZZ4jDXWW80Xt/YMI0mgh+cgzFzJ
8yE2TqKyRgzJTKvKeps23i8Id5qNmI0U3LNuY1LU/QleNnsmLxIo5P6R+N1b
111V0aIBsw8tBr9JGb7UNRCE2enbDNuhaCDma56cVUVx3d5A6ODi/dPT9CF3
aJi+segTZ3oxiEV6qrVaHsI3TynTA+kfYKYSLiYfZkgWVEWTjn/Gm6nzZutv
6rboV7+qvt9xNNs0BsgLjCYDSiUtOrrJJlbbGY5i2GfkwyuPVO8Zg2INK8yG
lfxkyaENXpgPhw6T2X+GwL4b+aqLPqsb


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
H63X/W5kyyX4I54R978UWbpSbn4Zh9Jllux8s16vD6MK9OYoI+hkCZ69LTkt
wzQkuyBtxnooIDrQX6rICRqbIkUGk14BtbHsFwS4GcpBFxdqU9/xBcRL6ABN
V4SNNTF8VOlg8gZOBosViqS18k9+Rq1Sm5VmntMxgx+jqb+8vJk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dqqG02SFDWNkZrLZeBpiH2Ec4goAknX6ybKSnyG+yA1PHTppPuLb1DS5HE/Z
4r4H4Drc6UCj7Uk8qjH+Q42V7Rs7c2nGBJhe6tW9pjaGvUhCsPknuPzeMA/6
uAwoqkC/XmXIpHeW8lrrrva5GDiBskaDaIhoWHFJ8ql618ZzsH8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8544)
`pragma protect data_block
BvwcyzVDM2H4CVRj6H/nsL97ALe0fIfSN9w0WMSslzNHMSnlS+p09JLmbP37
nKuk/pji5tAMg+PMB25pLL6f7WfYpwfVCz0Y6bOVaiizIWBeK3JOw3elHHbT
y+93ewz8w0e1PPdueLk72ObCZQdLrcDQzWjGGDtergL0711GNpOPY2HSjR6B
lfof7U9Yv88wFYdqz+LHL4NBnhXzi9MenDvJ30iT5y8ApMqNf+bgMpHRFLOr
F1vtXQ7Y8C2jNVN5wsWzhN+Vm55TOy5WnOhLBEjTExumsbAfAIgOl9WeprbI
XPUgqeMfzSuLmzlw2S006U3YqOB7rDhsX134DiUNgsMQT7lSIWPIpqrjN+eN
xHvROAMRJ1dWqDyCKPfNQ3BlAR7xpMBz/3j/7kaaVKsnR1BUaUxvZbtYI1q9
LiY9io+Eiw11Jav2+28hauMZ5zv72w9i2xEnS0WNeNRHS1MRNcUWmEmapR5B
L3BcUra0l+hmAQObiMVelUMFlDGLZQw7OB6M+vUMY1QusBs3GD5J7pinh+vL
w5tNO3yLE339fTvgeukve0mZydqecofy/rfIRXDQmaWC8EfsC7V3kF5c7dOq
Pdq2XDHXpNfTL29qFRGO3gab2Eb85YYBNVeHJqgxAbgVxmswohA/9PRcorNX
khx9iwVp4jMClPR3kZ5cDfH5ER23QKfcVRw4To4DjjpEap1SKhSqaBdvH1Pj
V76Uwp5jG+jg003Ekp2is4ZCn0GukBvZZkIfpGPdZt/Pi1fAFwL7WIwa1aCU
XweB1hSEvA6MJ87iscHcd/pUOfpqd3Eamon3eOfDTAPSE6U/fomc9ZLJI/KN
TCaskHzaAMRtLKGZ1Ym7CpGiqCsROY1LD1CqVvOaWrEtwQz9yeU9qXX2BTPz
s20p8JH4DeeFh38T0UF+YU9+rSn0I/LmqTpCFw1sB9nvXU9p/UI44pP0hR1r
Dgky52+ZzrggdV8VqhbDzJkLamBSUz8l/Q08t4XYmZkykMWmHU1phvJ/3RjR
HU9gcWJn/xltykNKhAymeULQQNy6m4Z5twjY/zD/W+ilzwdhk9XDL3E8WHrJ
QpZDy2XljPitU8rL6OWtwp7CQ5bqzgz/CE5aLxFxRa3YFwuLRRWrtrj+FJ7x
lFcM2UMEpguX7SNbvx/VCFRZH7V2ufONXbBzuof+ovkaPCWnPKWI701caRYc
A4YNTQS3D+T2SRVLX/o7Qr4nKufhHNfhpA+Yz32ZrXJAMOQXyiUS4VbSczNC
GxDKYmWmUEwD2fC1+5JoNCfnx7kVFy/vzknYmagbaZ5Oh4devOv+jf/KH7B0
/EgpbbJ2WWXXivgedbQhhPmYfFdfhKkK+yw5KWfBnM50e+s1m3Zm5y2VBz79
7NEcFJJZVkL6opyvgGl64k0nb2bb75AJhRg5d+Q4+5LV+kmTd9B+4PvY4Gig
KgoJyKaWBdUIA1YBXRAAZggB6Ij6El5pI70YD67ALWjqv7mUWsZH4EcoFiJM
+iSRZokzpe46WQAKZvcx2CJW6W9UGLq5pZaXiSwy53QG2rxYcEIOY6EilUlX
454P8A7ghAGp0I/EM6PYFCTQbMwHJuN8+3juNZbAS53Y+YXs0tWamfi2Wqme
8h2BTFAaOuMoUW2yX0su9fzL3OH/NspUPsTitSnQme6pUCmUXS7wVY+4cxBN
LPmDe+wquYEFIgfhO5+AFggx3kFdjd63j73wgjX7Chxgd3yd0iZub0PK0w2l
u3GJXvCmPxcirBQ31UbxzAqHXlGZy4bWQigjZCL7vLxO1LtxM+MkfHmGq4IF
r2TSrvTEDWRN4QQdu1MFSCO7+h6Q26JQxciqzsIrVzt4PniFG/lGrvdov9kU
GJE6brJeMh/9Jzy96Y/vHKhQo/JEponHEd6y++e9lb7jt5MFoQn08wvkbZ9y
KYG7ibPavDfEvu+Xyx8DQgp3V3NZU6lWpyzHFbTQy9qwbPdTIyWsKXY7zP8I
JMBP8kIo83b4Mj/XZrPi3g1DbFLT5FsBBl9kzW6CkrWSockoDQhS8ngBJprg
Sa/QyM0Gh1ZbVG5vR0yl7kvohtr7AESRQsfrL3IZT4aS1gv+TvSUx8WFbgU6
IuiwZ10r737b71S8kVuLrIDRxFt7vWvXJaQdWXVI4lYmNjtKirwZpxfMYTL4
znrGMA/eZm68hGqjo5lGHtB3QuHBpInAuScriRDfWq718RvUtx0RrAbKUsBu
ZVL65UQvoSd0vh2mbu1/cKFsCr7wFIRWeYwf4PSRFx2Dhm4zPZr5vILUWfvc
nu8SVPiLg+TYQ9AUhk+UO6jDRjEtSS3gZkWOqJ3SAGEzDUQIsTQuZZqH3JNG
59GJSm87ASeE5pwWW7w40PD1yxmMExbFxpxNOt0v3EAKGOVBWa/n3tXsRjsd
OObQW1bTvYo739NEpCq3p1tzkHyZEXycacMLAS3Jr9VhKp93CHhYxG20gO8G
f0+LsygAFTMx8yKgt319pQv50Bqg702WDJOhv8nafy2fB0khytFX6B0XEr+J
0RJxsZ2oxS6meM5AatdOgi1W/JDIWWuUXc5oCtSzSQzIxoS7Ph99NRPk41Sh
t/A5NcbfYBGLhXX+ZX8NXcTat7JaKh6k9InLgEPU6mez5OBJuNk6S3MuFgnf
2BdHReMczuzwWAUokCbXiC74FZTWo0UfOZKzRTo8qT6UNVmG4MxWkUqCVaB9
aZnk+7SCa+AW5TA+VA9A03VXIBg/mYprMcV90jGrkB4y3zudPn70Lcd3sLfu
t69/TP8B66FHqXI141bLj677NzeR+zg9Ry0nkRMyrA7oknsWHZO2PvHdiL1o
rhVWpJp47ly7oQA+EN0Qyq3VfY4QVjAYmtlY6m4+85egXBIn6zojZLh4q0uJ
GmtaROM9uHVTDm4eCEn0cP64/5mGycDnltAPM5sZkgxpGpjQKWYnGEzxz/mI
Cex1U7X7bv0lM1HgViDlvirZwcMmgPqWYAaGud+4LQ0f8YNFVH00n7Dr/wR7
akF2Dk3dWL/FbFoXciGB1QmPxYFW8GDVJng0yiVbTkAtfwM6D6M5DTKl1LVt
9KaJeAmyCFjM2UFpKgPX6vsS9VASgYtB24SXm4g4JVSwRDk7cE0P/8x3WFBL
3W1bF6GbaQDZsKDBU8gV9DOWESUIklr1sHgo+dX2YnHcVsA6c3/AQ7vfLu9Z
lAFxJQDn/PB41UwSRlMHOcAM9zMq7VzvmIkPMkknj4LE/ZXkXZpyvXN0I1CK
cxZzaNEUPvEEzD8a42BsWRdmwktRD3Ct9zPYUu2mt7jyR1FuIrtA3B9WhczI
Amu/HLURmD1DaDIsIxWjMyjYWKzIg57mAQWhOPjagn/FpJnQJvQ6lPsmEYjH
y3ohuBTJcu+5r3YwX7Nyp4avVZ50vAlZZwcLqKHLF59CnbB6h26vb7zoBGq6
j46dNOTf/5jqSqGo/cv4u8t7oXSvnBtTcRe4Rk/EB+mkCQk8hdK2hWHbwhAA
MVg6PTFlcucknWAsBPLonTVMTV2MqRKUyK2uc0C1i8lTzE9LG0/pUM+1Zlgg
CnbweNdOo062J2KuD2SvCy62KOJo7Tfq00JleL5KlX7TmCUbtSj/O2oyj5AU
pMD9V37cOLiaAkKISHilrS0rbO+5i/H52WMV0IpARxUzb0ReAhqHyFx/FSzn
aqzI4qp//HLS5d4IzfvwRvGsGcJ6CYez4cYEpKyECszjigXYHrQXdoRSyQ+B
g4+Pzsr6EIgO1QvzWW/h9r5WNBR9myaMObOQ39x1KdWmRQ+U45bX+VXKbtsU
y+KSdicwReUHlN0o04SfyvbQzoE3vq3KMY3nkzmtsCmmIz+RxeW0vVFvyT10
JByJ2Yj61GHOb9H6gXo5y8trnFpFE1xhjxPgjsU7Gukei6CWjJOr9Vb11kV3
FSV0MGLNANxPdOvm8vBTimtCagsGrwcFynDZsGAhTc1Hk2sL8mhvPEylQYCS
umf2Pz+dvULDDp/wI0FEU5IrJ+dcvcID8vYsPQlqrj6Z65GDqPONewtvQ9T8
zn/6lCsYQNrt0H9veQRI6rLpv/sEtw5Et91X/5UkR5RL2tbzgTrB5vzspqwV
+4D65GTjRrh8C5QQ55HlYCiq2Cbac4szcYSC81FOYKMaXTpn/rErfIagbBA6
lt6FrBchkCYqVvB8Xyx1ioIEcHdFFPX213oeg0FxAM7DjMRuvOgOkId0m5fr
bEOsb/FD8HUrIxVZt5GDioiBcYSK6nyHYldaIJg7Bz8fJHiDhfE3vRNQdaf7
e/DwwloAlAN2iqOY0EY1oIlJ7DlTGQckFYrpuDRE5OaZTfYsuYm2dHsQoCoX
XCrZRSBxAPvVwUKiXipAZaHEEGMhEtYcNAouwncYQtfHSTI66vNFwJje8BZl
oeeMaqvTfVQYHG7fuASt03Zf8H4ot/uxZTfJRFHlg/dRd2tE/h8sQIltVvQP
tGvuxo1dYP2ffEsPA1UDNTd4hafU7lFx4z5YVM+cOwyo0Clt3hFuJGN63EI+
g8US1iDuzRx7JCqyYECcbeZIEb+ozweaNRCmuSc2//e9SEa/MaZjw00OT5Ki
Vl7hSvs2jP+ojn6LPTLm5Auh7MSNTbUeftt8a5DFJydEOnHHr4vODPFMmqly
swtC15WaZyvyR2xIG51qOtEUkzZLopajJzIaQUygcH0BgTmerl6pRWb2lhKy
0z/QfYQCpdPN0WDqTwE/KF+YHiVppRHd49ka8lADbtaNMCXv5wcFL25OMED+
FT4qEOXBwSfYKw63HHUxpnMKxgpxZb7vZgJ805XZU8+ZLaHRtk2NPsmJLITQ
kPAS0miCoSUhBNCrISZMhPsu9yl7N1bEcg93XGRqAs9xWHjWVjQj71YLdaXL
0WmrzHTgbXSJ2eNfY738t1oJXujTRGPGlr92PO7bBRyq7HtOPNGDcDHF/m3f
8V9w3V/snZungZwtr9PgyL28ZwKMI5hbqFjYm1pmwJhMznAyNBepQvUqYSKA
0Xmde3dUkcNhAu6WuQrBNwuT2ZEudvlrDS9xdAYqU5K1T1hdP/Nwi11Z/AqW
2dl3AuZ4O84u+IZsWlS9lYojF9jily+HWzsrFhX39H4cAGBUPMmvsCW2jHJ1
quRM8Z2xlfmG+X7irezUizwb4LcvyFbXsXfmBgz8WoBRaHCJhh0LvY8QS8H7
B+g9nWx+DWOUfadzYFKIOT0oPb4YfYCBPQpwvuTDv2AO0RLmaGpDhdULgHGB
fghzlo57Ky2Lw2c3ImqtbZzlyFpjnac24g+WnJ4uFfbeBLS1t+UehYn9El0v
W6je+FqEiWgq3x18CUQ3OOEcf/LGvQuuT8DVJAzA3ya/Z+eBgmckM9Cytyv+
+BOSxL/y6aXx1ypgo3aM/dILyjxmSJbk3izUPIPt5ebGtLi8O7lkiMISAOaU
G7PRe0a49h50SjUZk3fuponyI3X3BZlWlAxqIkVKTrze+hEaIfQMKj70xepK
+SLLnYz7OauTUIO+E3BMLQSUs9YwrFdQ2uBPYigWZuyJw6K+CcNCxMVvGicD
Mh3UPPIjPI4Z9ac68hTET3xfhqcdtO+Ax6vDL2r4JbWSuhyGKlfCIlpx8W/n
KYcRvrc/aFiyBYf6fa53GFqz7ey6gFfd1PTB7F9FiTBf3VT3jdlXQ8BIzUAr
NS3CBUCiw3cRVvZyc5A5JRbhSpRseaXec6IFRzZ9kNzYPdWtRiN5a0Q60eSF
zG3Uo2WMS8Jv4D6ifqeU8vwDu0cmvyb+6rpNMi79zGmhNpcpQt4H+voFS6C/
fv5kDv5pTfIaJofJu3iUdseG1YQIzpONcTHFyPjMbPzZgSdr5oxoAfkJCrqX
oB9iMc6l9oGTuwzsesBoGxt3E1DO53vH2bkx9Kv3OFWmceXzhlghx4x+dZLe
Vf2emH4t0EEVZI3omNCYF4jF6jD3138btQcz22MDlA/9u7IbaGPfIUj6QHO3
lNJgzzDAGOIjuuLl826GVySk1OEtc+d+0/CJDap5u9QGQwJZVG1r9Ptte+4o
PhtXmbCu7gJXELymTr9ezCOnm6a2YbCBT7H4hAYok0IAft1zfLzgnF8ubdkl
Gvq5DdfsKXGCweY0it/jtmQQMSgZJ2B9CvwrGunVgP1WHDbwnjW7Kj0SC3QL
v8Jqa+D7ymmk39+MC2rXn/BYMdjC3oHEQOmcU70twcW4BrD3p6/OJxIMXRuV
8HoM/THdRwg9gm8GHa2eytUQYnMVSSE8Mw7FZRLIkaEPVpb63qQGLILFI6MQ
FH/YMRS6nov70otkhVigKUw6v2dlgn+7gnKm6omVA5gFsvLBowApXrSJVZ4y
1+FnOS3gtQudHf/bAcfRLFi/QQWeW650n5mhXb/1hyFzLqaBPZU+31Pqj1VE
POwom41bIC2TtzYJiO3ZLMM9/hEwDjPll8/5oQZZ3k+6snRJPSXGXL4JNuaz
uU/xFq5+Avea5LILjndhalV6bnKjNj8wWlBsRbORSMV0qt7jU6aMtkmzkGgT
XYAZQwjwrhn9ckUPukHk6dPlQ/3pwpsC+vmfnY/qG468F7NOGdsHMI95NX44
pqboPkoc1m6eCX7nmvj3xK3KVtTfEumKEQqycWxGgbqBZA9Xx1VbFSmOQ/3B
GA2tDmmgRLbTY8zcUG8o/eZQSf1XRMNias6nNP6ORybG248fW/zzX2DDk1lY
VfxJllLGlWVA+OkHpGEfCSS+620lzQEOh3JEx6rmrFGhz40D/UegktHrkUVF
GgQOVtny970xVWFNZMeGcEi5uRgT9Z5Ac2cffdgMS9Cpz5b2HcjQQIu53oJV
9x6qzuxyMWGk1x0Ts/owJsnRtJZhACYC0YXMcmnHwpsDu29x0YoBk4jPPMzx
6HoXWe8Z5yvzj2TFgaaOf65RdEEYdk9vpDkpBdzLPGVNhAOocETJezj19GCr
z6nEFwk1+7QPaF8RTSM22AR8wZgEdj1HqjWnbjD0/O4eCfj8+t8D//KkCuQn
QUOQ/PMmavKoblErND7QF6Nku8LdPPMzK0h0Kd9j9PsrND8L7iYst/t+JXxS
WI1p5AkY3iM/vzH69W8qOj4GFPvykmgz5M1aSinU0VIt/0GYHvJJY/1Dh45E
4ISIB8gbptn9NGc/Zt2Y0mtUruySizBzhRA1gIw5cxloiiq9PFq6z51l1sjh
QYON6h9x+6v1ikuJTepeG3YHV63KrFT/Z8SrDHa8T9m9qHEoo9RNb9SqjCaU
O1Omi58GhHTFg+p2H8FC+BHaR0YEsa1KWBEXeeW6ix3sM1JiFpfVW7Iu3YDu
KcTLNZ5mRL4cSQQEwutd5fidb+V+wsovaIkAgZdiXa8RJFEoRHDEfKBD+/Ey
J28PH6J5jMoKXEQkDyHPc6riD5z+ML/4fZctb7uWizjamIHHYsZDX5PAB1kj
zksrF3HaQqSyt/+vlWVlCYjABoS8YDeD6U4Efe0PmJ3/eYB5m7g0xreRmtgI
7BE0v3JTmtKStMaiIvyVjBiVf8ijgrCyLWPvMqQNAU4udpmJJKG9tIbPcvNH
ayEY5WX8ATXYL0KbduOnDqQriFIhZsF3IsrW4i+km894xuj000SFyy0QDEP3
zOzZVtysiGPSfQt9I2wLm0XO6KkipiPgVxArwtKto6z7zmUxJBpdv7HO9ohT
NLk3fZiaCEoBTidmCbd3sO05gPmF75S+4XkxpwWpJ/mIXZCH9Cmw9ysdv9UL
3Y/9AiT8/wSWhki7JF9xrTC73OgRrN4RlK6g3y5s94IVTisdfyM42RWvuTcT
Wg+hHJSoqO0IP/cHUcZEsODcoHGRcPHsQwGwkxNl4aS0GcAut5DIY4Hdu9JV
01HLmuj2gIijcNZu3V+/OkB5Yt6HNyWDuIt+CVyEGFZiS27vMJERuDZWmXWs
SociRf5iVx2aJ+cGrc5YWQEe85wim2TPyuN+BaeH80yO0krbZ9p5xgQCE6sQ
mctWlYLldnePGyVPImvf2y0IDZ7QpCFLU7qrsCZIlHdQ7WZEP60slpviFnd4
+OeVoJbMyuqw6kYNRsIWnfWp6AwOuY54yqM4Chj7S0xARNFRQFfOerBygu8i
7SRAhoXTwWC95UTf7LaR22EJ2RrAaBU0JpQ6T7u/ZeAC89jdeBvchia2QsT1
MsR/oc4XVdIwp8CIbb9vCNhJVghC60PEuD4/CKOqJGCWIarYW8+wsg+smoau
yb98FgN0gOqGsvcwbXN4ktkImmPPi42U9q7cocoRkA5JpXc4TCzHpwRfJTc0
yO4AREJ8mgdpSyr6J71EddBnSq4XmP7OLg6R9WoIKKPp11V86f9nIr8glmqr
GAtj2v6O1m3wAqOoQhMKkogBYTG1uI1O0THCwbC2RlAsnkZRLrYDReMoMBXy
TDWBmrjV6+rBZ3gz3uKSDYxCPpAO9kRf4tsRam9Ym6Yys4R7C8XzbIAXCD3S
qmXG4nmfeMjhtiXcYBiZKjqtYU1nW1XAWAM2UA5BVqg2jfC37DqZyzMlJbzr
ppn8+FaDCwnVQUX9dtHXnCFef1iPHBEpOUKQOU7rlu3vaT2FUDY034ZIlD/R
dlhvIw4BaE4UBemqoyTLp7crpEU6CMpYQ5DJ9cATeFliGnUEeDGekV6SIsKp
YJStU5Rhi1sMOFm80Z/nVku3laCPirsuqpMGmi1OXevC6HeP8arpebTtXzGB
UxNAi8XjP0HkN9GwqVHg3bpIiiIBASwZlq3JUu/HGZFxgBJ/wCiD2+4Og9+L
4MiXY7QZKQ3BNpYzN1H6rVyZfh4bqqwvy0f2gzwYRelXC5dSlIJLOtvajGT1
JTYL6WNBRQBDmI1qWwIJyCqQZfckscze8TRJHEgoFJ/4ZHsaeVR5bD7JJ/fL
wg/9u+7ssscHk8IqBFp23z49fAKXP4I9FWWyz0pwk9RnzlsSaoHm47fSdu3u
MNoZh1raNCqE1QJjdSginQeAjPX01OD0x7T/zwCBl/LJESJHQzW20B3EIqsd
vEWd4JsNJOxExRBn9P4nQVKdY8EkSVga/1oay+xCSiTZ25SM23IbUBG0p6nq
jxhGsucia1yVx42PGX/lx7RYN0KF1NDhtAGPF3K/5O/pshb4gkH/rbNEc/gb
p4oUAQniBcoBkrlleKZDjBD7OBJKUAfjxKer/Zm/Q9u6aXBFGPPqLFGtIDvC
4ui1DunRZDbdPfJZkHVATuaWMPbOs/JBKLIfXFgIDJZ2d2oBWnh0cCeNpdzW
CeAehi9eDwH2rVVLxJ01o3mw9CMOrJzQLdX/jiqfn+qr4ssIBd/uPbezDW8U
wnQG0D55HcOLAtoFx7kXVJmOOhdM1pOQ89cfmsmvii6HPxQQWvjUzBxIx86D
xNx1vpMP0GM8rG9w9aywTl3g/jFCUHMYyGkZyTX311ziXT8JWSLqz3oYLkuN
r3U/u1fGM+xx4KvyNqNlWRQf6kAMzxuJfY6fD4BWUEOXPds2JTAvsFiTvBQa
7MYF0mtsr6ujdoJWengYNCcftxhtA50nSGPIWLy1ZlMIMs5eVAbaWGMjX6rH
MssJzJIuRSeDx78uNpVWfvHH7U1K7aRS2gCY3cJIbCHKzv0hU3De0RDtWIw6
8Tfmx5kS89M8+7NOwds19/Mo1/svpzgo0Zkee4n5vf39OeRUpZt19wSQvOoz
AWTPcMoVuffUijkw8fjVp2xtCQZ6uB04lnLqxfbyFgohIejhM7ZtzSrbhmmD
dwEVzBnBqs1d3Cxrrjsbe3OSd8rvmpD6mkHJQ/FSn78sSqDsSKaLddYt9puc
2HBS9ZKObRnRWgeGHS71RgBc2UDDVc2iZldACbac+lfAixioTuRrRim956Gx
C9Q8C+ZONx4sAZ2XufCBO7gOy2ZurZ3l2Lm/7TAe2hSk2Y8mvx0Xfdbh+zUi
zxW7rSCSV0/ZHnmcgZdbv/RHPRdoAb3vWB1NscqlAHpPdlMvp/DT/M5/No0e
NIkIhRe6Kq5wy7czujP5J6QTVRq6VVva6P0enIXUMHBBAI8SLRj7ViN8i1l0
5YMHEKX0mWXGrBh6Lic/El6kgZETSIhA8/cJRoosqjcJLgG84eHe2L0Y65RA
fXc9uFBL9w4Trc0S3dQndajKUfbSZ33w1qeHhaX3tFOeASkZVVdJV1dcQ/sR
zGoqyumyC3YcEoCY57Tk5gcCFrfDIV4myAvRc/L2BTMz2brdDUaicr4qo6Tb
ciuo5BunFy7xHx8bFjWBgCC3EsKxgLXGOdrE7llNyLqIlp0fLbI1GlVgKyjr
v4h3uNuaVn2oMSLfUFdknCAyvnZC441FIyd9yFWgRT3FNUWtAIxhbrA3uHjo
58sonszOsYg35sglBULWJJQUVq4I+ybrNphudlkEANjctx7C1sRXu23zco3+
mb+Pntd/gNyjvx61/UdJqfNJEC3DPdLL7x1E4t4doaP6JTAURCj12w2WaQ/Z
+jEVTuDsmbr9r4znHPSbbof2BFsW0P3pnIM4xUWs0+ammQbnrptc4IfxR0ww
ov2eYO4BXM86Ma5vAXTHsbuzw4He27pgNUg9rfDJUJ5icITZ6lT8QIHgSB+e
vyAEhY2YbUKPifgLGkELfV1aZiTwzA4XI0P4Hd4zCx/PpV9a9twrGAAi10Ln
DGGjU/Fap8jT1fO25qQeOhY2nUDmhHOMcAab/r+QE0AHJzW9993nI34HwUSh
geCpydLokvXXiVp5e3C7mUyGBrNHArWy6+s9pfMHYF3Era1EX7hJFStT4Fn6
cjmC6+9tODz4BIA/c4RIojiqhO9hoIpNFNzA2cEVGV7Y9AGZHCLaEbldQsq2
gNONkCW4RG3m00AaH43RF/ZY/ZKeqNN0cGyWg5PfIpSEZW5b8Aw20JNE+VUd
Tq3515tU3UdJ4xY5aenEnkNgflk/LWzaqwZqzZ36xsPw4JCCgsjtQPTXazcy
M+5OCYT56X6L00f71Wv02Qdlv4EakaCXb2CL/hjSG+xcgIjDQHaYu4k3M05B
MxQIEpwZdqK7o/itzXqtowlpNjzEWVK3qoWJ4VQvIz2QtDiPzcuujWgNELPm
K5m8ae4c3KWBbcUB+JKEEyeKYphFJk5y7tvi0gkJBsoLyy2lqe9p9APV7zGc
TuS98mdOkFcJlrQ5vxLwDzK8jvBfzwpWxMlMqTHOOTX3uDSGxOGi4w+WTQBd
NFvQ1BOLHiWSIUrbevmgParcPRa5k1MsWT1pvKOWL0ylITR9zfu7Q7pjkgxx
nj2lhvwB5CTimCKT806I8ePlyv6OlL9pPoCQiuVGZqY7b8sBC1SO9mMzzTdu
kTdD7TK2VXWP1b20e24rcAoGjEyFf5BoMvYhsTfz7Jxz9Q3iy6O4r7rLneGo
KVuLo6cav2d+b56z9+CwK4oow3FFnpURuPQtC4ZQlhF51/wpU2LvA0FytDeL
nUYH8KMjfExmatilxIoKh4WqPyfz5VDBL7iksEF1hske5EvFUjNk

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "lK4MM9NDeLrdcSiRM+VIuNgpOLUAzWAt6nzBJ3Vw5tvBogzjtStM5gMJjD6PMmMyupOFzYouKIpJuOZh/11WnQBMmqEc6gvbtnHqfGmxFaxYyOv1rddc1B279ac1WEgUgi2BHG6DRj+tHk4+Vv2VvppW/Z9gUZ9e40aCxOYZZHwEVb/SJ8ximgD4Fihl81LOgt6U1JRoR0S/yAHMZXIkaoJ6FVEBkPAD3J3ew7MX9EzfFHWmiUS5rP59PYwwT+929JEL4QAfNQ+le+Tdz+MX3ZrBH6nsqaxkIVY5ED7GjyiikdXOW2Xm7/jwKAS40oVQ6VSoSO9AwrYVP0ZgkNePvGfuQ8iszXgBnd/u6tFsw5rJ0kDwsnv3g1q4cGkyykszKp+/RMJuYvKIwkrsQpekb5G3RMxAVq47eNgXfirMFTCZlYwFtR1UN7jzscbWRw+pH6gCfFx3VWQMWkjokeFikhheDifn6eMEfXNpUWc8TIFQsUgubBzqF+pznWE6jKgm19OnL7++mz60TMDYYowUAPxi9/wjigEdKF0pTyqiaAf5o2Icy/lOrrB7tBPTMOmngSl7r95Oiec/zXZ2Q3l9QiPwmD2IidLMIx55nMFz5OVQIlifG0n3D5z64Q5B+ebK/RKh1Zh3Gs3LylAP/834bYl893EtlGPr8zMPvneOHvtaIJ/NYUrlbB4XIN4lkKBfnFgI5HE9qvlqtALbJRG8Z3oDVN51M1I9xQomsoYQc/XWAWmyDFXt3n5E8TzEPU4lWtUvp7jj49rgnmy3bHQsYky821G+pdvKGwWN2f73WzVZNLJno/39PRgcVNrEgdfbpp7bZA594c9vGz6lHvgO11tGpFpx2oM95NBJD8GzcJs0JYxtGKnXNtrrx1K6+86NQR9NiI2Rf7hZEbAtDP+OEPhoh+ypiea6WbG7XxeW/O6EDCl/x3CkxrXvxxwN2paPr14B2TccWM1fqg4YTFcNwhUtGd79lHl70N/AuO1Nmd5YyKI3lVCBh6DZq5zZmQ8a"
`endif