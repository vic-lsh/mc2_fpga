// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cnPZQePs6eLZZkGU6A4uzmYvtGRjSzkogdmAnodtBmdYO43T8Kqze6FWKxHt
hxqJOFkcjoDigyGbm4VjGDjYBk5jvOad8/3K7yr49NNgRY2DOqE5zIjJ91SY
k4ciB34MWhzGmlokpgu/szFYh5h4zhTKv+AVAMvUOrX6jyRMG7FkamxmfJaS
LiiO4iNuUVIhMbfi/xNA2UsuVvxb3iR/BaV2Rt0NmehvlqS+LtldAFMziQK+
Q/c/F3qdDmtaKQEPtKBa3MQe2mzSq4t8/jfO04VjvkIWLI08ASKbCg8sC1Nm
uAkHIjGGjf5Tio/kb32IOXqfmmsVXy5yYN7SHt1HVQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JGVzoRajR/CA+i+E2NZu63oF/o7syRvQQXt5Y44ga9Yz8/4d4pBifCEK66xA
Y7Recq+NhZDi+CQcZBN9RVEbB/kalNLmalijk2LT+uSANAXfH/IJ/quULi53
bcXR0EIomD3LMTS6RmOHfj15F3Bhsd189mC8QzsjFET5MMXHDrIGaBD0A8XN
q0h9M5aNPy/TWVuKSUFPPPyRSNpvbRlB5qUDcIXAGxF1leV9esI8X6eCVlpy
VLtxGF8orEw7OaswqGj2yX4Fv5alcdPRYhZ6igGkZ3B1pZQbd+cHL+Ac8j83
jQtPaW/fsJzlx5LcRxHMDZULi2ZL0VnejqipbfDLKQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LgdUJKhLUQqWWpmnmBkstr1J2/R91cumAidxtKNSJtjRTrduhcQy6SL43Nqc
C9XSXaw33562TRPbobWkZUVJ12L5RA6nBrYBtcAezchyMwTbWhL2u59DRnKB
FFcIAruboHAxWVO6HGc1Hf6+pq4rbeCoZmtN2yb8b/M6PL5pUAwyxphCKVHy
KAH/l7AgAWSIH7XDbo3dSweZsLHzgegja3m/8rXR3th5+zxNaz4a6QWEqal5
tmi9ZO5hdVFhBiCEKUTW0l7Grc62kbGO9qs5BC322qVZYe7KZuywTfXlNstg
MwdQKPMj2ZysUkvIZmGT3N9ndTDW5BPFlWwY16CXlw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fJmx+cRywoy/Kk81932+u26uFxF/z1Ko6bc/R0fQcgU/dlS8bbBvHduKSKLZ
XV0/ecDZl1fUSbvAPfXehikbB3VVsi78vzyCzwTmHQQMrOvycitJAPH5/deR
INhxvK/37MycTU3m5Rb9vpBkBXDPOpN0pbyml3LdkzbFYRSnFMcuEg1pVX58
2zsYTq58TUsn7Ap/kg6Znky61bW0sSb0WQ/afaVIkjTIa7r8Pj0KjfXGAHFF
V3bLqSwhITzFSMQ2EjGL5Ilwy80JeNrSLISEwStv8J9yTEUeJ4vRnGAEDjfO
WytwvLlSqTtkle7XW41sXNMQOQo/wbMkXfETazCfcQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
L7IO9OLbXeKwm7LNYxnl90uRK1ckdH5viSwFJaAd39/ab2pEgBLeMj1PUiHV
8lFqlFhYD28rsNUmJIcEfdRqWfT5MiwM08s24RecVt1BCmdUDZ5Kz1Cnm+kP
ijY7aQuVZsUltIzMPH5Rxw9FPmLvyg0y81APdPAhxIC2KvVi+3A=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
rZuqIiWi0Z/Lp1w32LAvWrtXNVJv97FjJFvSOIg4yN67aFBCOuDvn0/mQW2s
RVKi3bAK0qH2bSjCj2eCactVjUzCs5+ifWptyY6tl9d5N8ZAI7bgLc2qeEao
jyQik/3QD/yYIPUCMYd74k0FpaOMMtRs6iHydb+mR3cruIbIezBD/LkAp1AJ
poeTx1UpMAMIUaxHxS8QLYDiean/Idhpp41td/EdW8ILga8NJtJViXXWRaa0
rzuzsNVFyFNOTa0RiDxJgrTOZd8CrJ3yGueYoyWwFH7SubTGjKfnQex0F/PS
l46ggxW/599FSx/Vc2gOEzqwe4J5NOn1d8TRGY9sDe6ay+9rZwnXTJRBdZwy
Awm3RMjWKfw81DWosWBiy+qm04TLIm+7kkBX7Jh15fEieS6lHawJQD3A5UaX
+uHNU3N4f8j416b2Apf3DzW/wIQq4Bcwm9GQX5KTomZW3mNr6Hz9j+gLqNcL
4myvfDroMaoVyKUe4SEa+0PCPZjLE5nH


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oIJo1kK08uZR2Hm6O9uK77pQzZfrxghI6go8nzUdIg3oJbVHtYLAdjiDHbhA
rh6hy8cc+sEUo5Ko9cIF66s+VEdVRkdHdYDU/Wee/p0QMgd4XRz9Ipi9X3bz
Fsh2njH/HnLJSSxUNV8QoUkgAtKQyZ0omDMA6OnV2rZs9RVd3rY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mNeRE62WFUgFRCf7AzfsBfgkqzpWl356DqM5p/2RMlvr/wjSalOTYte2wO0z
YzKA73Xww7LCDSC4A3Pq9DoyhXqBCGpFltVqkPLD/gmUKZ6reL31qJpDlG+/
IIdsrTQjH11z5/NiV0kq4J/4CXX1u+3am8cvUfyvxwMx4d0jhi0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 26496)
`pragma protect data_block
Hxbm5cFcoEIQgmxPnTEsOuOgzNnyVg+nCocXgU4ftrH6NJg2NzQwFBhJgpfh
ycTlehAvLebJkyAOQFYGKCnhQWfh4UeMWgmAShVbGqai/rPJG0/9u0DuqwrM
Ll9FJiV2QSK8243vR4ZLT1xuDLJ1Gp479nqnGFt6IVudG8V6Hw8qXehhMz+w
YIQqzC5RzNfRFLL7I/ANJqwGzuHqLFkps3vKTT5vZMIkVXRboSImE3QRxFDE
3uAUuwmGHDs75vBznjCreE44EV7K++K8rVgHnGCZVrPUJPhmXfAOUDl1urMj
PUqvEGMMXbJ05LBAvUKejWdnX0KEAaaFxiRmgN3NnRGmbVOZcNR+sfc+mx64
RwUa487lxmhNTJ1UTP2O21S27WFUnAv4oP9HIGgEwtsKAXkFmn8pY+nTWtdN
8PCpdaxwiamiILrssMwcfTMFzgkXTK8BQ+jE99Y1kBdZ4IrUb5J/SbvIOux/
IRbQBz1dcepY9KVRVF5a1dKD07ccT6AGN/P2+2fUVt6TOebh3+HZ5Uryjos/
Q4AF5/GI6kDTyQQCI6ExnbLS5pdvtCjhFCMvoH+GfKl1ZZ+Ow5WAd0NdrfWy
tVJYirXgqXM6ofT6bU3u/bCdrKQfe7ptfjIKXwBAix/01FqvxxGCHkNVXCl2
BK9pD5s/Z5u1nBwrJW2wmxfuc4UkWeNRX96s78I0/UkKVliAJRTSzU8Glj/z
QMAyhrsATtnqUaqz1P5DWtr231kUXV1UzV1xbvO3tch5d1VOtkIiLsT0xCCh
qNZsJdStS/qL5mz/6WaEQjOJflCl7Dh1jL6mGuQ/rsFmQgLaGf0Y/xZZMe6Q
Bsjq2wmH/HuRjFHi20RhYpeOLqHaYoNev5C5PshhoRzgqiloAdnneNro7HsV
T1bXYXP4s0x3pUGL0vaRCgqpw7d4h6NzgYW4+sM26l8bo0LGMW/paGVYp4SY
rwuFlRfBZc7fkdhmXiX9E67WyXbWH7gJWXzw59Qs46soXLCDtzAQRwKL5Y0P
I6CeBX6QzOUXizEUgq1/lwU3W14rCOsZH947V1v/Nq3LztkPBiaAQEqmqpb/
RluWrb2ajeREHldXqVQOkwqUdWnTK5hne1axteCVyUVp8JsaArK8vSHKT1HY
2X4pBWwtr19w+8HlRf51Y6Jc7bGAew137ZynjbaGvvckPSNpokD+UTM+sueK
eIU1XxRTigNLNtFpwcOH4rWwgtpwDT1rSqugtGFjBQ2daDdG6+9dCB/dJNij
vWaIbFUNCHqfg5MCw3VEnbYhgogiEkiAaRJQSEsh8A1EGq6xUbnI9vsjbk9X
VSc+cUcVm+iuA7X+G+0nFGi1M+DHFeXwwg6qS1bAkocHo0WX+4Pjx+/hOysr
kg0yWSuP7bYvjWpzchjJOs4+lBoIIWx60VfDkIo4QuqqUhVT9IpmmFSh/89u
i1jHyZ87MV5mV3dAizjeGWw7MzXRyX6D+Xdl9Pt7i5ro9aHgfW5KIjwT/VPW
hitN4FxXmG2GmKOMvpjVwLTLp3ns5MVpm/Q6YErOzEZLT6qX6unzQ84m/iLt
VeMj0iVTydDMd/5ehktrZGWoKv2OcJpe1EJHPOeyzMLiZRYeSlr4obCH2NT+
Jsa3A1ha2Jk65nr6Lq5oIRaJ5iVKpw0CNRLhwTIzZsoCmfy53G8jR10yNcmv
CHpkyyGFI4jhDVX/bazGjh7QRQnrdTmAONjxOZjTdreQYyeevebtEhs7avxa
L6QjN7JNwqrTQItgSI5Y3tV0u58gIFxxFjFtBjcFFbbGmD1Lt0PYWC0eJ5t2
CTvdaQ8T6bthDe087EJCOyfzsGC8EDc2r899sGDS9xH0d7ixm4ZMr3AO/0bd
kPBTA0lbgjmw6SMfGCMDfEii7ZrKVNNhVG9MOgRZ02mO+9OuoWujpRVGPQPR
m063XNWC+DRG4rKs8MYCwLzkgYgPszlkd9vs+lTJ2q2kgHjCHqR6uYmdfvMN
KkyW6E1bV3GcMAL7ZmrZDS6jC4+BHcJkFlDtna5eiaBI5+xyJIiF62Wn395L
CTNfqNm18GqMuG5QDdeur+wGNNItIVdYFEiYEoxSegBQ73DzNiRQIkLPQd0t
CvXNDAhOEaqcypsML+y4grXp7m5zavF3Qb5Q5GNNN/QnIeVpZhNx8L47BkYS
YAxBgAT1sSc4hxZ9Rdk4EGo9BaatQx7YwqaBIXZ1Qa6PI6fszFQ7vyNgMKSV
mksDMrGhDRMZDRFN+QFVRjoS+0Y3xzYn3dyKTd5tOrJayU4vRBYIkpKqWKMu
ymcbiHrqi3yx50inAGK9ljCFpVChMK9EhrYHiMTrnY4Rz9iRLQXQWPnodYcx
FAUEitjbFlNFnjn8lqlDMF6l2oktIfpjYpO3gwqHVeLtU1XIKtvWw1pPK+yD
iCKd1OawD6cTqQg/ivbJ7zQRci6ikq3W3riMAx6hSnyG8mdSEVo7mk6ABMbZ
pnXSQSfrXlUUm5kS5mrj2uum6+aAUeD4AA05MxS7V0LR37uDsDoSyEZ5jlGA
yWGZzs8T5WG4/Zr22oL971QBlYAmusJz5isA6rjimefm2UUj/Rc+ajfzqy+6
Y8KWqr+dw7HmMKAicrdlWID+BOPBGzUkZygUhJL1D23DEoi7pXGtNs1O85du
Mib14gye5WSZRq9TUmg+gwhBs71pSYw5dI/k3WE4fgH4d0ICxvczJdDrWmcK
9kSaqOR1a4BOi2AIEsLN4UPd/nTBGYpTBoGgRKRd/uN19ZDagipiG8IOFqOH
euDZ7hhNvsS9kPLmTLLvd4Nrc0Cjj75uOtVU2WLQMR7UGvoaVsqWzn1w2njW
N1CtvXu/lcse6r5wBy9URFR8+B72hd7eu8DBewMxwMD7x1n095WfX59F+zh0
BWs9tbUEYB0RruKp4HRGwWt3TxqbpsTKKKenJGpJ+Y/DCY45y5ZxFMv+355K
oJ7jwwrDE87RD/Dq8ELTa0jVTh0ZRenj4v7TXWscmG5jC2V1NA07BT6yu6nu
8T4M3oPyDpEurDJFP33o01ZXFfJTo5LR7e19b8A4hXB1hXzIGg0dMG4h3yJ1
lwTlvwlIeag8Ci9OgynRoEmLAVnyR/LIGlA2E59i+L2enpe+2RFHg1kTJtQy
aloSR0hOemynQxNFcPofRjn5ID+4k5UENgTCBTRzjWhaGcorehIglJfGQMT8
Uz+r05s90DDkYiCPxc6g4ZC0l2BFBZRF7dGtrXhdb6nUzZQKSNA4ezkLhptP
u1fXH7s9ay5FUxEYZpfCCYkEe04MJcs/60pSgxLPnPfWSelYoD9OQLQeYR38
m15jKtN4+duGZo13tDXjU6ctqalEaPKDVG01MQA8GdqEkro8QeebC6bqLvZ7
yEvRnH12N9gYO5nwFKUZjrBcj7E3pGxY9T6OHZ8Q7TkSqeVt82sFHwqFrJop
SvJmLehJRCmfqR+QYkQxSya7B58E9vTBPg3nTmnBS4IjVIBjOHHMIedNps/w
tIowQC+b8EW/1aiv47yOeM49C2zSGn9K9SIkRA63dKRnCjLHzMrg2JOh3Xsu
Rkl99f9RSU28cOXJlLRXYj2d2X3qYigmqkiiodox0uZKK+WnD9gXVUx1VPeb
bY0S7N9wtm144Vfo1DIr16TWmI1IwWNhruWOOuItefK5asclIxLYpQsoM9Ps
xWyasMkmgvXsyBtROBHcO59eYxJV3EHv7G9Uh2+kpuFnvd2EeU8xLjfdgnI3
NyRJWwwqjUs2NOyAc4CmR/i82Sb7BLncz8GXJA4fGM3/3eOQKFchNmnNNpCG
oni2t9fk4WeCHW1PmfW7sXXk6Hl8w7EN+o0Ho0pk7kqpqtCp0McqxjZ0QB/j
sHJd17YaJgGySf5TGM1wKM+QlTDlAsIDyYq1pA1DwRc8gK0hLS6X3L1eoo9x
CHlfcSDtmcPmMO+tazJA8gBf1m2U724AnnR2DT8RAxhEwuVmq6tHteJO01s8
TQkqttdocdquNWMYR0OEP1RpmZyDIDw/jnQL0ZUlVpUk5FzRCvMy5+Hem6jn
5Zc7sUoJsAN9gGw3NLjL+iNFUg+a6iZUMA0sJAVLwMNh0X4s/JWboqNHx7oz
pD+ziUd0VQODK0Cxrp7bcP7bDtAHf+qRNkKR8BNkIa8AFB6DH7kwSlyQxD+7
YQDcRM1UwzjHgSo4fYcRPyHGVK8SXxmA+h4101ib90oV0AfyUJHbId1xYOd1
14CbXuUYPvOK5u5Pc7agiKVTRQyyeH1mqkdQa9/cJt9K+FZooTMXdgR/CMyp
4NpCoG5W+bmwoDPvlOYXCl/EQH7LswjkeggOkTY2f7AY8CJM5RUJ9RGQT8uR
KZcg6z9g+zn87TFRC3iX0spSxbH5iXcynfZLNTRXFpM8S9YCYEU2pjbYTZt/
+HRcetLhc/FIh74Rmk1riIuDQ2YHMKkZlRGyz9PoufyNrWCxiY94GExonhAu
c9AfXyNY2fYnnVfRbM2+tWSJYzfSOFl+yOnagWOomhQioqXqHJKHnz1cTNSA
Nu+rLdTmEJkkiptcj9UxuKRscJFQh+KkcPDov5F9wkWx6xi8te/6wOOdW8/C
uQPl4wphsyCRV0Iv0S4ew9J1MrlKrdLxoEeZwWF78WXmU6xgmBoZgGA+P63o
8PsgJYZuDVdMdKv1drLV/KuQvNnHImlbra5UY93mNFMMSkbeKBA12Y0fBUcG
acDAayKN4g2BziLA8Pf2kpEx6Ru7ElJIvqbPGs0PCrCfzI5ZBygsDcsoo0lE
FGtVEndnMl6lTLTpwiOSAAWc4lbxUAyFxt4sNQ4Fj1DmkB4zIftW91Jl0NI9
llvlne68W5xsx9wlusQW6ftaccnCY4ahAssb5dUBnZCjeJNoHEO3xfdXxXo8
FPRNZ2yN3D9LJfPj6vImrjR5yE2S3t/GTmaWa05+pIpPrn/aF2VNgtC1LhHx
i3R11AQR+iAHfY5l4LyKTnWiNEjN7zEYzBczbGow17Da8/FLlyD/BUYawh//
ukPT8cupbd5DzCbIgPxXKTJ0Owhc94rwYi/apB9DYQxraKUNttWQ4vPOfvQT
dYdTJqak1HO5Gfu//HHXXwmyTmj27psaVNsrt9JDQzMeGmlHJvucGeSRf1Vu
hYY66SIpO4oFo56blowccHP8mqwUDPeNz6PHVAFuQTHPNu73uEhzLYuz8dwD
pacNLbxV5tfoFHJTe6ecCzVlDxCd06bPhy7KFBO14vRYMjwo8ahsaLRZR+Uo
lwT9nxlLWfNqBHu1zyS//zVPtWznttjPtOUiG+AO8zUGVMsvUGUekUkGM6xO
uMbkIKgAsDH4DD14yMq9jLjKIm4X25lBv2UAHsdmcUusRjXDIKVgMBdkdZ75
z7YJFn/BLmJDqPzowui2DFS9PddMVp6Krfc6odC4Cn+0M1KfvEe09MY/7tWm
DalSzQpNrNNmJbH5XdU+/+rkL40vpEbLyOOrhRpXvlB/2naYVgH3ME2i8PiW
OFBnG81+O7vGXkEKHP67SW6n+o2CcFoKRih3+urUaHZWhNlq8n2gDZ2cAQTs
jSt8X/v70NWTgueuJzIfk58oX1jbaXRH+wIZjZPwd1dDwxCQ9m0MbBo9ZHSi
dGK8uVXqunoQBpHplEmxoXUpWX35najhOo2DHPl7eR/0c86r8BThSZabQvWi
nQSUpFOl9l4ZQUL6TI3hEbBMKYVf0LWwTyEyHJsvVCI8Sc6h1mCG4OlWPfZV
ol7DTdMdj/YMCOjvb13imAzNevBqeHVjgd+ctDanMf0ob5cqWDJVVau9itpC
Zf673vM0nCBt0cegmTKBHhNf1xY7VRZu8xPcmw3f0dfIMV1xO4AMAMWf4WGD
4AEC64XUFnnf/7Q5oObfwu2dazxulAdB2Eqs1fxf1HYp+smvTlFY/E9tV+Wg
EcjFFd/G7nbzvhOgzphfi+1HFnpf9QzI2ZoA0XeDKEUor4j+J8WwjGAxPUDQ
Pl28633Q5jhTWM6dgJP7gflvADGNmt9uaZkA65R3vmE/i/606JVaMsPNeIN7
wUF3qoBOTk3cBjuuUhbOoRB0TueOgO1NtG8nZjZoweHfC0lpvmBRFbV287qe
UnE1pWhsEsqQVp7F2igYstznv4dUKw0PCCgc15hvdCatV+YZM+oIk+jrmqYd
Ah/GgEt7NERx2Yd79t/lFjhTqQXsWD+YZA/IWgWB0aHMXOqp4Wg04wH1LDxb
VXDD4CIjYq+q1r98vQrjhMqnE/pTMJwvxHoXNk9ie5aeX7DAnZYaPEgSUnQm
BcruKzz9OuzomwVsd/7guSeL3rmwhUMwgrck/G+A2Db8ohhW3cnZ0m8nJJHs
PD0ZZOv6vO1aH574Rj35/pg4AkddoA6GJFEOzMhbaz+lkfmOMWEo8YH1Lye1
UEgGtpApj+RHhvNmhikUcpSRh4yXGjwnQDQ6SNslCgo/CPnUesISBsfyy3Hp
N7MKztCzoXnGFVRr5gGwb1CmGqDuYt4+Jl75UeSRJ1gl2Rguo3VhLRMdG08Y
ynWPWf7XD1Gap4vagVf3tfPxEFqwdePA1AhQtw0AE3sfC4nT01Zs1mwCFX/Q
nEjo9MknZ9oL40gs7bavFtmMBPF13AYCDoJfnWs8gbG3SbWoX+SqIvQTj9zr
9cbDxb7MrfeAV5z25YOGh4PjgQTulvn0whb84gzCGcxoEXFNqR7LquadyD6p
BbRanBdO4vaBneqV0Vxelr9RpU2rZVRIJzV3TI3UYVv77QtbMXctR0Ah4Ih6
JsF1+WckXTdx1RdfXLvC2dAE8xeVJsYNeaY1KWzTIRKoxTzKdfQmUbAp2paU
yHOnnCwatbdRWA73C9/WNekwoeFsIrO44FKNiueZo3Idx4P0FRd2XplaRFNS
fslPIqeRc0SLN56VKu/3dZpYLBSSmf/UvPXIEQAb1XHgXZVlUESqJVQmQFIx
o2NEqPqLJX+QAJ4zlN9w0CdRb2rZRgyYOTh0ayMv3xzp9xK3YOQmgACTX67G
dV9lxj/JtRTaxJEXqVXxrY641iWvZfEgtRM9c0iHo4taS4t8mxuwwRoOjSE9
CmRbow3PbPJMgavwlXB6FVhGn5oiac2KaqHMF0p36Q8Q3+Wst/lx4Z72+u2X
dY2n0xHYwLpvw7t9gvgxTDP30xTvI2/Yg/OILJesgYYGGjFgD799A5IOyoc0
//DBJkfLHQyCLEJN9/Cw1ybCL+OFUBJ4l/Fxj7JDR1YIBOsIz1JKQXKJ7WO/
4xGFGQBdGbOdd4je84b6nFziUtEW/dM+iFezVn/Ahyl2juN+BwcYfgHMYXsH
X51rjtgKfJC4bD600Uu4SKKGgjyJ6Qi5+ynvrdDUyYAHwNqkEIBEXXonKYIm
UOG5PWhhjGtu5n7IJMug+1b1PVbiogRTQ4usv9VDb4aG4X5DJHehwB4kQcgM
d+OjRtvGf4b5heBdpH4ez9qPQf9txB5eu/Ps8XNpCDB57oXe9Ea36AMCps57
FrT0X9TjiwHdX4n56Go2UuYWHJZ41p9gsJ1LIimgdMO6EZR4zyVGyNPI69Bt
O5/D1s/1MvnFovP+ZdzQSP3a/+9I/z40sZ9UL7GKA0RmkFJs5/88W0reS/Wf
nPumF1egR41zInmFHgJpZn6loZMtl2yiD8H6I7B1FL59WMHrpMKzcJXPUucb
leyEriihASLCsYhPVXpXZpmDNa16eJayk1+UgbEHaHCijdJmbsPOw5TJzk+3
n39TCOBlFQIUxfJOFj6SIP1chU77C51fwQ+J6ZBDw1rrDH6gDQ3lot1y7H3M
UhFpUUjGFHCwn7MK7oiL/ePGJYm+1/0HXkpDwCw80LEHXD7c9KiYN79u8oCH
LF67/7AfN0xgbgZ+nsOOwOu/c5Knu3Wnvo8nBRwC5bizcXll3tHVs/j4bbU4
w9nKLTGyxtVGnqDejyteQ7mEvuFLGVzW8kSVLydZgj2aIBbZhlwLNbWVcKN6
KxOE+DpqkbbnTJc/gUU8oojy8TolfkQbEPbKrmipen7EYpVNmN9z04zfm8eX
639000+MK7SUkLSah8lUXkaVj4Kc1FoO4S2a0NgVmldSx9n63p1vtNLxL1Mo
AtNCCMJqJrY+D74x4n5XKPQYJc9nfct5HgYfGQFvs6rvP/WBxmcZqeoF2VL1
X6cwnB/c+yI+8f628ov5FqokvPLxHe4SYx6hBqBbH0Gz66ZmTWEJV3/5u+QB
ISu+xGLszYtqs4//GI4LSeen5FIdM73LFh9tYfLm0iMYMtQ1j4X1qwzwdxL+
ne8tIqTSwgeWZ15ROxyyDscpf5lJllmJLBL1Y4DlkrYyLJ8EU9gKTw6Epkz+
t1TNfyTsa8W4jQ0PcrvYWa4c7M1H7zQ9VwmpAnaBmaildI/R/+JY0rSV7/Cw
88Y/LLQmkkOevzl4TY94TNBS5K0vPxFCZUIsjphulPMrjmnjhwVWuB0heO06
3s5W1fQGM5sbCGLgdX3kYMyWa4gxfI2v3EP5HAHL1zu4sWBHnWhA/OvWUx9p
vf6Fm8i7RqCpTrc4E4j3Tz7ps30G++B/4xgzljNQqRvxDGlrioJNZ18JSVRd
T/uBchNePZslcTGOvUqyAfxhc/ODw8eMzyG8xeXXbXJE8TzXrBShb+TEFlNq
JKz61UVzG2TavESTL0lIpzCTbNXrVLhmLl15tuNFgf4rdZvMIrjEaYyNlRLL
7cHIJS7aDxQw8iMrL1Tt338xdiaAdWTIKyfceyA3O3WELPIbbFlCeEamxwE5
PoLyURnbHto8OzPx/kLm8yDs3u5lWGtb7lhJ3r+em2bNn93T2gC/jy33ytUe
muR6GbB2CwKponw+0tCMQ/igfEJeWGcxR+loofZ5Ls3SfzXek5Y8CFLJEEPg
dw7SPgX3ddjI3yTjeuRf2Tig3vrCF8Y9QjEyuvMDrMS/IYSz4/x/t3xyoN62
N4GMplu9wlLCDad9ianzZgFaY8jWrhtqODntMuq7CxNkqI4G304KWjkctTMR
M+RseS754VTktFvrU5ptx6yIaXwxD0G7hx0DwCmpboBxNr+CTTBk/eXPxV9a
XvScyet+mHFFY/0geuBp375S0DdE//zSe9jWf8JB0A/0uRMgrrx7vtykmdxR
HuGmCB+lKxz8luTmuPxS4DtMxZhsXRseWjqUka+I1Cl4h9a95xa+FaAXEptZ
6HUt/Qvio36OV7hiT1M0eVIbv/dWfNgEbcOEVZjdfgH/UDoxf31iOOl9Kmy0
+EDkpaKlbSgHBYxnbRBmoqoAJsBQLTVcqCOwokL4yQdKJX5DgGdgIOP9fMWh
xff1RFOerQPXc+0ScqMAjKpMhsB0xm3VlINsR8lCECMPonGl5xH6r17eKO8F
VnYPeVI3v1xpTBal839F2c5n1Fl2WnIC1RNWN7GE7ZpTmllRvpnxLD66F78h
VyJ4ObgmruM+JAAdvXcoGsJeYmzn9kUukgyQaqn3M9M7O4gq40LiWGf3tdq9
2rYpo4YrmXGYF8iDsHB2BwvQz/qAEkGs7eAxunYaFCA5bAuwQ9JEDHUq5hen
ipCX/9dglkYYBBHAEIayhHMurYRBbf2t1Ryqp7/C0qU0Q5ncobr+e6fKrTlw
mr9Ndc0BH8wBya/P+CisLERfVDu1aafVV+4GSRl1gToCmr6NZooVlCz14ik5
O1Fgn8xigFa+U2iVKPX1EO9fWFijUA7S7co/nd/qB4n43x/Jx+IN5ybi/sBv
CzSTgLFFkdp1rFN68hnEL51ZqcRGrNrejeioQgMwIfCDNLas7a1gqJCu7PXm
3vaGv7UHUgXijxAq8Hngbuno2fmCHMq2e3UMFVicj1Nx1cmJDsvz8n8aaflp
BFDi2JgJe1v+kbYZNxPAmWC2D0M9z85Qy46HTYUUL125xSe74jPt4N89W861
KXkaTAtMQ2XGb7jVVjE29EeH5wmaqTZ2DF6N8cfyKGJzsZNUgINALNcyBcnj
un+Gc4qMazIFPnoZl6PfGGUOqQYwPJEsih/izlOCWaxyScTTaeWuQPdEsCTG
n+h4VBjGB1XK3H7x2hQmKBrtN/YdEOV+3JjxCHLM6gJgasGCYKn3Y1A40b2h
39a18xA9Izmp4hg4Qu+40pd4/mj1FW/W9C2brCzyLgUfslOs+dLh3DmlgSxq
u1PeIT1PBQ4Ifs2GKdqqrU9US2s3CwCixRaZbXFXH4SyffzubYKiCWRlPNct
4pSyN/LDRiqRiMhHh8uimonAoPqh+WtjNxgOoXG8WQt1KEWr9XZnNn5WxKwP
vq4RxYsqZfPqgVDxxlrsZzV45D73k/NmP7G7b0mgLrUGApigxkcUZQKWN0Hp
VSHBRxnoT9P0QGiAE7Puikg2h52+Z+c92GA76sRoJkDvY4SbwSDVbeP0SP6r
w5G8NKoT/4cia5AAfm9K57UcmaAA2cLE8b8NYQRMa5t5oSvkug+DNPrkwPP5
GmY3br3M5IU/eCW7ZIwgfVPBKe+28MVSq7UD2ttU0n96TLmeZmZnjzugskpO
OQG7zNjVEmXVN9iVUKnOfNNSef54cG8OJeKCxmfFsN6wtOny6g/iZsklCkZk
KxtJdBn4EPdHYNI8zhd3vJMOd0HvNbptcFmV1POXOy9jonCLZkk4JLHENMEk
M8mPwuGHwd33h5AHcint0NLEZI4rge1Cj9X48zzC788PgvOw4U98V3/83MfJ
pWddmGTum8/oyCpxjahjbD0XS/aDHjTzUqoIOqyhBM5F8kn/F6jyXRWC3uNV
ieH59oBZE4PDGIzki1yN6sr1tXRRf5FcnDJfWxVpnKH4+Rtd8JcT57XCtJjz
GcRbpPavElvpSbaNymWzQNtuQLEvhVUlgRMzjoVgADaAxh1sBEvFD+Di1wJ6
uJ1rmD9HyNGauy5Zdoiug8QcHXe8Dz2GbQ0k/rz3IY7hg06FnHxfHIwgFDtx
nT+Ab6XM201AWMI8ULYf/j3Z2+yNSqrtj2T0PK2Ldp2g58+RQaBWP3q1zSCD
SEXgFDNkWw3OR4/pvRZbYwjK8t9fSDYe56MN5ufhPeokf1geVP5towpmopPY
MxSn0MgvMKwqcXsxvPXqSjE56g2nsMm12JNbom9mPH1Zgq4m1UoXcFDHRWz9
sBhUsqe/3CMgctqEuA3nfoHe91a/kJQ6igc7WAfz1420+a/QeXYcCviLBPtf
NZvvpjpuJBVDCCqMtjExsFuBr98GOEe9JJAWBfrTMtS5EMS3ERDLufyoR9Ha
59d9jzqBbdORCSLKIZ0RRuGynD0dH63TQ9dqDuP3H6NPPTpJHCLPdMkyGRr+
0ke8/spXyWtLF6VTOJK0/yWwlBLCtJU157zfd66iehf7lpNeYqUVboN2vjAO
jH5DER0A846z8CR4IwipGAXd6vrg4Bn19uYAm2+jIqSVHDMloGwa75RAMW6U
XyX78LWLGitnDr3BvoAS40gApDan0s/5mE7CEPCeAanGq/fFw/V1n6sT763T
7QxzKwkQV0gCE5rpVN0cqcmp868K1eshMHOKVKpQSFfhl2DCrl61mip6Qkni
thGBgXzfk8/DxPs0NYzSJedwG851zVDsq7H+yMOCLgI0H6mpKnKf28c9U6rW
o74xu6aVtDN8P+nQMcyghCCIbvfqe5q0noWTHhiFCe0N+jUXVz1jOBrUqHNn
aRgSeJ4RaMJcMjJs0z+9uPI8VsmDllej89m5AqjtHx1iv8CIAqtvx1U2g2yt
uIibVsaDlMCykfsGGsqaxWKnuqh9ON3WrqwhVMdCfs5quMtpYrVeZQ2ze8fv
eWoig1EeIxT0/mJNeOFnRXL3nNoHiHTZGv3cIMStMBNCxRsJZvz+RSdhuKkA
G+e0PnG+65SCBqDY8hTUKBAfJyLJt2CJmEzTPbAb4T+//asCKBKPwLcs/a9C
29pFF58Nx13AFPYn500kK/QLe/6hdp8MwnE3MbXRJ/Yd/CWN5SftdaAuQbCL
IJBZ+/oI/HdhmTf+ZCPMeTUFqWMop/RE38zMHNX0aaeVi8GYFDiw/alnjvbj
ZsW2v6h5sNh1o4nf/SvP3874U+4442yIQZKJJD1X7YOdAze5zpwaW0TBqfTl
+qdBxm5roN+qZQm3hCdaf72MM0G+KF9/mPBptQ2ulej2JIQR+er3GiFP/wfN
SPt2aKHVKc6wHJ+G+Fg40RU6ZZFXqeCxb6tMI5Ke9DVzCZXVkTEwS8SYS6bv
DgN739AJg44CUYiqRTbqgUbp+RsN/pV9fWC3nBX7QD00BgP5zCbt7IgIjAle
f1pkXTliy8xXuKKv9R//qJf5HcJMbrg+O/aRKctjWzcIA+Ic26nxzYTWzLMo
7oIIpMjt1xxmwzZEsPgSREStaIgRw3/H23WBkqU6qln1u0tUdNFRUNB1xnLe
JcAqqyvLzeBuxlVasBO9w7oRWikNzN5aE7wZrU8Bsp+SgLPzzXCDyT6csFBU
mJVi7/petltth8D7QcB3Ve4qcehMlGEkr2rG+gCZAgLZKnJC4h6fxo0ek0BV
lKIOIwgAQYNq6YStyXwR6n8UYgpvuujRAYDdHRdVHpZakOZxiVSUdaEDybLl
YbtfGmRuVJfgDc0nVP8MPS0NCZWIjDvB6t9OvVkAXlCcUd23yHJysVkCwBrp
fWfr3RzHoX0AkCV42lkzs/XCzigRUdgLI1jTQ7lIwz2V1Q1kT0x5r0p6kM1h
pAQudXrAqQBmt3Qgm9yiWkdTHnFZNKbybJVuqIgFQ/xuQ17TaDzWB9oLzQOK
auyyfIClANemWusuYWm5IlB7R2fHRqQTkehNqYgumKLnzd9lGTawKd5Ave/w
dYPvG+1qszTBn0sC4IPl1xHNvioHAQanwnXHBEcKUBYlDpwxZ3JXoUjLAudn
LFvZh8731dcrL467fE1vTxR4wGLVfTFrHBuNVpQi1hpznOn7LpLnL7wrfmer
A3Z1WQEWaWzukWBsBbAZpKTcTQ4sZMko74zDNs5MzRjmJunjlMoOesHkXh1g
IUx3Jw0AXaQGt+0AWipndbFOW9laBg5OvP5igTAI0DTM+NpE79B9cKr7hwyh
y5+t9FKwgu/bt5DlViSK5E+xu8XaXMP7wpZYEA1U7T/q+gsqg7RedsUt42sz
aEh9qpZWGFhtbO1NpBIBA9vyN7Ra3MHTBV1N5GnSjDXoKDvqDVP/T+2ZxO5t
OUO8HsuYxLlbj54Qxe7Tih4l1kBAKmiZZXcHQFZzdUB2Ac1XSp3yg090IGzV
bTe3Dq6TmhlvIgcCijhOnYRDRWCM62pAU8yBt7F8rh9sFw1kZdMTLK+wtzrt
yMEfTSNlZ7mbfIEUkKYSeFe5/IEH/51F4diPvCSV1NVZosxLNoGj12B8VgRc
rLPxVp2AbfdDCcr6zq/eYgjheoLwuOJ+7V8Yeyq7zdKZXQRDi69agiZK8Tn6
t2oQLQFPXPcjrb1YIonjv6qod0NIK8YNaZ8e9EYXG8RPd558hPuukq/0Kpy+
3aiIsaW9OKpvicPMcL2fIyTZRLmcvnogYLK7Lfacgq0E2rLPdrKAqfO/jKBl
qBJtN0yy/v2U72vKEUHrKKOeM1tawViIDGY7QlbzeCcsb1yNttxNcR/uTvUj
j/j1uqnW8yHDNuDu4WcJjViiEazido8y/3kSCj7xAjbleENpql4xKglBR8xr
2E6GiqPiBUx8XTCkVRuWDRlP5xmAiuTn0Zg1JJFi/esRQ+oc4gTF+J5AhJBb
5kcxgSiVgAThtNS0pmlH8D1/V8sZ1aDLxc8DwgYG84ywudo+8MfKySblLmRG
DCO4yVeESLA9/hy3+5CjADKcLXzbu2u4nxZjDJrOL0jW3Nr38mOl/pR28fvF
MS1Oew6Gzr6P7NS/Gw4aqFWc2BACervUrvXpWAWWpo1G5BS69duyF/11DfWM
5cakRu/Hatq1bauGXuG0jVl0HtETlei6MrHYGteDkWPIAxUPyiMDkTx+9QNp
KKyaTX6P4qASptJ511QTE2o2C9R5+Ngmj5+jjssIJXnhbzNJpgh6HIR09KST
FnISkJJFzoHdqm9WEeD+tbW3xmDmhwWrCKm7HGTQRLdUOGRyp7hAfBQtFgvM
lChjMPZdu/mRcFWCJ7I71t1PKEGODgVNaLGudax2eZQO4bQyIj271G/psBfW
erCbuIrjDW5A9xvQSGHw0WiQQYI/n/Fqjdvfbnzmik8ignLpN+PzdfkrowOz
7z6gCgM8OW5GQKrkSHAzkliLzTgqt0WI4zd5gAxOEBZa0lLDYlrzuY8JGh52
zuu/ZF9TnPWkLq7Eoj25bDmUbBUBWFtS/ChQPBOIHS/nZo1QV3auDmp7DtFD
SDxIOTmq63RwPBK3Hs/YOlKjnDafp00EHyY7I3exAu3aFaQST+qglIxSrQ4j
tu0nTYh/h96vhsahSRNasQ1QoTvih0OFOg5EPcmYp8jRsrvzLdLPLnAGAd1d
k4XsalUjwrHK4L2j1QXhKUuIZZtNnYaFPBMPXxVoEVUZVGPkqIsvpDBd36Pp
9AV1ekIdmvDL/RdhJ4UPNCnK5ZTIcDbYohH1VqlniMClvvRa6t8hnY1RVWL6
lFL+s08FstRqvTD+3JgnuVdt8Ztx/QiGi54m1Lth74XMq90estRPj9O756EO
/RUEGldrl541wCJwK0yZAtROECHX+WCAz+bZiqv8rNr657/ZjbtMdz9pm9v1
J9GmEoV7buKHVofO+SgH7Kk4mi0HgnmBTJEpDKpFrl7uJotKqoZsZ8zGzV3Q
CvK9mawXFcd/8Q9RxBCYNLaRXCAO8Y719SiTAMMGatFDh86NidxvIXlTGvp4
EZ00JUFjmX6q1dh3uuqucDT90BnXswpBRMSEKthrztDh/vkUKJjwmdjiEFTA
J4z3By5vL+fjWlZp06cWmf1flSl+qFuka6t4T3h0vKOneX46L3H5VMYMCkJc
mbNCQipiyagh65ZZVZCv8SEG5MfRdqvbDlYnZI7nhSyB6Vf+7MJ22g6eKzxw
mu4HdIjQIs1XwSIiO3oT8cDViYQWy0yLIX6GKUv9F/e0NlLLl1bhglZfh3dD
91edxIIvTbvojv8TyHYugmn62L4gSRDd7dTlRSb2dqxQ95Wo3dCIYnYitYkY
PtETq5Kl/Poy3FgkU7z5Fjecm71SI+tX6xWfra/bKMO1TJfZ5v5/cjRjaVMl
Qyyqd9XISPksSwMqNh1dbPKtxkjIcNjv4l7Y0onAqTZF/GQffyFqSFHmgW1K
Hq4Jfd4WwcZokP5adKVLUxd9IeMvJeUHKHhjZSI1aY3n2QEUSbtBr2OQUbBq
osxZAR0LujbbWIS1owgkxNlhMCUFlz+zciSGCPudYGgJbiPiKOSyaJLNnp7z
9CPMaYOtQWoPPM+fKlxxB8+1pvai5Eg4/Zyi9UktJdHcxXYfE1Ub9mxFW7fd
jz+4w8PzRHLpn5w41M9j/bivXJrrzUDPnYokVWIUZvyZTLe4qq3GThlbU2lY
eT8eICLqEvyj2K/VZf7H/wcUpHv2GECb4B8WFYwY2LFIu3YscuMqLKiRGBXO
dKoF/gb2XPOPO/jGBkfpGiMbnTpLuy0kmXIKt5JJJvzaLo8TYuX8jRewjsnK
5617xHLw6cOVoeOAwIOJiqLuEmBDSmL+G+2hFNy6BsOmPuLCjClnCdI836p9
7xKya5GFuU/jnoE3KTolkMxOSwZKfENjNLbqBa4AIk3QbKilx/v6cSiRgnKL
yEmoQ6OMmax0UCMn+6Bs4nQ7DMszPyZRqf0v8HpbAeb75BJfVDOJCLyg4Ig3
LznfHpkz60CRMLom3M9+sSYlAOziPpcLoLACm1wJFxr4xp1sNXgCHFa75OOp
1sY5GoGyYGRBW8RXQfBWl+WoAeqyVAQnqSRBtJJkwUCZeEGbNutro5RsZAp0
f+oNAnEzyShKJtMYztWOkisQO0NkjLnCPXP7VDROtsR2UMS0OTjKAA+GrA5v
E6wfayYSjJ4vPRCcpoF78ZhFscuNBCxNCncgotMqQb2ObBo9+N+ZuS6MXSuz
TUm9jUHG9til4d9LVS4/6DTGEl32D2M5Jl92Fu7usZo+FVNDg02ZzVmoI5TR
ZFCM4zPxgTvT4NMGRYOMVCKN54mDa7Pk61yiB+Rbkw8TaCTrCHY6YV0SR0hK
49W7DaPIoxZZlIioKC7GUB3FAYoqEXxt4+BnksKPhRKTEEeaFsRnEICVLx4L
3pGe2MPu7wxHQzHX9qegdJB0AaL2orpiOnT9uxjc2etnVmNXzx2UgaUuT93M
3JAYYWExE208UP/2SAbZZho6u08usCIqaxeiR704EGtJwu9Ty1mAYcYUy2R7
GiE7p1oHqkFCuEDafIhkA5uSQPFCU86mChtPZnM0AnvCmN25zz5s9zhPghRz
MRY2KmdQR4rwgo0U67uQgGx2v4rSWteUB+mB9zi519xNFyPvdIa9kRcdyHOp
sbVwNDXmGrAln1j/G7cAySgEzE2qtD+em5CHHb0adgZSiYcBzowKMDghfHo2
Ddt8qeShQk6h7ixeiTxkCwxq8U+k/3iVPqpKJMWal3XdK7/TGRQX5hptJ14a
V4CrwT6Xg3ga3KsZJ/lbUKkGW6IY978xdDm8JYdYZfR9jwcDzyyerl2Xz/ql
3UK4miWC/ZkQMiDy6yqnrLz+BGHiKLmmAySzOMHKj3t6rPz3c53cWiTOsc9O
zJiLaRjmCb3l7uiwVUMqA36JU0hv/YKJLg+pMfgsmy850mjGnC2auReCB0aD
x5HYsIyTRn1Qo2s2spf4Z0PlUPtkNXDKKJPA247Y1HEHrPyqfOZiCngYNWy7
rK7hRlmxp16B43Lek1wqtm2WSxwqQQkZ0H1PKUmNIDUIQpchcUsUFoh/UXuA
wjP4OXvLscKqSkSUx6o0JH6Nt8F4lOP4kehF2QlZ4CGAv+hQBpcgos01iILJ
MFQ+iRQONT/4b/g9dQLx7xsdxGTBDTrXTU9dl9D6tRTUZStiF3gC7bpE0kvB
ESVCmcxcTZBgDSXao9XdC7Ggt5VIW2/nIx7XaDM/hgK3PiiQmNOZCX28YFRy
3vj60M7Xi1V61wuiWUVOe7OnaqiYSO5/1JcjyRxbh4hy9pnFiuttBuQde7G4
6+l63c9QgMDiXqtvCpuMd9tHNq+h0rXobbP9nu4Ftlwy2jzHscdKIZ5D90WL
z5Xkc+nY8cF/uO/BRtEsxomekyY2jnIR8etyzR+NQyDohZim2UaCHq2Dxqw+
SCo7rCtzg+MbcS9QSbS5pCh1TmJqPvPqcUqgf97hQd4R9rzRcYbaM3tJiuDy
fXCx+YCdxlUMm056D0HqYwHbgP0/eJraxXRV8vDCxvlmf3gpcaZ1nLE34fNN
hx6wOslCYOMN2wwveFWnvwH1XFGVPm13SvSpQUpu5nuBbYjJkban89424UXG
vz7oKHnV/IvHm7cGvz7iQpUaxFh+II6IoyfLy9On/TM3tGEYh9TaLDDH7+jB
7OdV4sMm8XxDEtpqk4aI0RWl2Hn8xFT8wVuDxh8nxhzZak69uZw9OvMTgdSP
azolMIS+XCWg0zoqjzSz9vyJzvFZvuiiyPeW9gQQGm39RiN/LeRITFi70dxj
qJ75UUiiv+1OW8XNlz2XdSY7TP8SFXhj0OsSAkBRPOAvyOjnz6M3KqkyMwA3
B/iyBYemLymCVCZHqaETU5cca1dZksA7QNNCX2m2XX5jDOcf7EgUo5Fz0p4Q
3Gfi2OM5Lwj5/PNXaMAwu0jbCVj1mQvgOdxiNURQnViZkzMiIlzK8dLdW2DD
oztiduJcowz6l88jMthkBECW91umYmFB3AUuZ5yJ/j30BOZ0REkccweExL8N
zXxsO6faxzRQChpsisMSgr/pH+WrEmoo5jO7edTIqfqZQwa6TPSEtEFfWeJS
yqGWgYAnBLtR+2NTJMtNqVGBkornKn5IjRsDabo4t4Vzksd9jw/SaNX1gJxX
Lbnu4ufu8zVAsk7SF5MbyYNw1+eQmyn7JDpP6vV00KBL47ds0aWOtmizxexZ
UiAOSkyQf+y3jv3e5PdcwIADucJAn4wr1t6HctGE0l10DyFKVamAjpI0JVw3
ccyGKyVW1hpqegr8sFkfHY5N3RQtnZ5WBy0u77j6PzEWlEntJaTC5CaqAmHs
eqYOSBuYZEyq6eun1+hEGWBclfwaqvT5jfKv0FX/jZ5U9xHJ+K9f18Ej8UnZ
f1HHoBfNXsb8h03SDcw/bzegS+UxLgG0W7SqCgBkNEHFGgbvNJQiVSdEeKi0
7oc8QPo2RL9rh9fGT1/A1LLQso8d/xyRDAEzzYjcg3VgxMeZcJ8xu2HTHibt
1Q/4dj7whQDMFKtlugRumTE8wfJJ+krR9w1fB7RKLRZV7nCHgzTlzdVGyNHR
AUnp9fIVFLniI7cq07C5JtpOqDQq0MWMriBVFLSPLxyWrr0yvovVqe21Mgj4
2wgOVQRljkN6SLkJVuUBdtyxLF+7XTId44s5jfKW31cYeKJwP4j+AjM4Oq20
0OKOvKS4mxaULV/y/YsUUKLRCkTuTqd3sXfprQIuteoVFmrWI1iIeR9jjoPB
YVIWE9HBPZIAfkQ8YXUGVt0Scg2+tmA46JeXe634YSSkJvhIBzi0LEKmbXin
7GtTShOICwKXIM4Q5uMJqUTKwTP3VR0s3LuSYAPgtgpOWwzt5FXC43YuenMM
k0mgLwPoGTPZRx9wX2wwBvEI7jFga+eluw8nOEq0kf1UEeMUb9PB9/D1ChZk
qqdUCgj6ayo9MOL5zpkKLHgUxpDHn0UyafhVljqvLwUra//tA8tV38ah5Aqj
sJqg1HDNfm3k2SaMHaJb4p3WhhOOjTs3AkvuNEEvdXwqNa7mIfYuUB4NFOI+
ayM5FROzZ/1lAjo1DH5fZ0khknSOLPum4PsLJY9O60Ipy/cZMnLFU6FZotN4
xw2mUdpcHJE4sXzpg8mnrRkqN3XSELAwDkelPEHvTcSSJBHE0RbK3dA1XHPv
hBDuUIzzo1bQKscOXTKrGWERGST9JzraTzxABK/qWVEdRbMMd7bdAVsg/Ehq
cCpdNRkJ2rrpdgn1aLtqc6JrG5ELW7JwOrEQkyCeEdcLRyWojDq6zo2gaHKi
B4Y8ppylPa/ptlrvdi8wGdFiV8BcigzWJB2r1iERXKxzvmTicLgX9iJ+UAps
n9TSk6NeuW75ZgmII4X5AWG6j//mttsd2cSvbjGSBIUaejCh/mpZe/I+wWv0
AuQnp3+HHvNZI0ifeN4RX1Rr+fWzkIVQIVVOm7NJCHzTftehAdKBjGBCPl06
Ijl3rJuXsDgpA/KLggjw6t7DnhmJcfzqYC29DTMX1IsuaamwcwzBonkluww+
+4UWydSWYYwnFpDytvUxB6xd61GE5PF9bgz9q2A5YFt5/8I7jTUvIdhTLnHm
uEnDiMCqGJOi9HF69DT59CM9IDe4u6zT2qvG44At49HZQiHqvSvUrOWN+Onf
+Q1JPr6XFx/CwU6SF3S5iYwSRncDDTbl0QPrEpF0QUflhYqBasvgAD9w8XYU
Zay9RIdRBKYpVAe/ti1LbrR7BqcEM3VTcWY+RN7CjyF0d3gUSwhhPHe06aqC
391zquCV/B+GWUYNzkEFNfzVA8sjr3eBlHontTXttnmYIXTEjb0J0vORg2F2
pzUBn21TkUogOocBycVT60DwYbB9DM3vy4Cyg8tWcb3so1UjZiiMaiHndB32
rC+TajpJKkhOcALT6VtCGXs7h+yzpNiK8sUdpArAqUmUBbUH7423pjjnnAF5
7bTq+4LWdAXk3lzh04wot+JLV92sG9nerELgTQgb3Ye4mHhmtg+pq7noQI8u
JlGKhguTv60BhgSojY4L0n39fNsg+Y2Hyzx4QHrAZo/km6lduze4VJNdlSs5
azgyeTtROH3j5gjaS5gKLQfwye0W6Q7oLTmxjONZD/2tbQawSRy/SOhfjabg
3mj/KsENNxExiQIyV5tS1wE+gB1Gr4bxYv4IiqUDb+3H9vC4+sMZXdnkxFKZ
oxBCKnJxsDnQiLuqRpH7RKaHp2DcPjWX6dAAP/f9LwCob76Q3FihybOKlZbt
Y7VuoOeTBRYJBnuutCPVGxdTJPE2pQ+hyU5NZt7mRdmtYmP1his4y1FVRsME
TXek5Y7Dhx8h5C5PbqWsWzDxLIEhD+TgC8bNGJXiFyVLBimNsc8zfZu8riYZ
9rXoBgtAUfqc0szaDT6FDu5z13EM18ZIn2k6fuosJUO7qJjPD2u1eSv1+2ra
2YMiimjUZCGlqPxXBvBNISoTFrPuralYuS/nz0NGhlXwbjbIhWyX7+42MuA3
5R2ftv7dQ+hPkSlJRkCgyXfPLOLeUmRXVmgTyo4z+ctMyzUez6cNnfInK+yZ
ds+KvfeBteEU459Xt3A3UDHS8WFGaJlv6m8PPCkle5Zy1NVrY6Xw2ffqRO12
Z48QB4BBEVeN4K9SfzGvaqDZ8Tpa6Pteuxx9ctFZoe10WmfVCoCHS3NXSEKw
GkPRcSFMd9pDS8xuk0rzg4hQYb9UtnpysuysQ8zuPC5RpBlHVvWjXjp9uYez
lN6PJ0wJGLTgpmvjrYR6m75sU2exUVL10ayNTn8tAa8SrbrjLaclkWTF50oU
Iu9l8HiIQDBd1Ov/ghiFzyyLR/t+semZBSBlsKpZH2dbb5rwRapcwImCbX86
u+20SZuW6g9CFqO61VbVOQmmP5fYvrwaSeKys9Jf5EJ4qNoO7JPzkfuvinF+
dffdLfh5PLvfCFAJDPu8njs/2Gtr752AFrQYlJ71jtezMlt2yxtfFtLp/ZaJ
kBex5HIXAx/zyICVdLNCiFsEJFFROArOKSz0N4Ik0q6N/hcTnKu4VeCYyt5W
yrURQ8aOxRkwJYIjO1S1MISdUymX+fPcFQnJ/N3cTnJoCk1mthGWdM83dAhy
BMLFWcV9/nwkt47VXcRmuzmJZe2T02AVKWvU+Nv5vUqnBO3AsFnIko5PhM5G
YF/8mjVnzQKjsQMuUfSOE2PDttkRbN55eAxBXKhBdPkT1xd49d6QiEWgpfk7
AyrThCrMvpHp0EA+OVk5+Qsss+vcOXkOTc4b48m489StMxgqREZBeaR2+vSU
Z2+SFKSpDMRcmzLpLqGgMSJNNHSaLcADhnRel1MVP3z+br+6CbbM/nqVVaYj
oHChBQ9oLaHB93oNNuFGA4FB4+VMaVdfbvOpQgevV2I/cgwc//qwWzcc8fxc
bu9BZf5dZevVKv2he81u/nnWmmBgS088awee87Sb5bIOFn0Wy2ZbuvFSFl7I
QPL9e9XYMEPOMy5eYBprotuQN9F7BQhs8LO2VftEN5yWAn4iBQ/rXcOjcjQ6
1k9QWmX/I0MvT3PuBFhQ7sHcjjOR3TDw+MVBeuc+uVhQOvdd1AfCsMawfCP8
RspMbW3WXTbSpeebY09XuuzSpnC5XMXWpnpd8OEGT8nO+5Q7+cVx6xOpdwmM
QXpd7Isd5IyHer152DAP6Yt9DRbRN9q7/7a8yL7vMgIQwXo4k5pprH65WO0G
FroIXiJzFJ7Yo9qgxcF7sLPAoNGqToT1ixDWyMILy3TzQ9VjXf3GV+j37+sR
6OmwBYfsrP4Ky6Utc3+6vjrbaXUaRWuxUWlh3oPIv5JKsEx4FQiJ4bjlp32F
45yHrsqRdpUv8eO0/TPtoTlBV598b0iijBekdH+CuO5wM0AEVUxndjetYzDV
2bbbBZDFW1taMaO4CGDsJZQK16IfxeOwumwp+a+OEWpookAIhiiOw8IgQQN4
U1kaq0KX6vNV4/5rMtxCXD20aiQHAsp1QpPFjiFvyC+sEiq9N5hkVGVMMBz9
Wp76EQgYpu1fgm2s4PLc2TLDleGdCKz1lUzdniSp3EVkBT8fihIrCvhg0TkI
PsPNupHcf1Gkn7QTRAAtGH5oB7MCrYWwebj+j8t6vQ+ay741fENgEcmiK4Mr
FZG3oE85w+32pNAswNeVYixxiPZywjL3f9UuHP1X+BQkRR7PebHsnJ+gpEV8
7FvC+PC85SLyrN+9sDaJC63SmO97hNYxVD7evFh09mvBBsD2wHKPllOwubkA
Rg85qEbHXGeqeme5ybkwHNiVETepU0SX0QkbxAWi4iTaTyLDh2vbTrN/TkpD
pSZTxpp0ODbYRI313WwwhhThAQoBob8P15AaQaoJzYfnSsDg5J1R2axzdWNm
7a4YUBE1pc0uFJAmBMXlrQLo8zy99InBki+s0bPFQ4oDBozUxDlGuE7xuaXH
nuyQloDTuL/8bMjVQcNPSFX98NKTPaK+p2ASl8pDOgnObgEl1GoDG7KX1x3k
8L/uQpWpTxYsJn5x852j6gYtWp87uX0BdalkZ99L0V3qfhOQgy0v/SBNCh8a
kpT4RG7G1pEJeVjnY/0OoK0PXpzuX98zepdGQwemhrp+e3ZdqzlLZpm7T22v
J7Kxzsm4BnLKtLFfYZOTXihJ+RIOWtnbpBL+yA5Af+LFIwCn1w5SQruhKRyt
3xEFK3anrEPAehBwuMwHAJbXEscg+u46SMmJ1AD1AgPgpDPbh5uYktPoirI4
C9BNh7q/FwzvnQGr3Ts/f+SsTRljR6Afu0ccACNzqpatAh7nurWXUSkfWMiG
Jq7E3qb/IOLghTFCVJfYPk4ZYi8ycVZCvhRcOPpKGzKifr72GhZxRp265kGb
MFiQTHxb4pPQyZSNBi1xxms5q83QGPgLBTiu3cPH7e2hauCJyRAAt/VMQ+e2
cpmheD8YBNPaOAC6MVGrG26PcIFQLL615dmwXKGOfTJA52giR4Bg62k9vmZy
dF07wHfpovjEqs3zdwSwmZ9xYRBrsJhsO07K/YncMvV7tIGLFOcgTTK8tcGw
+Ne2FLlIVbWqvb4uPsYWUHHlQtu+S5UGAdrOBlVlwcFGeFM7KHL6WyqtLxJV
TtTqhSo5TLuTfcV54CYck3wh66jjK5juVCuSVUhQlczGhycKGyJwfmYdnkFn
RxDKt33wX7nIprHrYnzt5qnc/2OZD1JvMGQzVsoSxpNwdoNNR73nhCIg/M8N
bYffP3liMQA5YLg1oMa40pA7pXfxSNmbfrdk552y70NqE4GlMApUw7vRLaVF
SBKHr76E++vUzj+gfDqixrtivYDQnkADN4w0xhmxL67HZotgPBe1shgD+idF
DvD9izAhDFHGKoD3BP7ch4JvbZYyY4JeYlMIlaCXTV39pNg4vVAL0dprqraq
tJQn+3jOTzov4dri7yMwYKgRO3BkZq7MMmJuJtgyxzrNnI030pJyz1tUCIgk
f//7tbYppPGrsXfYAownDFYfQJKqE7HYyJ4pQpN4gI4TCeLHlbk185JZpfj0
iUBw/TrqRySZYDosQzdlDdEyM9EoL+eSUNFFhu2W+xdwS8V3RvGvt7cbw/6/
g9upnQY3aGAJrocNgqdrQLLbAlGyXC8RGOayhNMHaUOPvZfWnZEP6dDcdlaL
jwB0biMod6hDO70XIFv1wNkHT7G3ErqkVhglotFZxSzeYWLWa9cxYBU3YD/W
lp64xBindE9P0qlqJtCBnPPmwEbRb7glYrv1lQux2uwkaCRVA90KXGf5VkiV
hrmmHFqGDsTIraHrBmGl5DwIE7IVS9kqH08Sxa8mx3ag3FOPulHx1PIRrvlI
LnVIbTdLTQ8OScdtl+veQF5mMw4GbOmzrBcTMuP3ep1Ld0tk0qQntDEYxz8z
Gz7kFgy4SPnD5Cy01pU81Fl7HLqCqXaSezno0n5M70i3FSvuU7GJG/TarmBm
AWv+RsI/3pXmpteSiI0mDBc1YaKEyWZVOTKRc9ZFqoyl8r+YqEInxA8A+Oz0
Uqsj0u1byuH2kcJyfvx4QbUKy6neYddQYDbSCLpH6kQCrlkNYVscPHKq0Z8D
8chwNbWdZXnlNyywl63s3gbmn+gCZ88oc2i2WmFaJ+/6xp2+Cyt+PirbAhte
7S1C/ww+Rye8ngN1WE3PTHN9z319nnuew9zSywgkk+iF/p/wzNiSqFBTqG99
gj1Da8MLWgi51vX8uDGfb08Cm4595NKITFrHLuOUFGGA3IflxqBrmEL2X0Ep
SifmwHk2bIl7Pmsj09hYpyJh3sivoEvJ3zEKV30LSyyE7T9Q5Anwem4zPGTB
mxdkwKGWLChbN0YupwVcMdLV58zzatdMtDKcsuJHeJqfQ0Ay3cct1oXHrYSx
fR3m4+IZh+T6rBfSX6rRAj01RCmrvis8Nz+G8lqCMQfsQY/HdKJgsof7XnCK
nuP58tVjcqRDtuDTxwcQDKza/ev8nAOqY8u41D2yvUVdsRU1oWvfuylB87s8
uNbgmdXpKUIAnDD782Q4fN0fASsYIWsLf/YrR3hCRMakl0mjfAqKyXiJ7gzE
1oNSnaWDMF4YjYT80eDuMpCb8RAI9eEGfCaSXoPa6K2wQTLooFETJs6tuDFV
wYfY2JSi7cDoZhb9AIE0nwwzhVGMq524mReXkuw6mGztwgdR813DMjegVtjS
en6R3eeFwpRmZl6aUVm2n7jQ3X3pMcjV7E0pNPk3J0RN5XkGXq4gsPbO2pBF
Otr2G2A9VACzUdCYdXkBBY0Dh+FbWUjJW5YYn7m9DbSnljz/ZIhZz2UBUn5e
XZGVCsZcd7K/AvUvU+5DDCSg8Xi6DccTOOQBHBhJiaWGmDlOA6snl42OR61T
N3hGwiZzF36WJjOa0TE9s6OT597lez3sbjNN4Sc7y8IxrijkQVf+sOtl8GKQ
4FUNowEY6l5zQZklZi+p6Jv/rryg0mwdjAcXlBGmSoURELRZMf5c4fRGHHsz
dcDc66stXrLK33otiv3gVrpuT3LhHrUuugVfWsVQ9E+UYjQ2oH3yodA0fBER
bYEiMvFSbBo/L2Yv7fuqoLPRpI/C8tYZY6CaQnSBrCJYAMizFeFgUhojHiZq
2zEfr8vz6zoVOrvbb8TtMXBb6wCGJOeL6vIuM3WM1vN97+XoRz74xdDcwIOQ
sQZRgDGcFFb9dKZNS+9AlkRBsEc7D4Lb4ugnCXJPthyOXwI/8cClwnd75zlh
v10+o5fCh0GP0gYR9m4UVyDI8Rs1sXpQOKRoJvuRDKjXHRch/zglTznNbmK4
iedPll85xbWSoj/KhPhilqtc8VccAQbjNwE8I0mNEDiRvKxNvZECtTvI+hhF
xGk40j7Twy1m6Q/84bA8brL/4VCO8NU0ir4h+fRkIKYUp3GQqmoaGNxwX3nN
QLYI9lhsv3Q0hbCBQBjV/R8VEEA1ojvtS8IASN50hg6URekKdlez/OZCXVVW
Qqyvf/Fe5Fo2xndmnqQjDXbSCNuf3l22jWf61oR1xozuDgzXOmlAGR9p7ygI
8cFSrg/3fh/m0MtxUjvFhauR9tJST+i+s2NXZCCTbhgbFxvoVdCvSwoKxD/m
BpgUAwfIL1KXoV/41fuVjWSIXQAAFaxVjFF3aqk6HIS9RZJa/7pjhscamNbZ
m6JyBnk1hv9yOe5E6SHv+LjZ1KbUgfdyZBtac2wpxIF8cXNm153rN5fZNTxs
UZBolbSQ39g/cCeya0XyXQOW5VIS/jcWfJCVuOt5dhLt8H7CJ2wLdSNzcgU5
fV1AOUlS0nd+yV0dCJxSC+lhazL1HG/1lERjRRkkrH/zpeD3pwPgUv9WT0oZ
gDwhwpekdvosTqkjYWY835px3fROFEkY0UMln+UZaz0cjCjg8YlTc6U2Gjkg
SCxUrPYoOVXQoUCPacxav2mtB/eDyY4/0XYJqktzp3t1wCvsqq3CUDOdegbA
oRtCZNhgaHoQLdaeL/RFqjG3CHEcvDh9TSxGeYJvp7rl7ghB9V1SMjKuwgJR
aRS7yCx5mKaTTbdsyr0Y7i4w5T1g78v/LiwMB8U8/cwt7Lfw20s11+Xbikky
4mAcvmXt9pQED4GdfaLub9JiDDkiy9lJ43hGQyHHfxGr2hLpSOeUDuy/mf0r
Lzgipgbv152Ute17nWlaAAg19JCELENBLLpkLpTYKnhDY6zb2NgfMSNZSMAq
OFHzahBfzXRxugnT0+UR+1iOchfs1Lc4T0tIuZ1T/XEAwh1ObDWuJrZR0Tjy
P1/IGsXeq07BQipR9m9S1IVr05uspaV0GpLiyH82vWOmqHmDp90fv6G/cnSo
nEGXsmQ/AAeg1GuQYsPmSPpFkXuSol7VAa5qZmPO21+GvzNg7Xmr9MH7DxVg
sqJs6WD+SB00ZWSqlvk866JtHulJXEXVqh512y1w5IH4gKpihSwQgN8a/Vxa
3TNeRH3ONk63/FxajFQ2Phf4ofPnS9OpFIzUBzoaMaS3CKA/8bXo1cVZO8O4
a4Zt5lTkFZz8saqExF+fHXCgGzRfnWwLr7dvFm0DRh6aYy1yKCyMXrW+9gIW
NKI4bryolG+SMQGn7WAeBgylSPRgjs9WMko2hnGfGWBJHyIpjTU2BLlKmBKR
kiO2ZTZFnpgyHMKxAcg3Hmze+wBq9juoRpl8HqRKxmz+meWne2Kwmidmps38
jSjaVpnXlSnRmv+EsoCSOI2hbbAUCtRZD4+Ih00fyxP3JB1SiHMXuWzaBvKj
6dIQt7lfOChXate/6C99U2ZxkH4RngXHe2o1HmEFt6maq74xEGiWC61HvOVB
E5ghzMd9DK8zjoo1t8A3edcKKvXru9NOerVuNcu66XHYNtFf+1iwJNXLtfoL
RHfuZRGVxkhJiHc7MUkCNsSX6aRUJUDapVzj3qFUwxsyqlfMxBnJW35dCP2x
IzuaeKS6R1OEKxA+F9SuiU8K1VJa+9T+elFno/UoWAHMT3FEzdccwe/fqIW3
nWie+A8uWv7zUrUd3vF34gHzpH7dKkp2tpPZ22UR4DxBt2dKys8tz0v6kp8w
hoM9ikDMdywXcKJo94Tul1BLo4csTwS7l4Y5RHOLtpR0CgthWEMmzWleBx8A
GvT6JkmK5FE44GeWmBj2Anud8D0YinrbrigzpXaqlEFqYWtvbosMZrbPdD97
yPJ0GMvGRbOthn87EWXsTVfh3oeVarX7tfFsrdFSlJS4MVBxWF3P1WGsi7Ef
9/cOQoi5bk3l7ELmNQixBFNUQw767/v4cP6GC7Fbpo2MWe0xu2B+vPUxDQFS
und9Iu/nwb5iRLDCcYVVu5EgbLo242te9LPygWzQwuJB2o/JQn9hkl1vP/y7
YJR+lDcSz6pPCT3RAJVKpWbLWVZAGD4mX/qGrGfofk4u8FKB0XoG4XptNW/o
CehSdowgclbE8Dt/5VDuY4Ew5MkQS0TAiQtp01HBTN8ynGa++aGEyfDQFrxB
ZPxb8wbOvS446Dgrs14nqfiZXOLVabPtWMylvpsDVBLjpA7wLdOkVzWA7m8L
RCwBQ1EkmMCchmiSeRaLpBe585NOam5RWRv0wfnsGeBguNsE9Q4/iIZo0sFI
GO6jbfwGOAcOXGN+qGkKUEkyvxxEaf36tqBKM8cNB0b6ZQmiLR2EtUcH0JvC
ZSkfIHxxF34/jvSX5iiL7iurAPiiqaSpe/sGYGm4eqfzFSDiqCLZUCUGeC/1
vTAzUTggh8Csxlu/wdRXBE//2loj+S9UunuI/JAfDbLULKd4YpZ/xdtU9T0P
wS5YcQlWDX522paBXqQMzgM+ViD2RYgYf6UTpf36r7wM0q0FC3FwJbKEQwWI
ZF7xtlUc7ec09WCC9NsJC5ujYW1DhUeSamZKrZinKe8+g0jp7zShkCPLHF3o
yKTnf/GW/Db2Betkr2HKDqVH5ea7a80fQoIPudWirELG8Ra5ucX2R9PSP7GS
E4qgSVX3OaA/5Vrc9r56AnByV/b6fcXdq4pnQVVgR9VKfI1EoFzVjXszNsfG
F5fzNy2ZKo0bJS0r+hzKU9vpJINdAbjkv77BU1oVCVN40ZpxNOIyT3uu/xLY
/2xC3/HkzE/m/s/+1SPbS0vATDTMe2aJmzLyp5L2uxEASErPVhEafuKitkle
bAuS0znOhJ9JI3z1Ehh730FuQFhCuf2rVgljno8ChhpzpaKkswDmGMVm6qM4
0rFXf+537pm9hSuLicMwXsKFDwDU+GlCBCThiyGegd2oQigONCI0uXkTM1Dy
2/7pP7f8Tv15sC2ABq2IgsqVhfdnV6eJ9BH9qDfwgT4ZcNIxH5j7zOIjsCwy
Z5sLo5JE6VS+126uCzGdfthW3UPtH7ALdElDxMGw7fomJ0qZ0Sw6VZhRjoMv
LMMi+iKLUB8HI94SfwXxCIVSaJWOvZBEJPJu8K+HRGBaS69hN9vCu9uPH52Y
GcuthT+qtK00ok4JASJ+7qpGOfGyjEBvL83j4TooshT1SrQhD2jZaPEmb3In
SEm4O2Ajr/vhUTE4wKoFo4uHXtWF25Ebky8Z2/TvV6EaiJTQxjaXs3OaG2C1
ORHGhudmxQoDFoLqIxv+HPhbYdgITGw3Zwcjk/PJHYqniWPbFG/GGFR1cwzE
G2A8h7Wx0+nm0Yev8ci5FGZu2V+mpVMJlqRhhcGywpQc2VPJZzkKH7B14ejy
5ic7sxF7JFDYWY8k3lMBG1eHsdXfvzeoL1hlFy5sTw2V71jIxur2usBJeh2i
RIx+zrbAUIeTcbyGHBtHsSSA6t1RSxwF3IkO9GGLMBln89DPBgQr4EMv3l9P
NftatlHVnlPx6nca6/YpEmsx3369xDQwNiFllz3+btxWMJJvGX0k/gb1LE2y
e9LipGTYWfF4MmBZagDygtFaAjc7yaCDiRZoLAw1lgP1ZYB8EMzM9aWbW0ZX
1ad2v3IPjJ1J/CXu05HePyp7S30PEcFKHgUbaHZVvMedVozYJJo6C/iqZC5I
nqe6vN+TJa2ZY38/7Qxh8XapsN6nJDlL8X2BHMvGcPdDJ1t+f591wVDVpE0r
5jFA9643If4mZloSsZb1CvjJVbkpMO/fU+/4jMoVF6MMacpfGWguwlLi6eNA
Ka39h5hebp52x23U9A83cxULBljY8Lb3eUqoYHPLK0abxmGd/aEbDcBeUu1i
NScPCP+LZ5YvPicy6CEHAkz9u+eZ/F3MQ+AtwytnDXbbCQP+y55mGAiI8Jox
HXAVAVCMZ1UwrqE3A3+KTjM5RYRhkSeKuMSp0aAUJjTqqXeguU7UmAMkuZiB
tP6gJRU5nUdYMH8w8Lxl1ZdaXfOvNPyyVQWeqI8US/IIHLQhsya8o/Hfjqjv
BX/0TPyO5Om4HzJ7BGhy7IqDTnTT59HInnabpJp4Q8z1g7g1bxzMdzILngUk
IHRgXgXEhAs5tBzW88DTKneo1ddlDJntcTDl1qUtSfZqk/ykTiIrHF0FxznU
JBVknc+mFqKiWeRRpSt1aU6XoKkTJe7UE/a/cSf5oF/Wnyk6KFE1EsPzcfxn
hZGc9j7FHbRJNva2akPA7k9KMVadhqNO5QZUyu5LrTDTXcwU5wrld58piaOS
42O30HFoeaxuH4T4WESsDHjwteSL0k8jlGo+jmBWYjUYLD/fe03VAVQ13obH
3KPShlWZVJd9Zpiquhzkz2eYQss0gnZ1qUqMTaoMi/m1Rkcml5+nq/jJGfXN
orWy6ihFzESMV4fwwo94lly6YmfSfNsnF206mG7P9biBWykuD8erELvy5sIm
LvJ7J+r0LrB3b4b61RG/p7dv/Oj9ciDB0Zi7QqasK+C07c2+3xKgSQZFMRQ6
PMIP2sMf1v4GlMWWLhZIjGsvVBg2FYjWkoP4tx+H2ZJiyRetgX4wkBZwz5kH
VXpAZe4JlFWA4jEqS4myCgcfFB7uqR+deURstwK/m+/YgGHCtMGQR/AWQ/rS
zoa48YttF2LJSRh++fXRP3CYy+NX1grAAMuZR55dFhlIfu4ugv1mT6kzEDVl
AlvKdTdlDFIn6B2xS3/8wdBy/fAAbsLUtcYwGELorqMyCo80XTErOqkK29Q+
jm/sUW1+xllSuoRhOpMZ623eVH99j1DLL6dAdMCta5CRS/g1ISKRDw8vCuXJ
g/WSyEZEWDVATtl07E+N6Ke13+lvUW2eeLBruz4avJffRqAC+3jIAbKQIXOe
/bEEAlI1f6GI+lrNVqOS9NpmUTgiFmnsS8mFsYsM8AlEjMRjj9EXbF9yZ0Rl
kPD/U/jshj7KerhkyAZ91fSjTm3Tuv9VohdxXwoSDkOcuRseu7oYW9wtwe0/
/vVsvUGkzaaHbNhvNoVqzybcTD22DKvtPgLTfNunILKwkkmcSpF6WVL+Shk5
T4nsrwUNIkNiwluanv7ehceV903+gbffsiISLaM9Xc0wRMr6Kw7q4ae4Jh0k
p/n9WXElhwWKYzE8ioDNsvzRvzel551k4jCfZt4H/RvFfrVS8iV7xPf7a4O/
iZZHjOIUBr6oaXPTrLLCiLfIt1aEFXUeIhDAwDM/hyUU9E+YQggAGH8XN1fP
CIr5m8iM5fxnxh+yS2nNzjoYWGkIRlw5cP9Q3ObZvqmRDn74lR7Go1fOXkPi
0eP/cDRfOXnkNQ3SEU9ei4KfGfGR58jVbIJAggyCBAY1pg3WBOZ3JnAoyEOU
jG+5l6tDO1iqNbj2BfhFH7n3CnsNyaRHe17Xuyl1oAgRf1emj8uaPyY9bwZA
L5To420bIca6okVQyXXNFnNbZIj3lg1EPEB+LxJJicaG0gq1epA2g8fi09wS
W3LjCmwDBUwLwqeiECCzhQCO/ZBbrIPJWpSfCJG5GFew3kYTfGI1F8v/x+dP
8bV82M6u+hK9eXIXzFHsTmDUMRHAUJcZ0b2KyyoN02l9eih8juwfsu1gQFG2
Cvi0zrLznBkzjCKcW00sntVDnYQ51YSStfwUiivphrsXKlBUSvhsbMFmbAVB
SO3xIfq+G8/Lyd3l5IFFoeqEXzbQIOj3pHJT4gzoVkjU9SGm4PU9MYtmLXMQ
24mvr55dFQGdVN7XEDpl5ylB/+KAGXqmLZNoDoIOx9IvD33nhAG4DsMsUTxG
LMoRmcXYbo3JxDgvF5IbhgjWATOLpW4KfEsFYidxLaY90Rk6Mkxu8WMs/hFW
PZ6Cb4pS0prtnonQXPCf8h5Az+BB1l9hS2dcxeUxHg6z7twDfRbNrnC3wh2g
cR0tFVR6P7EeTQLi1d+vrqotrUTxUFmzZ/LYYWnw9Wd1gjkfhBh3lbXfCYtC
+h9YfI4ObGhQYA/esfv0GNCGlLJ5duTt7bIuDwmdJAU+bcMnA4wwi9yo2FCJ
aoW/EoFm88I77knrhN2NCRp/DA5T+uvBYJzpT1ubMuCyTIyh+YNzTNEUjufn
wAz1xEhi03EPS/cL7siOjwMVQmcH546tPwlrBP38fbvsCbfX9+GGpo0v5XN7
YWSsWbi/ZAXPC3CnBkHOMXnJB3GT4Bql77q8WgkmhRBdoFgfPyMU9faV7O2/
+/4Co+XZxzmQYKDIHIqGUAiWjw8fRnPGYVYJXuO/ZSZHo3sjuiZ8gn2NtB32
zdUZQHvWO11qjIfkzzfEZf2LFMwwd8acI5L9ZPjHLEtJRO6CVmRjox2mt9jE
iB675IAVKJZxf1CoLT4gxI3xZIu/X+xrC8rJ8L6u/BkMn218bTJXT2l+GanG
sJkF30CCR8rDvBr+LC8hZ4kzhHaNBrls1dgtB98yZD23RkegFImXIM2N2ADY
ajWPAsxRIzSVxYYbM9sLRpvT3EAhcP2cCNOGVOYAFQQd7FsmhYJERklEv4av
vbnLJFTZfRBeF5fAkSvlOJCXdiwR5MYDo6QZ3qELsL1wd7DWRtm7GXKRu9A5
xzgh+bbzspAgGt6nB9Gv+FGolk8ukG3WOkBSz87P7eb2uERbZsMKKA4s51pf
IMtkM+fB/ejuLT9kBlN+BF7Y/VS6sWdNy0l/F90WJ6UwE7iXgUPGSe2njQdT
gv6acfLAh0PPfxng0HJhDR5HEnP81PLj+natCG6yhsc+dmzfMjJlHSr2I3y/
QzczdYIo/CAlFEAM7CPjRxrstXDsgO0EktYjhlfelTypw6jRZdnAiBXSmv86
Juctre2rgs7clT2cxxujRtO2rHxwK+58IyC+zYNkhn2EadHTRI56xT444Ojd
9iv/9Onf4ONGd0Tsqq+TbfjsgQG+cdXy/wxAGLonxfg5vGwMYsYs8GtdPbIG
Weg2IVErAr9tUnPwCZsrYI4aHcZzWzuX5QA6kHrwQpsQzrIIBZQNvxmnfeo6
r6FNCBpNDi8kW7YxEvbUlY0FpcOCne8Owz9zqZkJFajdLIuoCtBQCQUJAaiF
5t3V11oTgrB1JL47HvbSj5DtYQQzasTVUTlbH6c3owX365wRWp06Vop9y2BQ
Oos1EXVQ6VREzKAnwG4+CSC4WQ1B0WD2leB4YdF50wy4t8JWtVsT29+dp/32
cQety5ene2f2xFCjHLkEtP8IEaYtsTX7qpUqNF8g73PzsuxP89diGcLal1to
w3goLTc4Je6KIXLLK7GcW4/aFOqNg62bNEBDtaUKZaKlEdt5fbu+7bEuP9eX
kn8MZYqWkBa93+rKVFXt15yzDSvjx3iALwYVh3bd5maemSF05Larrm6990Qu
wTdrakdDvsILdl6jF28LzmBuN3925HGkV5Hztqo2IL0S2faR/3SmIK53tsU1
++GV+3syNu3ODjBoTrFNnDKChyhpaTlJUVPJtebAE86tNkrbXFbn0cDY9iBY
8DOQuauUWyCcK4Rs+M3gfyuaaVvT9T56WnRswvRRFDaXmqqzy2Ib8eDeq7ZV
A4HPvykhldhTlS/Zn4I6Okqt9NxqfAZ7NA/4TCzCrnCA28VPN4hPCFs/kjCt
s7CgkjXEaQjH3gYGMh0d8c6ybE4Af64PtsBbx+9Ui0FecjgAiS8vMSq/2IxZ
wsrQrEe1uCdFSjzVDpVW3R1nQC6nR1YA9fn7rWJjCtDOfrwDiiu+pNsVWnT6
tyJ3vysiq7McwX1FIr8xCPAc2mwg+lNttXzCRJ4Skbp4CsiKA15CWVAZyOGy
Z4tUbn4LbjBDJDRZW5EMYYANei8QCmj4Q5dJtRDisc3nmYT7d6Dz6RYiKhQH
H0hRpDLjMzl0TtTZvonUJqUsy9+hujGdr0E/03gsZdPipj0k3IqTd0e/uKhg
1LbrROucJYA7xz1aeCw1aNNYQOEb4W/8Ga6QYUkaVZ1nDvWDQW1ldiO4Bwgd
JG3Zp6Z0DAjamj1ru6PgreyeryCSa3rHEF9Doe6bGZo0dHiJjNtwqES+VWYw
216XYLvWpRqI5XVEj8ezRL7lj1DDhJO2lxTaEU66XXyEu1ZQ+zGqQwfMKf9/
QrPHiOuCc86Lz7x4xHjQYDOtnSXaYi43+s/+10H65wXPjB9ZnHaoNsQiF3z7
0eZsZE7tMCIkIMoMf61rDJgw2+7yGOWyZsa/UIQusv4j7U6NMR7GfJTd0OkV
HBEYmjOAdyPJddSkpAhueR1cbWhUWmwPDD0Srl621BJ8sIqUso8Bkqx/LBj/
8EE5sjXbN30n7SyZwKIrpvDQvBKhGFneHWte95IZCajHpq5ZG61kLSxSZqo+
EHGCpo28Js4w8L3Coq5SVNeZT28XbvORSYcAWvGHz8YesxQ3w1UCCD2LxxUJ
XjSS4/xqAGCuODlv02zP7mA4ZMw2XJ7R9tNKhTxa5CZG5hnKoyVg6fLjcqn8
Eph4TNYahKZtRSKoqEfUu35pXjXKMOmdoXMQZWSS9GDYKmI50db0k6GTeM49
nXZE8n7xgLAY69DhPrX1pHMt2Uifz2qTCimVLPnco+gQd4M44hQePd5ZamBd
XuA9fo0Uag7xsQWLPkGX2iPrccCBG7nvp49SpsZwH1bE67VvEkWeuMrSc/6h
aq766NDvPGsIot4wgnXV6qpWlejaprNsweIOcDko7WpQTk79eKko6cZYrRyq
RK4xIRY8YxfpgPhHmEasR6zX33tU/lhHWxJrht9ott6ctKp/uM0TnDYcZRoS
dNGa5jp8Lh34SZvfcB3CFnIGseNnV5jFud2rRdX4ot2+jfzebzXf/v49/nO9
uGrq3KIY/aS3kcvvXhr+JeY5WodBp1qpT8X+UpB5/UDQ7Okou9Ux3xpIVwR1
pSoMnvEeUXm6dniTPEmZwwyJQagpop5Eo5lTi9gRqYdMWuGEhrDwOM5EI0MD
X0yNU4itnzYmGJaZiyM07gED+S8hRrHZAOZNEz0l6IaS2FPUsitwvYgPpxIQ
2SY+S3VEfIwD39ubz0bcCEtcL7aoHKSJtw9dwudJDQnCR5Z+vlIWBeLQYmYE
m0HJCwWjfeuiBKx2CerYsQ5XdVBfMMbiGjEXWfY9Dv67meTedgkiw426ceze
W9ccII55WXwkvv6yGHyISMToeWUd/q73xdnBt3EF1fUoAOqjoGe86gl1yY84
26fvkjbHaSFrulJFwgTXzEUf5MB79AVyyMLWxWXzCOlKCiAymiRcY4xLbAQm
0VBchvR2NhFMR104h5tQ6UDTsnCT86Rk9N7CWifPq2oUxUjJsxsgssEmI8Sa
gkLHEzdkDupM4S6H272Mdf1SMSnXX9enPuZJHtKa0REq/lO/oiOHT6eatbok
IK4QX4v5Ll2TK0jggoZXFrche1gkDzpnPzNjD2+a3PgQr1jyNNixOZRedtiw
OrP8qIcJvb+6heKELPb43CeUdBoTrxwGOqMZK8Y9vZ+sKl25CjjesKHPei94
OhEl5Iq0J6t7kXzR2pm7MuM+cyqJTXI1fduxP/DQHJPs292WoCoIWJIrXq5h
/2CL/jCbbzd2Ypw2kll1oorTyrBZiTIVSZc19F10olpIdV03RjANuCF1jDRl
viGkMmMEUR4IQBxg4jvPxjLVIX9K2Tx7Qpdg7fgvEWySr9XofTBLmAFryQB0
CwebGohJU3WF1OL967iGl2qWrnyBTGsUsC+IFy55uufPzJZTwGVP9JkvUdxx
AUM4DNulwtFKfVGkia89t+ULVsNOq51jYe/eJ68uR9YKmhI08KaRH5dvjTHv
Q0SKVQ8HTaIt7Iv6zaIyjB3CM2q0crrJU1Igu9ng3MF8kgz7vppARdyvs3gX
gfJ5udAX5oryenqjrdtQYmHMmO07CDo0Xfd55eCT6VKJ2QSbqMBTaZp807ms
6CqkAKeQiI9h6I2js6WgROF8a7fiRG8wvDx73HCsk9am+j0E3OyBoqnE3ZoX
ehv14djs9Sh6ySV3v78xU9p7yPboimsKLR/EGaXrSsgCaCWrYLwNNNmwyGAJ
bb7WdLXfRat8wC/L6ZJZxioPv9lbWfviacQI0g16Uc9VJ2m17T5XwVP/qsgy
jr30vYaYHwj4bmj1hqWKlHzcST98/mYbjfB5Quz50MJmEHaD5VCoysyOG4jY
DAzxLEB3YKMuhpCoVI8kmzI8yvg2vtVuzGrSR3jxFHW7sIvgIjVq7Ewwn1YZ
JTILebfftyVh5Yrn14wnYCZAuSWthf8H2qvFUhjKQSN9dbkqHJ9H51rYxsXD
TNjkd1oGvFHmVC+QIdVN5vV3uOoFO33wHQex8OaO5d7MQqtNxEZ/NMrVJcHP
df80H2Us/eTjS3wJ2MCsoFd7X7W5RUOzqVwKhFJdN4/Q7AVCY9exCC6jxXGe
FURCpcHtjj3yRJ9rfYbKPoo7RlBd8OpvFaR2LfHSW4FDAqlPKT//3QMHPZgK
sfz82ZE3cgcBPW8qGgTQo1JFsKvU4uUzJ6yPaqolpjXy0krr

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "B40jvh7ud/ahkCWXo8CJP0S9JYnc5+J2pwOdONjrEnmjRzb1YpxBEP/gM90XdEQFf8e+9j+GJABVN1VA/EUgHmy986oXHU6n9uJJjaeBsR8h22iSaiy//95eH4kKFakRZgkZDqWp0dX7AUTwRg4vZKk0rom9cx0xsiuc1Ki6fTzxDmmuuNW+yyxk/luKJogixDl7f05H1PhFx3JTfD9y6cRFGovJ+RtyYHOBbLpk0whfEKTCdnooYQ3F3IKUQO5KvydzcIC++Ym/jTwE8vGGaEFWGxf5ffl3hC8grTgVtHSSa5lvYMa/Epu9kAsHDsCLiX9YLu66y69+BSwtbMkJMnZQfz5M2Le8rpO5Hot0UmaPU8qZXDJxAhUQsqL5c+uzMDFqVvTDDY0K51pdaW+TIQjZXSC9gP/A186AF1SpfMVRfyFo3IoaHQa62RYZB6ZARzd2vd09uN3Sh7DOqgh20A7mAY5XSg6tnbKqMGBOOYBocinoRdC0qcNLJOoAmXlsw4pji+7drzlZYFCFVaDx3AThtYOLrycGPATwvoANZJBJ7mhLLILnZ6F9+PXXfLsZ0hG/ZomJ+VUG3ywMc7bDrKsertCEFpFHdaVJwBrc94T0ZE90zctl184ExhOLDBJR9poRCFAC+Qz4LT3nRiJ3VVg5zgm0rf68Dq64t+zdxcz47BcrpqC9tsmmClDDYY4zT6QFiScyOq71eaL4XNQNMPC6vb3XSrN+h0pbh7NjB2LEJbgT7rsf62Gr9zkqHR2AWzJCQ1imq3OJKMp1RVvOmJ65Fn3MnySOoxGXGcC2DY3PHs5fk8jU0PLKQa5Sd7ymDQjnjAhbV/sGDSmfsqv8SobpH+PIq/VCKG+AELS3hFeOckUY1k6qoNm1bs6cP+nBVjxku3hdXPd/b/F+IHElwo3vXb6IIg6eeZaZKv2JNmJxkiYoAivuEWCmCDtyp5RGXbOp6sxlC7hkDApsc5Jd0fKOy3IzFBepjZsr4AeZe/o1bpSTVwQaplF8+FZ7dFG4"
`endif