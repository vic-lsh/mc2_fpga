// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
b2uqJnVLdx8Rlq9pldQuHUD2kM6IDdQkkobZZM38AhKjDTqEubfuU+KCscJ5
hzdh7AtPSPs/zLGK9XXgeP9zWrw9B4CG8Wi+jGtSsLc8GyJOc/pL9cjC6UoD
bA06q4TZ3dcxfmllQ/NYWIc+yaU0S2lqkOpHkDX9X8+K+uvqnWSjAOhTV4jR
W99qCkbKHH5S86rrC8/1vhh/7KuFQo4e8na20snq9fmNvFNhcgOPMY+DKZK9
9CdgbPdGUvK8pAwIS56v0sy4d/xIKDw5nUvbg4FQgy1XKzu1LDbFbLxK6DBH
hxed0GNCrAjppB8vNadAO7VACxZLy4MVma2YLKlazw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OreqWVHSZlP8wsFgbETh+eNJ8PC8Rr7QMU976+dgsAWqUezP3/xtExIxPxwz
V802sxbgraHL6wsM7qu3y7qf4Tzni49wUE11+Lakq06RYWwshQKRTGPzrtHN
/KHfbcCy/3ehM/14PGELzr4o8f7T12QHozX0mULw6OH7Gf6PXcqfjLwiNTNO
W/WI48ypsR9kTRIAtIbfhSRb/elkdK2bRKsmPfmDrSO1kyEnt6WqgB644XEc
yICCZWJoH1spvr+CgwHxH7FxXkmXQa4bnWqAlYgC7G0kr2/HYDDdFPUaOErl
ElifvJJvaOOCLQ2tfb0wmoM8J3ZTQhPF7oYZ4GLB6w==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WRsc44egXWLGbZA+DfzEFtA7QwDXOoenmUVN6FsdXMeE6SPJ56xNjzwi0Zbq
zg1jTVafGpzy7TSIehNRzxAdeUYp+FCJy6ywOdbWYH0UVQpVvTQrA8H2cih+
w6/TOXd1hA2ewZsmG1MRNYN8jD4biJiFET4lQz/24Oer0Feo/ipNnnuryBYK
ZfCbmBlqJwMsYTErTb+QLWvEy0fb8eA/2X7Z7cRciHj1qv59ZIZlCjB0HIPt
Zhjou95pcDTJloepnFFLLKxVoqv7ubxycDwXPUmQVYp5O0irxbKJlNMMMRYU
X3xH0RWtpWRwxyqORyhglwWG6NegnD2pejfhrRDkUQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bdfH+T0X2sEW3msFz5BGFjcm2cQWscTcqeVxDY8HiGonR/0pKAgsPRkbKTBh
MqJsRnEjpYRd2zx6sqdx3FOgs13Kfc4YwDsDFP5mtjpj2sRTHw6MvUeAsNug
AWeL8iWzT3fb8qc1khkWRzBAfB/M+9BNiTWQtBnEqIbfjmYkKGFoFNhCpC7s
zfkZTFjyY6BwpsU06r6oyp1EGpGn4VM9pj00mMCqlif8OnUfXgvo+Vj/FAH/
kd+4sg2Y1olIDCpzm11wHEg9X3YX7JBSoLAyVo/svzwE9O5p+NhT7rLJxB7W
EIfM9QLtMYXObbUa6SCXtEourroFn1hINXlOeYIKWw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
M+D5NGxmmUl1DYIl8Db/IkbI5jH0kJEeMIOuRyF/uOdz5Aws8inJWnoiOVQW
lP0wSr8cC9fiHFcQRKN1hbLHN5NG3tkj+vgZL9wikfy/ZEIiXK7k5Wa7IMHz
L4vZOYUcarCbyQst1bHW8V76sgATlwKEapqpJ/epAJo9UrOBtf0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pRIDHAMJiTgKgOj+FZJzdFdMx9qicm9uGhHmRT5gdodygt7Qgxf+Zukvorpo
h2TAohwBe8xZ5gAVm29Ob3lMYCeYeI817dlE9zCQ5QUoNBSbbNc6s7HLW5Pp
Cv0CAP9RgPhGvwcnFO5TCCUdovBlaiph5LJxdiEMrXjUEYkH5VCl+kD10+kt
wZlCxNBaYDZKr9F7PsuioU/xmUu9a/V54KvkFzWoyk9t6cEaRr38cfxXCqM5
SwXn/RSP9QLM6hgqpV+B/DegV7LOuT09vEAst9dQbvDyhTOJh1SudaVPySg/
GXC+2WkKCUiuvvuASC18BK70KjPwAF8BPrN0Un+/TS4k5eu/HsBoxn6f3k9Z
M4tRxIAbXewQkjtNzExTJVHU0OjiL0ukii5QKTPUXHhjfO/ucefsvfdlVCeL
e3qaihhCYJT22h7B0zA7OpFzEXOKuzsaDXS8nK5nbKpxuWSjvs90riwOCHml
0ndKMH2Y8Cbe6cmQlmOT48DLwDa7S20P


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uyBGK4+iWMB7mkwC0o7kugxC0uEF1wLjJ2pT7DiXHUPM/FU1bhSpX7WzcOUu
3HgSYCLqLMb5vjlP43yPBDuUOkw8bXAz0BbF2p37mKJ2hfLWlee34WzG1msK
fWHh5Exl/Dzvw/us8mNHIuOGjqqmP7shOjrX9OWemSe5Wm+m/+g=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uar91aJAZg62KiNjU4TeOW4cAYLns9O8CqP9Bt8lCxETf+4h+E19KLIpFqyn
NiA4i43JOYmXKrEFZX7CbcZJmSB3mPz1VnZYVA5tQ0DyykurrVSXRDWSiU6O
gejN/x6HlxNOKkHG1VyW2mxigO8hZMix7WV39WUpJvsWqGGyr10=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7152)
`pragma protect data_block
PYnMgF7TfeBWUaxTuEBN7ydSjqQmla52fYKUewoXQjyd+aB7UbYjsuebdaxN
q83QhAfkLSc4edqq7NK4+Zab2yezOQyFJLOaR7WpX9vZuRfzPppit+U/kqXB
nr73d7VaO+ew2UsRk/NIpOz8N9HXi+J55Do3gx25eFt9u5kwafT7gDao7gei
Ew0LmxKs+TiWY30GBgEWZfXqtY1oQpKPTKfWK6D2XUJX7mnS/gmkDf7fEVBg
lMB/xG3LXOJEVCEpa9EYTriR105wQB6OSAt6ZCyvLJI9sEQaSlV0P+TNpeTG
CYiCIsJS4Ur4QAR3MM3hQEkZHwVo34q9gbX5RQ14vSO0G98/YLc4hNRDLqe2
r5pSrwtdcGOi1EM7ezt3lh2YT2FMG397aWv1IyNrn8pOS4hXZVlKM+X6Dhuq
S69uZ+snftETKHgUirDkmDE6/G87zmqVv9SQ9CnuJbkA3CSjXenFiAaw1z4y
7X8AZ9e4iPJPWmJegfWoKLron4felm3CK2i3qiOy/zI9W4JBVlI2B3Z4fnMj
vLP+Pj2fsSm49BNDOhc4oZ7C7KHZ3MbZQOEWrI5lR9WD9QET3bOg8dzEXyDl
09onCHNJDi0f1j7XVKpmrWt6NB6Km1xpCOgwhnyJgC7OGs1ufWt0KvQJnwzs
4NdWpz0pC7EAFSz78taM7OJGaDWWqZRmPXOiDaoi4zIVHqj+s9jWKAkaOARa
VnLJan+pxPDptPSjGXyUgG95Rzk4bQApgz1iT1cG/e5LnFZDpmETylQkhS1N
lxQbGBa8dfsJGprD9+gSPpl+kR7lu3x62Ix7xQt0FToq6Y1BZfStFpc4/Eoi
TabSCrhv9Wy40dP66WYRfwZ0cFhhvmQzdLgbwdU9+/hwwQ/PidsS2k5NgF+O
5VHiJWtE3BJeQBn2hWGRJpuQMaH68H54RS4ok7HB5w11QC9wt+2ye/uezSYM
6+WOV2P18L/xKWuv3SgoJqrbnRuITX4NcZmfRMx8MbxbFq2d7Cs1MazQSP6u
qjxkiOP0F+EMo7bw63b1nTpgr9u/gy0wZyaTHnv4Ys6g/8E2GJ7liDkW1UEj
PPMEPa2GElHg7aTOaJBRjJU3Yp+76ZkwqneKlMn0g+fdGH/oqryRSchcFznk
kaVQOm5e857JMttWF6THCNfyUlKjXprVtc6XIxYMK1MI0ZQAK/rm5iTEsbWD
hPxmswMbeVOfcQgEXz8H6zch0HKYQQa8nxMS+WHWN/WntXb2OgLMM5lL3AdP
PBvYVsKX4uoKLmdGUdllhT4S4WpZafgNaaKFdhYaQmDDAONI1U0Jhy597Qqd
4HTTN/RVyF8XLMN6PNXhsJgivcvA5DJRVDGCvBxroMhPYxEm0TLrsrFvtUDN
C5z/J95FdovKbooRVyO1OkXoH0eDRCKY7v3edPdXDotgf8HpYCYlESvCAqUh
iiJDOq6GjkiaQ4ziv3ZqyuRP9QQPRN1CIUg2H/fqSLY1wWJvi3yEGwSkStKW
EWsq8qlYxRZmiepcxbfA/nlaMiGqKSHPm+XY7e8McULCQnqmMMG09RMQXucM
XesMpjQWpZFPThG4ZFM61tn7OaNC+6UpCKtZrUpRe4xVo4KVQCEpxqiKq7ef
PLjZ2oT0ACM7VrUYYt3nSg+gub9YzsbEH68yetmVCK4cUlZ20UHnpX5tN+kk
mQNhxdV7vf2kV5lMZURCrnFAmmfQjyAfyyHM8HtyktiuYmnRAEoeTUCTvOuJ
ZrHINQgmyolCXKbKM382Ws/GbSEjNv4D9A99CL4GN13OxrXVZ7m9R3FefLhV
EU+0A3Icb6tcH12vKXWdxG+4k8+6n/1gEjsr+BDZs3BAOxOPudRDQk3rgMeb
YjarQC0aRO3Oqn09FO3BcI9YpiGUh+YNTRsUam6dDQPuwpIbLNVigbvYjhUJ
0P0oOF/lojGI4Qgz+5m0N7vUAhIUbTRciV+yx1jYZ0INp2PO4AvmwwMLf4so
buFzHKiVX9cNRO3eTrn4ZlmPdUUV6VzfgVUnM8frNS7JQmFkpNUG/OuL7Goq
Kc++/0BXHPXNK5KGtdf6b/QxHpyUDgrYvmzRydsMOMeA5NLnm2MXQXVHEiJG
yYg4aQo5minQA++C1/TKwiJ5PLofdsEdV/gn54KFdOW9B5Ygci4r0XZnZsfc
oqAxGMOSE2zh2N0qYNKtds+bRy13tA2V3cDbU2zC1mVctCNw9xkKQtfMUzdK
2KMEjIg4vy/M0X2O/nES2lWlluslzinsh8/dcHLzLIxISawXiJ35Oa6NvdkS
GZDAxw8vfOv8s6Dz15OKINhYclVf/apIw9NF0iZh/aAvtyVxwQLszj6uh3VU
bO5l2vdBvGV8Ql0ABNPwIEvHfYunJGCvj82qb/aCbBxMjii8a/3I9NHTtTcJ
JsdwjxHXj05I9+EFVDGmRLXSuVeePerZtWWyvThk3xypjWOp+lAlm4XGOFF3
5PovYWYHWwUjT0R66Ceoh8lw3fAxDhR9zvPUufhi7yda8w5K0IVHLTStINSw
1kVrSIIm9CQTjxXrSkuXP56MJPzJPkUWQvCyfOA7nJUlJR4S4A6GJoL5D3q6
wnPHJtlAH8o93bdiwmoi9oy1CoHCXauS4DxS3s7peDj8dzYCzKhNw6E7FOlg
5y7Saa9XrQxKg7EdwUhwMKi4LWUmF45glcv9NIPD6eG01+H5yaXOHgTIZzwu
ke7/W0OBWdEWAj+QZ0cn1qfHzJNvNEIZbUmlzkCYmg/TzTLJw5G3UC8JUZM3
XEIWPOlSG/Glyqg03/WpG/Hrh3cBcRuaozBaS1+1tIJ9tBQMOk6pYOHJK/I8
QijRUPZmiF7iC/J5+tvpF4AJPPbia5cOCLk6a6sKIsya7dF+Xas9+YEAlg2P
42U+DAe628NEzaPDTJ0JCgtNUyZlU1VCuv9fNAxl0UH362Az9ajTw727P+iT
x8LlPoaWwpDAekGVdZt7JdRe7QzpR0i/ONj7O2tSIAOVBd6uNlbSfy+rsiZ+
5Q/1T3bDpsZR8IK7Z7DAWEmFpES7LbeLwUrMhxsBmDTN8Tklt5XxufvwrK2q
/UGEgRS+yCzSUBZnh+YKMGP8QW277cI6bK+Sj02UT9ft/AQIIboJvLthZWjn
HzJq4ZNhesAIW5chb7HWXZKXgE7QT73tdB1h0Q3t8EuCsZKg2qVIjr3NGJqi
4rBPPg+RmaWkNlqQcdlL3M8SA7he735S55o09Px+U1WXsKIGsWy3fZZfRQVB
NmBVzQ8FNk8kmFsCbuJ3Uo0J5uSnNdPrZrNei9drcm5kW1NsQQPW8Bv5cAfI
DzN3zBZ4V5qvwxiHyNWVb6O+meNy1+l8zPRtveDz8To7KU5c/mp5/oddIcbe
Qri0jIjPd0h2xS1S7ILvHnZaLIPyRb7okgTdPgEWbCpFAyWfvhthcEwDLgF/
yCYlsXDg83t0rQjzxRwzZOli3ARKm+Kb+gIQLU6VWEPRR89hpOb4Xg3T1iY8
h1Q8891ZUWLUOxu6osQE6q9+v518vJQkA9rrJOZvGrAN7iUfrN4ZNSn3r3TT
qu2sZia/ISgTJZwlg3McLTd7kLxy+1qGOevbeBTbiutjLxDTspHCx90foSlY
Mxcb/3ozb8EWt/0Tj8mBTLMKU+Pi2zBJVUHIeoVQeq/DCZypjNPPS8WTzj4i
6ANGsbRa7orr+8+6XGzl2EspVYneGgVGw0RhWCnF0Ksg5X6Sh7U+hMuWMiQK
5h7ZT/60nNhkuqvH5LVn+AeDgmJfik9BV0w9wqwskwuqaB2gZ1gefBNalpKA
hMFAVYcE1x212fx/e6QffuvSqg/fr6S0Rr4YuvKrj0VPJuEz82oY009xXUvW
umLoXU4N6WzRJ8fuT6kWRFFnFykHSTounQG6iKlxP/c+dYHY2gSGmy3fog5X
0uMoGEwtxbRuOz8sQGsiSvSKQU105z8fSv4ft4iAQY7sHMhNkdtVTIj2ML2R
Mgy64mQ/a9ZZA7aTUeD996LSHrdS2djjjiMU1T/Vss3fEeazTVJ5rg0wjPJz
HunB1rcC75TJqB7z7N2okijtJlya8L+sLxx0oboHFbU/tJRn7N5nBPF0b08E
RmEMZbwwXr/Am1PXW4BlCf6L/Lzv/BIgtk6TNJj/PtyKQlXBWmK/xpEM/PMR
M8zR1+5dn9IyRDtZqW10EjLfi5zViD/Jc48bRsEGPEYbnd0hhebdhdtxQyEA
INLoh0yYor46aBGmVibIokqlsoXs3VvcKdd28v/RDti+StRVAOOwEQCfZufv
47gGE/mwJIkK2bJy8oVFUJ/t3WXIqTagm8ChItenUYkqdrd14KT8TPnj/a7l
IWgbwE02AwzO3SYBNKGgzvPpWDUEtQfQXhLT25mRFUdgrOJ+EIzfkpb14rVb
evL0e7kOANq/TrtRkw5vFL3FJeyIus6uVUsDj6rOgk/M+EBMdVO4RoSjGcKF
2unV47TM9/sVbYXIqLdLMKurZ8Wi6YFxSboBrEzocsmmTBaMS3ihERNa6Kri
j02nHD0auNNRhiXNwageW2JRWBBV8Zmi9agFVDtu3UHO38cB0sjBN29LME6T
awZvdol1zgBjAxJb9pVap1n05ffDE1Uxxt6FHwz11htyQWlrJ/jDuJg1fUCv
ot8BeTHAJF/YpBWBBPxptz+kqbPSeNd1NDC8whgA/u7suP3ul0Fcv0xZbsUA
7fDvdl3mt4ZgcBxkacPj4YecpLekqvVUkneiXTffEKVWFkvON10RTZKIfVPr
fKSpTMaF/S4oc+hkLeRE56bnZNt0bAbcbfgPIqZtv+Mm2lvd3vvO+5gNF1f/
EeFPEUNs9XlGyU9X8vFUSHIb1wQQR2n9rwesFkzrBVh+7dHGxrEzSADh6Osi
G5D6jtv5w4/HFWkV/ctF5p0tP+sY052l4MN4kawoB1if9sD3cE4+UjiBRiiU
pL5LsFqhvtF9JrNNZMiLB3NcRnXGpc+kZg5g7V+i7HfLYSNp7nqB61X4RI2J
gcQvj9k/d6FA33tcnYydZY/SpkA51CiXZu5MuSdqTi2ug26EFB8RA1CdVI+Y
gw2ewdMColxGQGEbQpmKgo72U9PNQMW8eWgIaUajUiLFGkgB5UTopaZmtnlM
y6kqcQL+75rOS4wNUi1j2gIDHSmhCktxWcW1gr14XSQ+VKLSb7Z/OTORiAOM
BmjI+0JzoNRCuHRnQEJlGYbyqwazm67S8lwjJa6Je7rVb0nLguBTzKsloJKC
aYDvZxH3zdHu499BDJPPhjtpzWcl6A9hTQxEnxU1r3dzMOi2EFAGkboujcDW
oRU92W9w/marPkNTcJDFP3KpMqHWhyeRiPM95PVsfbptYv19jmPOUhXK3QvL
8drmVinpm8Ccoh7OHIGDRlzCjbtTZl8Fno7KQZ6MtKxjdKNbpL8cOe3u8baQ
jDBua+MjieB0Gy+Z9dAS/Hq7EWsxv87m09SSz9Dr5pDabMh1gpuv3WKlBjkd
apLM3b8MYQx4HktNc98rprXzpwOAE2AVIVAKkURPQGhlg3mI9gfTmf2+ox3S
6xecu3l1guF/X+3DnAc1b/twLoxG2uTvuEtXXx1oKcwpcFL0iuYTIPEQ47UZ
AyHoi/UTb02XeXHtjBEdDmZ9rgUkTJNDpbJFxwThtdiSCRpcLI23/1NA55OJ
YAAgxfLWug2vZsX5on/j6FATDAmDHzewJwVKSIgOhu6+VIYXYzvsWSSpVoGW
C+YbECa3XGoIJ9K20rYevRaMYkUT/yuAJ9S1oSHB/anJUssREf2FCRyI9y8o
8h9vzduieifQ07WCo0baHN0goQ8lRU+4ZuROcHgg4zQ95ZggXxQJxWlrhCyj
zyyoOLQY7TUWDd5Fhosd+OzzBQerMzOPZ4ZGBbl0kOquFjWN4dbwEEyfzGs1
VrFKSjPwguPpvlf4l3+SZeBsi3XbCwaiiYFB8mgmAtt+4UySmUZTEzdWentJ
6vYEtdd3AhYHWqd08dYz+Q0e9BtiyYMwTx1fwYnFSkQrDcigz0FyiOQCQrTB
hl9TtE0rVidH9py+tm4TdkJmaYKFl6j3JQmZzVdXHasPUNPGhNWVZAlRWaEl
4/8Hkp0Xaab7PgRUIoB1rsTVNaTtAG0OloUojhRgmY0n94N03NPT+delH3Gg
Oaie5AKYvuYZfqhsujXPVc0nAeDz9NLXXT/A5EXcoSzNGD4Z8lG8OnTvajWN
706Nld/UEl91k3cUUG1y2x3UOir+nY08uquKq+29lNYoOMlvcu5/T7FVIgDJ
LOn/mIGZa575qBgqE5OXGsismmX7bzuR4Uo8Uc5FD3IqzFygiPJWLlIWVCIi
4UNabk7PGbWWqWmAA3DM+KVl6YoFYIGKSiu8YfN4KPTTzlNRVCK7YjXIQDlJ
2aXj2V3cxhAlEDj7I7JSb2SMqmNy7pG7SCd82cX02yW/ovxYQ4JoeULha701
3R/1BOhdo4VrMRb68EC5eLpKC+ZUGkM739nBNumK+HoThudf2wvfoL3p5vRA
XwuU+ebJPu4qcDncEhG/CLdUIiy9RvdCA/QDVu7FFICfuzlqERWkzCS8YaEt
/046wbYFqM2isyUwMIR3oC2yLseG3qo5zN4UX6o3mIc43qkAciR9s7ffcQ3Y
kkVJe9+Wnu/Ob7aABGTOD8MyolRzVyGq3ql1r4Y9cU1SBjGDUTbSluhdLHyI
NUCYyXoxbjcMr+ktDVKXK/iUAG5Dk67HUTi5Nog+1F5v8sY0xXF/SbPyXJmy
VCboHhlaWJHHyfg6MBik1nkou4EscszZ1ike63ttyfDxbfiNKSZmL4ZgQoRL
OUKsWhuq/W0gC/6E17S/7Xg8Qcyom3jdCZX7Id64dVa2gL76ysaHo3YA0Eb+
2JmIVC5VscRMbEiH5yMLplkYwDc1qHheIPg9iju7I1u4JHLXK1uQcCxVjPGG
eUxdjh61VoQaxNSPdPB8mEFw5Vs8vyKlvJnB3QDaMLga5zZi9nhoxdKWzjtc
0Gf+JpNyYtHXbgz1ajCgWjYlPoMaLH0astKjVyXYxnxSkc1NguOOYo8tMCJ3
xByj+Ut1Lc4YHqrb7QPAXmdWgbGSHlvrsOQzbrt4CYrRuJcgi8APXqJM7dmQ
SRdv8sofN5+/tUyc95H+RU2Ae56m/ckpOKfWf23fH0fZhOSrvOMOGS43aHlN
cwf1YT8Wlpy6xeEG2nnfbtvz2OHYES3c+28G/W5UTqitLXeZnU2ikRd+Z715
rsY5QFkx+cSgL07L856v5nbea8g2FvFzPcZM28I+FYvu/OJFYKmF5z3PDb1f
RlS0KnQn4FXxIJwGB2DfRZjxwUBRoIrZy/G1K8n9dmFaDdHYnqrmpxemfNhf
X8mFePweJesKU0TndhAFav17a8OoUSHqaxLoS1WNYzAfxFk1GxLfq8lg9Qsh
F7G5ERLgcgtxAMJjM8DLACU47B85PVQ2jRNe/G06gZoUPGMvU3TTV2RqzIkh
hzNE2YkDz5oUUyw0GFIKQq+bH+beMsQGWnY+DVMkRslM+F20yyl2OXGv267K
2w96+s6LOHH5Q/jtLNiUNkWJoFY0B5cBrRa+q7qizlZus1UAkGgWKVGcsSbB
T4x2xDLUp3KxABuTeImaxRBA4xirVl9eQU4DkCTnH03IB6tYgexRLmGVzXG5
9eR9i5xOUW+szGuCbOQIj9dh6x9Ixh3NrdXS3mn5mL/KG2DB1i660NLJQ4z8
QhwePhrma/+htfXDwzDwmHbTEWJTEdjK+9llpltzI9kOvHZ2WeuGtSxk6Q+a
mwFM/cP8QnBS9utTKh6XWuqeR+wHVGhx1cseJsGl0DM/0bNZp1wZzEcPz/RD
ljUEhFtKURMa9pWNik5AMEuDonSrjuCtVdJmFkyQEMFq8G2SjezMYaAgcWNz
m+crO6lJeRYtjQCskL2bV/Wwo1f3KRmKqPMnYiTmDOtLLpyjEg9VrBfsDEV0
duMlUf6TVyhxLTevCNQiRYlRGgqVq8Aa5bQ9ePFCIxUAJpZMd0IgQYAGtZet
UPqT//3dUJv3h50yiOo8YSS9pA7n4SK/kTm9ARFhpmWMkfGXZKjcMC4LXeF+
PyUnfgFjDqxEWlUzFDOA0njgBqZr0SRLy6yTdIBYVsbqIwon4doDnQXw2oTQ
Ic34YpQjzScwcPKZ9Hxt2GIe2/+dPPmaCDadIk+y0DFZFWdv9g8ifwKEMjp2
xEa885X4TZmde/gH7tomzoN9L7omHtAWWSm2OTMtUcJqfxKajwtWwgxmRE8P
+GBEYTBRG85ZEe93bnDMOSvuzumDaiIawobYqbb4Ea4t5OQjztNzsO/R4fcz
5/d8mmc5xhYt+8LSkE/XmFagIkV+foZNUY+5DqAAeOcs/efUvlBI4sOCP46i
n4jSMs580x4zloV8gkIJpqyPuZHGnmFpHgfqOhhoSQrznYQ0LLz1enyXFHxT
mHS8+VBODgYd66yWWUTnzT3d5dY2i9Qjeq0UuRK/OKEiRngOEURSM49of8md
sEBiQQl/w3J01WVombR0OTnPaV7CZT0Mm77qNL020XcxBJobXcp2pKDSJ2k+
IS5swpV2D1uSN9Y3RQlHV+V2yQgscomXlCePgAoH3zB9ZDlFeXWpxAtm3h/S
czu6EaevoletYIUomAUyFQxnWhUp8ni9+XbgxvCpRUinW2i5UMM5dsARAJD2
VHgKWg8XQ6HfsGcw12dUuHPaXXQ+Oj7rIl7QLEBZmQzlDs3qQO+8SP68emWu
1D1rzguxRRu4yxXpJW4JfVSoPI3ekVvsmrwpDywrAlas1QHeXtG6CH+pEXZu
BTqo7KlNM+pnJKdHUAO9G1TtK9GvBQhFwN/JDBllhl541yhBzRhn1QDvnwYV
Zz3YwfqXNCRn1x+1o4biD76oSWh68UENKej53CgcsvA1eTUMxtBx6lLjeTvh
sYqJAdh40ivIkEMphGCBAmfW2Qdpwv20S3xIeyklxTA6S75N1Kjo+cFdiV9d
xEKL7REjbLOcmmzTENZkeIt7ywjUxNm+DNqcEH7Ryvm0NkTSYhr5+ZtXosv7
6MGz8omAJwIdtM09idyGbdGsGtd4bxTncxwQX66uIKJmC/QmGaQfvjdc5tvK
hObuWO+BDjT5HNaztfxRq6D0NZ4977ry8pt+EUjFV9QVICPQ5oeQSOLg8Nfm
izr5Z6lgxk33SY1a2dMod/qAu00v6F0uuDkYILL4GW6tBH8Kk4GuIuZ065eR
BiTmssFz6rSyMNllbEa2EIvHFr9u4flGTN/H1GCE5wekwZ9KDcvQC4JQ9e8a
ckJG9+dcXP0eOoOBEYrX1Esvg9dAODXRNffv2iLO3dtrm8eixY4+pYC+RJUy
8UzfmyH/Um+QizkYMn5QanKK8msg+rmohBiExdlSwCFx6ZO+Ehrzs7OUFRlh
06EMJsZWUn0WFUtZ0BVGOuvfetkFH5zrKC/jt+TVqR4LF8Pjo0RwSPkosFAe
kcX6bCPuf/XI9YG5zlwNL20T3kiIkw+NXROkBbvZ3U24s5P4pWoQ4WxZGksU
2LV3GPCiUjv6CSYIP9Zz26TUgq0cziB6EbENJoapCoh5gliE8dE/o4sg

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "lK4MM9NDeLrdcSiRM+VIuNgpOLUAzWAt6nzBJ3Vw5tvBogzjtStM5gMJjD6PMmMyupOFzYouKIpJuOZh/11WnQBMmqEc6gvbtnHqfGmxFaxYyOv1rddc1B279ac1WEgUgi2BHG6DRj+tHk4+Vv2VvppW/Z9gUZ9e40aCxOYZZHwEVb/SJ8ximgD4Fihl81LOgt6U1JRoR0S/yAHMZXIkaoJ6FVEBkPAD3J3ew7MX9ExNjVmwTMMxYNl5WRStoF4+96XeLYGpKmZLasG4t/G725jnYmmTgvdfsjWpsG2dwNFjJnbqe/N3T1Sa/dtUEhlL80hNqbT8c90hfDqG9u2hT1Zpr7ggVUoix+ho4V5T9sPGjvsUFD85cRuxLGiFjmVmAGfGp5KSAW/Iph1BHlyw008OzD2zPv5IYqyKYoQCkkunGmBiZCmdc5KALTSWwnLm3vL1nTQnlXNKxCVcNgWQ0NabHyBW17c1gxyGVT1BWFZtbgEyZ7th5B6CvLryWSJdUzEBDnP6RDn1RyQ1RCv/t2FpkfQ1ixjjChk2YHa3qzr1FMvws+2fiYIGj9TYTZOwRmSVnDhsQxLbooaLT0shjr2/9c85tHSj3QehcauIZLz877eAqauB+oldnBtxrq94CqAsv761m/dkTVrH1+IdgE+C9xY+98T6tJDg5RSX3+H8KauTeh9pNJFGQRauux+NEOvtRchL0GBVRshzzxDWUHcXP5/KdR1utnaDr4Y9h8YX/42eHXyAOlOELWMnBxShYesufPpd1fC20zROMmviGNKJ/l0SpEiIg6al087UwyLAB7PqJ/LQjYtqZNOxOYvfgp/Z6XO+B3MMuSVRXljO0qh37eqiOPLqOoNJttgJ3o6OpCGx2Ty0RvDpRHQjT9Ce7J56PSJtQ0Calg72Llzl3sQvt1vhyMhiughYJ8BYpx/wteOmfN94Sa08JS8HalQK58Vzu3YIHD0tY9yahwzPTrRr32X753wDRTYK0Y1lcAvI+U/dpYK+ChDZ7Edd/Yvv"
`endif