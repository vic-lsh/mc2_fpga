// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
h7iUPEXHtrIPlS7ipIKp1Ly8q+lkA8Nt2kXzdxmk0i5BBbsSkYYiBP+1Ukbv
lVResDmu/EO+dSuZ+UGCGYITcfoMV6ZREeJY6Jo8W0CbMJQRat8ATSPbUVkw
Gqfy4w37NWPUMh/MyKdrwA6PlMLI6+fSJC4iePb9r4yS4nomdrmSsQ8UlK0m
mFisDMvFZC0dNJV7SeNe2eHxnHMo1tqDVaugL0SvXXQJe27qNoTtx4oViaHJ
cKvypejhv9c1CMHJjeQautAzsMZ/bcCnOOHGoKKQMLyKJVfwmK5WsYYf64fw
z1wJe2Mnl0Aqm7IdbhwPT0mso9MvTdwy1UVldlgoxA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
l3KVnXiHSax6QJJXjigXpLlOOYHLPUg6jr9fpqN1JXqz1ksx7C694lgDOp2/
nlHV1Aikqu5lAhwUgMI3RmuMgWgudLofc32Utc1pFl+CoOiG5OkrL/wKkPlo
+nKohmH4bBNIj4uGny3y5CNXpeer6ozeNi6+6vNyGW6XfvLzOopBA//TIcyK
jIR8Uw9IKRmOCpsLvQ1k1YjW4p+cv2ksfb/xE6An3B/PPjxzAx7cWq/6V7Gc
5U3vz9iQbfjne2hLAbYffvpZl6ISR4TtUwFrywKu7XA07yy+VSWcHPpeTtJs
4ZoOhDjk5BVr/pDrnDcvu+QNxWXA25IHl9ZlBUt6Bw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
uojPyBbl+HsI98j0cLaxQSRjkao66QYHVmdA3gwncimy0MhvxzpOm02klqJg
52dibvugFrSRkrHmIsq0Ga5SxqDmaEY0ew018jt/H6vxgAt15Mw3dYXhK93g
m7XycitiV8I2xi3d2eTEwd9KB/OARxfut/OsxuVtENWaO2l5P5RMkFrbDe4p
1BhIAmT//7IJBzvP/QfQi7PaJ0nnIbfSZ+hwWwX3+bMQsuoscK3Q88fIUD4C
hDPfitPqiIRRuWJMJa4L9dS0ixFNLAV3RwtkFusnga+ygLZ7RRQ9lwjQEFBn
9qMyayBz4J5YWUzUjNMWFFTZejC2LazyNYXJ7ERfiw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ricgjoksVxHfs1g1OCfsG+V1JlwT2nrInHAo6zA8OgDFzQJWyIG6IdOJl61f
d0rxl22VIkejJl5J41j+4fQLQMCcSyTtlhattlxVrDMgtlfRn+kqrvC0Om2D
en7nFGT8p9YAhTtynQr96vVQuK2O8HYnm3SqFBb7PQhMvCHdlmaXHueFf3XY
HhLzWFiY/b+ZEYO8d0bDCZahATal//Sdg4s4O4ESQIcQMYuLKjLrBxeGgYR8
U+HCn4hEOps6fRgFi0tMfey6il6f4Dp2e1RkKNkb8NXTF9OlAJwuOyLzdKYg
786a3AjZhnNsl83YsCRoLgFq1ODSdOxd+PdQosw1eA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HOvDKi5XD0OZQI51GMq1+uHBG8UXg2juUN62hWI+DfeFPUHlB/7x+Q7VJNGm
0x56apg4tH9V/R8xBK+KICtU3l1V6rRXLihcaaF0lEXKZgLlx3rnUlVrnmVn
W0xsdTyhL7lGaewueBL2OGq75lMjqbaspSBtmwUPCtZOkneIZTk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
KLogeZ0X+7zMa8pdnlPUmeR/aSMsIRY9bT40zc9M5BZu7AhXeMzMPDImqwQx
dQB9UqHz4nWMPADTIQ3dkwwxgbzQMcDtWuCkHN/FKcQ+++2JEQNfT9i6wAop
uzrD8ZXNr9pHc8P+HBqfLyvqCH1T1a1YDUt3pv6BI0L81nYnZHTeWeKUiHpQ
R8L3bAPNmAu5Cf6sEA6kdI2urUfQ6tTu8OohQ71s879B8JSggjpoU70qd3AM
kTrvNZn0brtB1i3xZpfVRHsvAd9vnD2ASZr2W1eYhzhotcoxO6NgqB1dfLFu
dlr3P1Taqmxo0BcQ46BuSpGHg9dLnLH3JgBU+HWEv4krALgq5A+tH4duT6+A
grA3Ym40LKx/8qxAFoTiTREhgpO8JAmURxU76U3Q+alIacqPVXFvSCJQe6mv
hG23IS7nnXWqJtvuWj5X+x+d3Lls/U+yMAsP3HecPVKW7pPGo5hTjpLI6yRJ
lmEo0J5dFy9YZ8pZ3h21oDvbBYSU0JwX


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ac+o+k42tCBpKKa8W58o5uK6ayUW4nuPxPIeat02VGuKusj5nM61Lw0RELSi
0saVs+4zv2R2IxxaSsgoHOTs7ULTp1hZXF76A3GQfTfWWIrx52XXyxp+2mRA
P2D2YDEgLLWD4dO+UxBUJ+UMo644GkhO1XcJC23KNTwfB3GXmQ8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lLSHZN2p3+13HXCS2GXoRF/C9Joujemdtove4J9F1MDPj56IOhnUATCqgtwz
JZxm2UpehCGXGVyMrR/CkdAkxa9ZXLbNJBzjJU+eo5S4OTKECBhI0m0G4IBF
PBYhrhjFyobERXqr25xNz1m7aPVUY7/KNPr6U0HjaeCGKFIoamM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7072)
`pragma protect data_block
yMggXB3qNZTKkvR1Pr1ZV2uuYJJp1evio+KYqPcZDthAvUlbGZYr/7JNRQew
nCjDEdSxF3lMysdNJbwbOxtJKK/XHCajgVsYvyqlxWVUslY45vM9Y/jhoMat
pZRIzJJ1WlYXwZ7s9dWolJAVSbQCue7P1kHOdTu0+H4jjLV3EwLFQncp8Amd
o6nvPV0H4y6Gr6uKvuu7CE5jlj61RCB1zuV8LHwt3EeIhPjRlUEPMZ6BxXWk
uPOJNEM/LvwFPshIRvEfc/c8NZVE+VqZxkzPxuiinVos2Nc8u5BVnd8WiqEL
B6uDe4H0CRafoI9sKWewo3XHNuxLNh7szPIpaBcCDFonXtAj6lU+Z1vpHN2h
hA2DdGk5ZCz9HbmLKxN3H/Ye+iJ7y1/IDOmkvNirhsxDKXrH+P43JaAisHC/
vtgFnedW1krAooqgKa5izilAN5LYCKkmihbNrwYknGs63iq8Pr+MkjtHOj2+
nkLa6r/KOfdUppnmUKuyOfj6OpBiCOAJFtXKIIn2TrSRqjBh+0CPM5obr+WK
1/NmLJxxIB+j5sJ54vNdkJBaIBJs8rdNFkU5HvlbcKrNDVQXSMXksKwITvnT
Cbv88Zur4gKUiQKOU18d34AfBtaE/a7ms4f3NlgKU6+QIHSLlSrhKe4XMxnb
l5SIeL72S+Ii7l1WGaWwsEEtm5KhZ8MUCwJ6XFjynB+dt9yrDB+HOE6CUrzC
60MAN8eLTe5XLNrRkptm4kIEIkkVdjEyjdvgN1PbYHvjxQc6DI+LtYjgGiSi
mWchNcCDf65GPLIfrJvhYQf6IwIbu7M53Y2PqeS4yq/pcYAZW+6/dF2ZdEGw
1K5pSea09Dd5los3sWQrcpVyqH5YKm2V1tEXvCi9isOPlnB4OoFj8Gx4tsxF
PGwd5Be7xP1lGnAhuGzpRB2OErMeF+E402ngvrIygUF+6966irsW1KO6Aov/
wxR9fA7OR0yCqcBW4cn4JVGfZlsYs5ELpdK/hHT9glHSiKPBI20lpuLzeAQY
TgwZ4V8X5Hkocp7nVwY5332u2l4Koe7wv5Cupxo7jJhTb9xsEkHobsnfTiL/
PeSR30IQ6ehAtZuyrthcvhvGjf5DCjHsYMjXfOBeV0gPjRU4XGjwQXOK8hJC
9vkyzJSW8qizDFkB7xFD+9852TiH6hkqki5ivrK5xD+jRD1X4XnysPz+cRoa
Ja+IgXnwnW0Ek+l7AoiT5gjPSnHdqQ7kYjLDepJhtmezZSxSta/bRrEhOpeC
jalRmwgQ1gjbJkrQi3pkv2E026TX846iVFJ3Gg8rbUwLsl3NwoS8081HSKuQ
6Yp7N1KntBFr7PKIgP9a2Xi+W7rJ+FsXeZ5GXjI94HZCkSgV5ScbJe2XmU7v
tSolql6b4QXBocecoUmPqgXISc1Yr71VwLpkBMrSa2MOhMqBzR8uUZtZYnZ+
wqIQzw1Wl9vZKruJO1Trset10Byt7fuTuVcZUBZgmMI7My4fBfSqSI7Ww2n+
T8gbz6Y8I7TLGFd5tgniDs3u6zbK+YgzNLcFnY/jCNTmNtn2/l0OYk0YdyPK
lnbECXbg3G7eeGFO+yqZ3G863EvK/n0w0KDuiLVIs5raW4oxVotjAweSIawQ
qQwjYpD49XymrmZXtO6h9bNvh6NXlLGHJ7aEH5nKAiKZ2J5fG5DVteM3t+sS
I4aNY1y6fDLiV11/OyhjabBV5XTphVlZyhZKshyCE1k12XgR+nHlzp8pYebP
U1vFhIa+jQVUqiC0Ju/8A4DO5N647SIhR71vXYNbAfWcIFgzJEe+91N9FgXU
sOKSqRBA0GKd6Xws4QAiTFHzAgMSmt/1fhRNycCg5lw1xn+Dd2kb2bwrUdhA
ZiTh78WEzoYEXCUM9LG6ckNIAFc4ZOvI5VGHwK7RdMhbj3qOgWpUIWhE0GoD
39MfdWnl4ib4dXAr3hCE7Tt4eOkOnLJaR5m6+oYZet0gn1xgKagMJkus4OMq
7JqeS2yEVkHcPN4gaqPooYRTqDnWJWdq1gXGrON6N+fa9lmjmY/OOOFP4P/s
K8r6BGU2nGm5zh+UU6KwzBs7V+l4SV9Yip4xrA7wd+i4CtnC8Bazj3i+JbQ0
jHBKbkAMdkn+L3hx1yQOkYkbCCx1/z/nRSWlSrXrf1D5qC6r/TEItE0lUNnN
zj+sK3nW3QSUjGMInfnXeynEZ48/H3xBJEBnzCM94tsnLxIHxqH06sYQItPD
vjmIlqUwTASSHVQZhVtGI7Nld2xYQiQTxWnFDOJfV7+OmhKKG4ARgG1eecXe
7OH3yqh4CNc/l9PCu3IvQWVroT+FmAGvNKKh16qJpazYJU4ECx6HUGK+vmmo
AwYpMOBbs+RH4/7pq9PdUMgJFmt6N8Whpw+P6GirahEgEbC0lCxjTxr5W6BW
g2+JjZ8wBQ1MYBIG+JEq7MyC6D8i3yufq4yIrIlJNEF7dsUImopHXrbSnu0m
2jZxW6Pud2xE7mXxyKwOBe/2TuqCS4QLopJXPcr/rX+ig73C3XmtTu13eFey
6e4YEEMTaMZ2IShvd0ZXZMVdIK7EvsWxsug11dM6sWxR5oyvOJ4xUaVailSP
bL88l3lXi4wssgyiIThGGZGU5KfYGv6Tr4p08i4L4IDZnYbrThrydGp7pW8t
fR3VmGP1/V3PKYu4wi8aGIFBgw9ElAeu4L86HLvU5to4gzyl25cCuQjr+E87
ur0prvvTHyl1W1q59kccO9kXe/vKJKeMv2P412LueIupEk30LMxmbRw8C86T
7nTRhdm4bCcXAbSAUJyXhA0q36Kt6AyTJ/ZtUmF86B0Qz5/UImbBxxLOZFdB
1VZBEG2LBXjpR1iOjyT7XWRUo+Ihq/MJMHjZY7IdxGIxo7zkIIsVDrlFn+Mb
V6MpQlpMhVmNQFZi+sKTQNeSjZ6EY0kNAIcSmBg1WrXZR4cp7ePGZt4pnAcZ
Dtfw4cqrFVXCe2r5ZEGf8DWtohBUeMxbwu0A8zWauDOroV9fVGTM742IX6AP
iuVTjLOP5LzGSj9y7zYV0WVV1xdk9/veQIIveeASsO8wcEDZHNw5RTENaFnW
p90K89w1n80kHsZfN+w1IzMASjUUlBr9bBGhFmiiCReXH0EjjbCXE4shfytT
v8eNypg95JKJDxugS3JGpx6tgdZQrwodiVRvGF5iNVJ5MIiiGLs14X2dYjjf
x5bYvmSEGoXydpHi+jUeVHIUA0AkP97eeHB4V5wMllI4zW3PViBFxFVDFKyx
45bmC7G1iAibkVICoubSwQBuA/1Whr0ys8VMhPs/JuZ/fw52M4oCklkCnJFx
wIU/k+RH0QVpE0jzP4EMCSx3W7AGsTAAAd/A2Kry8KoEO0AxAl11q3YX+Z9Y
i7ZkArbAo48/ZQMH1DrQzCag1vR2Vjye6GIYABE2HSwEoB//QzWdt8zdvEQF
PoU3xVk9hwLjF2z9aP2jsJccADV/sbrrCLvFb1QUQJB/j3Odwz/6Gu2rAe4p
RvgvnawJvEneLSMsRaAWb6rjEFkStJKouf4gMnxxYrPPK52AXARIz8G2O84l
fjwXPtzK4PsGBO1Py31TXPIegHHmWeZMlvZCLQQkgNpTNh9/2VUBxW0OyRgR
n/sjHMjS+KIYAq8CijNaKg2kOtjwyYuG3O3pTHIIf9LgH/KPfCuUxiC8CVv1
EmYeRKzpVAmx7Yad+ZIsjQSuztByNT4xcJJFL384nN4pO/upzRgJSqcjBC7t
I1AUC72ODbfslrI7W+hTWs/PaSfliArFT1SR00Re4qdomhwh9e4HViZqzKe6
/zFD5zC60l2hinKAyrexU1hKzRMDYHuGE5pdmuaa2423c1YnIPutRHWHfRKG
PD9zUSh8f/EkCPJn7/Vy8R/rpMQl8xzkbJWMYaptELSdmSswrZNUn9RIeu0+
cbDHmwqA8vJpJtrt4/oidRcw0p88I8K6Crcw/u9lDE6z4njY8WmuTIuo2Z8X
eSXjja+QQG77JJz31ltGbKydp+04NxlxnAw8kqzN/62q2GKjDn3daOIbZKeB
06NPveOgP3i0msBFMjflXC8ikP5L4KtnG1lEoDmI5tnbm/dBdWR6G1ba7gn9
7uCA5KXKsQjGMUfi1raAwmzol0QiQ1451qekeCOZjqOQJbebRjW1YZREVhvP
xgRRjmR8O0/87GI3mFM01wYsk6G5OllPVEh857YUpsurmK4chJEnbndRLnO+
nR0DtClFpBuSWs9bVylP8954dS2pYy61be8EGgBk6Z0w9yiRX1+8zZ/SRfXS
b1oC8MXRl2edSpBCh9aBITvZvPe9RrTsK+WMxz4hg448g7hrCp5brfFbx1LZ
uLEcc2UNVSasxfpAyi+ZWpoW5MfpGts0kSoDx4tzO/iukQhuwqXIxs+gDbGh
FxpfwYcCIZklH/ECeRHSbXaZYz3CkuKubuyc7MFJnGZg4k/6+zUE+aLtOoo4
3+Z8hFQ1q/AwAmhiw0vde9R3F8pQOTeo7xJqNg4THAwTL5M9QJsa/zUxNoJd
67gqBEWlpksqIfDyY+m4ckA9MXhFV23Ir4x1s2lhI88fiVjobXX3OhiBYxp3
bNodyLCunUe1eRa9kPLSD8FMXBzBbACGoQdpJAWyZhOiXbA1R9PZq22OYBlL
T0Kc8PukxkvBOTqrxGKo4eY2dUUODu+TAkvldTb/9n/S3Y8uRSAQ/x3P5eIO
RVHzg/W388vBIHuMw7wRi3PsoJ4zauIX4JU9B5Qv6Dx279DOzxXis3sBWgOe
J0rYyYP+jzfZbNM6x+xrxckVbVKPXoV0HkCOrOAIQ8zgm+6Si8vJqeY+FOmq
tSIDHIDHcAL+SacSgqV8c66M0uCuIFhb8mWNERQSEsxqyihez/kiAPM1aWgu
TaM1IiUPKBgEOLnhW+vxiByHsn/BM4Gt2kjdNpZxs+NIhbnr/Qdw4Rh/NmkI
ns/CRjQ8H9Hics2y/NevW+rABdb1T41nBbg4tvnqMogK/mXszlm4+vaZeW/I
8URkGblfA4/01j1Qme769JJ9uw85Lz9IqD1ZxHdFT/S2ZN8fWXBIl5LY1gb6
prpiAQfbO/1/IU0aiIQ5WDdNsXPkribLrM/igYs+vgYnRA4EuUuheIIIRoE9
un/UQFT8Cvl4JOUL9N3fEwUbFuERZTECtFPTal1d+goyeUNs+4bGPnI3tm+D
9c4evKRQchLh1tZnoddzhJeb7N0/MFMUt0x2qcBc4z8Zdpk0LWqz1uQtwPy+
/JtON5RlcqQcqjbuK4pJROZ8xTBuu3MzM9YpLyz8FTp54ouxKfDzkLNdAcj0
dHVzIGoRvfIkdWGjCt64hFA+Qh7hqafwYdE0sIIHpy/kAQKF0HN9WKviLLgh
e3TEgVu8YWPx9vv3eqxwbNftLhLuK/59F0jjNSOkB2uCR+Sjcheu3tLWmb8l
WrLPCMIfLKu5WvvInEHH7mGuMv0wia8iJeowJIT67bfJZV9o2fMb9wTbPe1R
Bc+PRDN6vKMqCQgDFIqwjk5Sst5/OFgu0uDZ+0FLTy0Gpkp4F7gXE2ms2mya
b1iCoKR43gDzUDYB2In/ZnOWu8G9KXkvMzUtp2EygZDp3XQ5MA6gu2KPXShU
Cew78gde+ou35WUWmzbkIn/WkLeJQj3A+dlTGkLdb+03EBTt6HgDT6JR9ef5
/062BUFdx9BGLE1R88DvOVJfd2kvn3sGdsivhe3OFKdHy1pHjSWyi0Lyms10
/D901Ydt9Nghgn/A/o01HkpPVMrXybg+h/9ucPDvaPYX7M75lzOeM+5/Xdek
kqRPtkG0y2bdWWSPo4pi+S9fu5/+oVP+6OZd/RHYPHOwhahre30SiWkpZSAy
KrFxpue4THfQ/aiV/oqStEnU1Tlb7k6b6Adc/jj1X6JZbBtdPeXNf/kd7T9U
A/GF7I1t5pnAASSMH0bq7n9pPhJm+v5gZn2KVhoRROnivWbKyO5/Bcmadsje
vXgzFkCtDehgGfacsNTcEGc6t2Xo5aEpgDXTF0/Ke8OW88jNEF4iUD97t02I
wlOf8Xg6y49Rki0Tul6HOl2Ugc1e3jw18D1TKgKo6RRjZharC6KkW4n8DSaZ
QIzyOCwxUe9la5sBCvzZbW1ffquvbXxAYpAqLp7R5txlxL/wZ/nDPor81rsq
qveJB60hZm3YluOyvVyTqWRjwd62UXQi6FKTE3QE0vgbwhV9p5HTnDC5nkpZ
S3A7gXq8w8b8vDElZj6IEfhvokOwWvoYZ4VnHcw8PuPQ9znH+o5fzL1iCLVM
9M4R7eqX4oy4BOXL3Qzr2yX/oM5KAbsqevvDLI0hF3n1SbzbGJ8C/T/iYugo
/8hgvQrE5R5majJxnd9OQtzvn/hZ3N7OMTxhg/UsVx0t3xv/znEF4BqFg6FA
nNbXcAo7Vh+nLO0arv/znkgW6V5fQ3cBELPMj582nPWPXoLDI7DcIZjX1G3C
/LGz/kOnEU+BHpmoeSY6+ZQdOkZKkM6UnYaFacAKLl5bOb3eEBRPtnyNmDJ+
bTWfkwxxynNdQM+aBKTu4MsuuDfoi9UtY7fHH95B/DKvfapaQAt1k+nZ88yd
U4xG+a9vVjHci3TVIYAtE1VS6GX+afL7RH/9PatJ1Pgt7rl+wtA3uyvLf/Ma
cBhp2nFk5MqQVsTuCHcz9Inavg3/YCKo+NIEf0jvT1TbYv82gubK+dBMqdZu
zoJtfYThPFZdj951oila3dVhBcwNwT28+U4bBoN2tR/LHRDTitGW1O7bR4O3
E65lrg4isS01+ru/Tx8NAO62n0FhdOmwD8uOKMhxCLWjEV6Pa9XzPRJBGP//
xqcYoiizN6C1+k5hY+VXwSDrkOXIg2kND02ijo+n9qqZjgpCFF+wO4WZQjYD
lqdsPfBi0caVgv35uIc8p4Fh8vEwln0r5dxaMeCxB3Pjy6lqTZTMt9oRDlP5
cSgutgCJLgrtjg335JtMtELHIPnclS4BzrU6Dk9mPdnxZLfMfUPOy8uKqp1f
a6tuAolidG06xHAKLiHqpA/WtxuPxDovd3jCk6g+c0ZxBC8PYscBIEahpsnz
6LPS7OmbcrUewf9HB5TAG6uTd+144m/c2cxPRWlkHWupx6MT3sTYnLzz/7V6
++u2M33w1f7TmteNqPY3mYNEcacVFLPfjLTpAkVJGfae/D57tu9gbtIFEuI1
QVWveZZSiqgQCFBKc6UdK27cnFZEGyUaXsyLlNshLg+PfY0sHxG8mQMTCDB+
ykOeB/RQalPqp3w5iirZ1mGL7ph0aPHc9J052yS3yuIlzpf0+5r0HQUQhKNl
V6w8h+LU3eVbs03mikOkdtrR5AWI9LPnuiYu8cRp2TtUPvhcYCTimOuO+NAA
oiVPDR5yf4DTjqs1iqFnKgIVhH4w7GMz003OHvKTgvxt+jeHIFLJB0mcinqL
+5egm4hHkdhUcEYthwmkz4wBhjIDi1lIvD0A9vTvTKzGjODGoT700OKYFXzJ
cv9pq5Cd3KHc2lyjtNTj5Wy//lY7yGjzvyTBdmOl9tsgu7KhAFl5Q5ldV6Dp
fLJOZ6uEsHm0JUxgcrxD1igzDEVFan+tvM1TEXD5s2qKa/LFgv2AGs4CAI/U
hazOfHjWiHVVTuUtP6BRnOumAQAfJE5Om3d5A6c3XMoDUAYUdKNt/2kwD39Q
2WAlTPGszQhYyspgJ0nlE+mj35xz5+HFg73dV1Xh/6MOpbak18GR1A2l1/yi
hCI6Fa3IWunQ440LRanRRJLqsJxKDfLnaR2vNKGA0aeBMYI16cxsYSpu2VVv
OcuKacsmIP2XI3Ei/eEiEGiSdECKomEnP28qTCNtLQC7mjdahufQ1pV3Syu0
hskoggvM5kdTPZV1YVPxlu3lfB1As0NNe/UB6Z5AmC2YWMEZhlY/DVnYWONw
7e5/iW9+kf4AX4w9VsRfOIPA6OvqQ8GI18XcG8h/zYSg9BSm94uIxdok7jvw
yKusrKgklS02hbFKggMi3yM3RRplmOHMKyWMLt8f4D2Dekgt4lWqeZtGgZPB
IAKNSh9SyyaIQGocxMfPLnnIvw1j1Eed3zArAEXgUecVCBUa8g5D6zJXDdFq
UxHjBOBfQ3GxqfUzXU+8PEmd34cvVSOJB3AFTN/grOPoH49yrG/EcHCkvLVa
Kt+Re2GGkLP8XGgG8F8bJkf04fZxzpJJj41JxGXvvH49/oCB/7elryY1fC8h
1ecqcNQFRbk0BLvBLsrNYlN+r91B97pEBVlAfO1XU2kVtFIXr6++/8FIJabb
g/TwUby6kMBH/hMiIpw22+fhcBTmTfTZetn7DU0prDUc+nPrV7t2hYcXEBxP
dqsZ2OywZlHqeTDtNaJQL0Q2sS4RcI/DTQS9I97RV1ObZX2aaoccOGbXw32w
SP0EDJyRMCgZXCOxfmbyFmnP9aOoiNKIKz0bpDJkRGv3/C+NijXj/iVQHRyN
eNs/X5vRRcI8LvL8JGmAo645H2kWU1xggH5JtLVsDAIkBGEl74R3YgaBGnf6
vNEGEJhr/EIGO1oplhPeWtLgXJOx9DVgEoXysPH9hD1KfKlCMh8cY8S1RQ0x
65SFtc+YCRC52ChaKPD2Pvpov95/DzpjtVuucwGaq2032tvM8GG1AEwv0KJ4
OJNQnwsmoe7qiY4pvtqB9Kbhmnj81d1hm1FVL1QhGejHh3WTaq9eOJB7XON6
M4Q4J/qXK9hyY5dCsrIFHKBob4+dagT8ODkdrW5e2XusPl0Ob3wuphW+SFkp
o8Nn9taYPz6YH2S8sKAkeEhh4HWmEUuR8QTSRJp/9c3W7LB2aUXNzbPElPzX
unoKTpDyjdsYefeUOE3+L7s0j8VAxHujZBT5RUIoesGfpshakDVFbWYrqhaA
C97b4+43tlP8IzhkcSJWJ30/DdWj/CXU54mK1vPrUlBkix4kpc5mKiv2V4K9
kbR+MVx/Xg/5nKgIPmV/+7iF8SVBWfiyjKE5il1ubtewCwdqYqvBuP1SM01K
VGOYOO5qH86PA/59XRzhCwFE43dmpIpw+TyWm7PHkmJua2e9+a4v7wjSdhEe
EsrxAAvc6IKkeM38/2fZTsWNmpgHZ37p6pQka8kBOpVsJAZbY+ww8cc/BuX3
UH2KGR1rwtlzMPPXR40Zg7L7ELm6usP25j/oQjsJbpPMWsA2cOQ6scujEKoX
YLb372LCvnAtJelGnGtDSmycGWc77V2WmkDk+ovv3V6KDYpf6kE2AD2hmvJd
RrnV9XA+UYVC9U2FqaB5yxMuTbgAAndHgDX6qqvKsPu1vlbn7ErdpQ1qNPy2
BmZrGN4AIlflMcSKqlODOcLmiZkqdLsdffJnnzguwfHkVMKRFuyfpkR/eGSd
FvlQGhceV/kHbZjr8Ch/TSpMj3ZOX3nU0zsFbpm9078N00hLobqxvwAPPJAA
Fki7k9oaz/G11fL4uiF7Ka27tvvrdlktHarrEs3RFdbbkKWCOZacM8zASW4O
FyTfKRaHSA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqfdJCIGdA9kJ9YakhewEd5FC9jzvQL7IyXwpv9yaMlcWS5yO8b8TZo828SX4+Vs8dC/QQNAqDIEyzLUjJXzR8SYbjEWeMLXm99F5BNW0b8EiEfwBz60PBF3Kc2B/jg/0wTdc2uiFSEVWJlc0ARx/e2EZTwbB+1VYL/7qZj5newkcPAIzBHm+NAFuR1G72kcQCrsOYofTXaL5kiEJ9pVFhdsksyjIZACADCbVd4zEK9YYztB/mCQCgsQIssqbH3+SS2ZWuFX1CGP6m6S0HhjthqFxl8MRv29qgCKll/qmR4Bh1JQ6DzdnTpb2DSBZIEnf1GnqRwQwTxZqfmENrRp3fAmKhiYkUkSQS+9V4OSgt+Aivqye1ajxwcQYeXO0vjuVWH367HrSzAJbkz3nS3Tv0gmLm94j075oCp/HPuYf6k9ci1LLbRhJ9M3omMz+tqIgw0SXM8U+UWl94+Hz5/ZKFEUigqQ1btx4bW6jFz/Wg8rrTBiGMqWn+LdyA6qJa94A4L1BNEqm2nEXC8rMlevbWcGr8396CFG3jEl8QVRWSwPPRWgmNW7kGf1BWfrPAlkVAKp2WzezD6UMbwisPfKAdFBOhKLbvh95aymKS0M5srZxZ2M6a73Sx/tArIx4iCSzSRazgYYakY+jeGNznPN5q3S6m75CCz2nX4PRjZcLSPv5nHDOMX5ZIf9hQzUgZmsxYWy9lupOXWcLHTPeiP0vNZDxQqTVUT0T7g7wlXAZO2c3sejsGJwuKpjrffOSC3KrAQR90gJq2IAHxfD1t71ScYn"
`endif