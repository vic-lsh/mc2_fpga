// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
k0P1xB5+cIF5geSTOX9io8MyT2LMzW1tS9YWO38mbjJ8MADLjKdaJx2bouTV
z/6dcQydjBRrtfpiUotlwZPy9OfIzQudPvXDmIWao/dqmCDBcW2Gw6/50gN+
LeB7eUSzugnZxCZaTvFfnefrOk8vEBxSztwJ3i/+D68TpZGihhSLF8UOOkHh
qLwFuWBQiLBR8YnkVu45tAhgLSm/pMsqehMTDa43mGPUSf6GpRKK+sPzBvH3
FAYNt1DSssKcn1s7a+PZlm0AL0x0bYTKoN/DJ9jFMrup+a4RyRi1oI6N7eHJ
g+rYHxtGtgD4hT56cKhftjy2HHJXa3PlICW8h7awbg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SRBR2NMCYsnj62qvE0RaCqTbfxxxRiTc59tvgzs9T9wtiuGm2zmejDsdYqS0
WiCUySya/rY+HiY7KUgXdPB3Mvp4svm8oeZ8dlSnFrRtD4Hsf24lQPfpYp5C
791OJTLyLEa1ZEAmJvna/2zJSOvuwME1hXOPxBFiVoKJ4LFnCwycCmCKbt1/
t3zS7qHhdkClmQhE9CcF2yeR6Rq8X+osWwhGfQJ/gbExvLYa9OFbvDLSlOVV
63Lzmg1h5AJtSdSDRNDtUt3IHvAKOlINiOPks90KRKGdqgSX5sZ13nrvwGCo
uE3cCxctTtmQo7PHSjFBVUydb8vq13ts1Y39jT8wZw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
l0cVVq9yfHU2fzVOATVMik1LUDbS/cmUTROMQS0Ja5KmRiguoXiqVln9PzlV
X/zvPcHXhzq5X2UmFE7Tj5Y9CEgKTBXPX4OcmXDyfdmoP6CIUccwTvkPCvyi
kCJFXwqUPC02gsWh/AmKRMfX/1jHDSbTEZyT6tN1DmqHk7KaWxdTEEfYBBsc
Z2I7TyCpDsODFpQ7w86ELSsiMupLmgXwx1oHiTb/cdFLDCCDLXQcGCRgLGYd
QIeyBHTbjcOP20jSPNZEz8VGk1i86ewcCi1I24agdPXpFYI+ZEdi+tG2HAvK
CdCfHBVbMukt7r4xTQpCYyhE6OEskzRa9VEbFIPIPw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VLUe5IYbrZKZ/6hpxp75/94Tkxrb8Q0KjmLGhi3/E2RQNeo13jnQOR+yhYCv
Q3Jdh41xBTVo4NZZ3e8/4ZVrh2JO0imyln3axjyzKnaOCcNAJepQyk//lAlC
uae07b2ef7cwHQGPv6cOa7t7CliNImqSilrwhoRG9J96EBxY7Ij14zdpVEl+
qUdPVRra/HI49jkA+ULT4XDZj2oNswByd7F+LJCfwR14insIvZOhFOhfUV9S
4CuZhO2szPs/iyra4nsuLsjK1MjG5itx5ZtBy1EczmPhEjPJoOa8pmUM3b2i
MpE+VIla3CLrdLQ0SbwHNMOhONQ/YpewVvOrTkOFXQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B6/o+TDJftEyaNt+0iKLl/UleyEMAmD7m52a+OrfNb4e7J+dfdTa4yOVconG
9urTPbyWsAUTtpvJaZM7FzB4EG+5PMU8X8PZq6q+4XDQr/BhRGIFDE+zp+jt
izUXgY4Tk8c/Z5iNphY6e9/3R1RsgES6oV3zEHcBtUv0mnAA8Cw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
bizgnfvomDO0JMR5Y7q/NTB+nK1hI8ayOpZglTrQjlG15fvpzSMkQKpuy0P3
ZApTyZ3RwFIhKAA43scIS2fmqUzNEaVzWJ6lEql4jfXzPo1h8j0PW6JBQ8ob
WQeOoxvdy2hp5EwFK/bR9yTgnKozw380gGbI3gBwbFeXnRetvU8ES/UgY1hA
Dc+cspuWgFp5SWfAMsQu4g8AphkQRrcysxxfOfwDTywQDaHCK8DGFf8dBf0y
NUyeYOgzJAikmo7udfuKqNH9cn5ptMtFpK0fKyXFUsCzLXsg7OChTdJ5iq9U
IKllHQJ7t+DyombkazJUgccKomSqUB+qJ6EdNTatyp1pc7Yyezs931/JSHwz
dphRkJiy2aHRwoBpviijvPAW6VH3tt1744avuX6OSNUGOIaibI8X0YMF4LBb
2CL5xU6BEwllQHT919TvAszd0HiWZKwtoo5+tI7Ubx6jgcX3jsib/G/qmv8F
VuxqcLgVEq1eurQPKyzdPPvICWSqUUo8


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nBY6/2MIgdcj73mWsz8pM5ZMvBr9wG4JMX4nrTDHC14N0cVSRiBH9YeIMVaS
0mwBh2hux4r+KkaPmfCeqJCU431O0+PL3zOrvZNdfQ8vN6pHOmUKLdEMKNa5
QF7S+ukmNnzj3cWPcF/nb9s1H+4MGX/Jz1Iq32cMZ0HIaMEHPIE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
n1feRU7LZ0Awdr2H1TAirwSHGakMVjyww5RbwNsgEBdcj9S/NnlgEzMsu/m8
6G72sUIZSqbFlyfrsO4+no4HsRbIyYbCHIkdIWk8eRvVdio/baWvUSaaKWtw
iC1V82fCkLi4ANHrh3xI4kXQixXo9hEP+GwELSO8DgWGfwcsbsc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1312)
`pragma protect data_block
ZqEdSH3WU4ZoqBAmPjHy8NN7K0anj02NDOhIsIKmcAyfLa5zAA3oTTgz2QKQ
cIhcvnIxYwFcwj9qKLKI0T+wo1yLPIaB59aQTWv48s4L8aOE3ZYP3DVWPfSa
Xt1qSMwsAtS59pWxVmZsuTuD6Ud2/+ru9mCIg+qw12Owb+/U/9TwfZMbBIbX
nw+1W3WEuawAL2NNIhSVy2TjMCtn+4aKDg6ltWgbBDacEEc8LUpqK9c8K7zs
Mjmz0iSOLKWJLLBp1CsPgc3V1d4Qucm8iKITcC9GfW1EBZzIypLkZiwemiH1
uLms7mhGHNkOvrR4mPY+xwguzGpQkdthFmDz3NeG7ZKzlozc3En6B+is5BsW
zXo7SVUmuU24DxqKbJ24Ky7mbs4tBR8xopTKgztxJ6n8iWMvV8I/H6El2I+a
4X3p6/T8cZ9Tcipcfu5rJVZ2DS5e/5Ryt9xNBSiYcfSXTI8QlbZcJjzRL4YK
kzpk7cem2QP3SNox5lWo/2d7B1W0iOg70zjDuvAb727jClvCBXl5IvIjVZnK
FPWLzYG5ztan6KKn3JdZwe/H15rP0nytHk0YJfiet6egm6J/QJ1sMW2lHGQn
b6q8cFHP2OfwSVHQlJyvoVxGFryIZeCT/Faww09ynMP5kR1bX28Q8lOJe3at
MbvDk6ebYc5WsAwC2yQpD9625tjRg+fbAwBPXwKj6iiIrDXoNBE53J5K4wid
/qy1P04eQvZbQtMqlAOegkzeAXF8psX7gGtJJQY6jxXWEhG4FN/DvJbODOvp
fTCRgrPoG2eonYUAp3fOBZTIjjjOM475RDlV0cdvrJvfWvVbz+xYFysc+qq0
1Ig1WSckKFxSqEcuyoW/BhZuvSwKOH2WF9MN+AvhHiCZAA+e2iadO9TA3Agy
N+EAxHpzxNM4PvwuRWPFF3LSrlVWAjimmFvlifaR2E3NHg74WyxF1MMNeKmN
htCvFeETjiNzWsea7XjmJvLpOKG/dYq8PAfRrZf1yKGgIaEs3i6265tRkWlj
cBMSbr3Sr7rt2TCdb9HI90Q+hmY+tGqCUdAByTXevn4Aq7YASfowZdwHX887
NmgdQ5e2hGM5BPRwZVH0/rGmDGqQ52XKv/FXPizRfz6QD7XJwP/iAx5PURhK
DEq7tt5O6aUib1oXrSKgr0yhr9Fr06x4v9vVH068usoYLgQ8rljujaNuCWHj
lIln267M+j+Zc1MknGuCa/Iqazxv+vX79y9y4EGcLIXN50eyX47431rdiOqh
r7AffXpu1v2C/XNqBczMUanJyooNuZGrPT8FJll7LS4XOJk1Es1QCgnJjowQ
xwz4ZYrsguexmmkG4BxsxAln4Si0l5bEvsIlcwnFej+rJBL610nu85FFO5Fh
TepQssqau6H5euCAm2MIoL4XzMcFIHcm5SGnkkiG8PJeBdSSYAOF29HhMdbd
rsIqWmKkW2SxyNW7Le7UIZa63rMDJc1dj6pO4+Op34xZD6d9O7+rvqL9l2gb
9pPP223E63TEQpkrnNcpA/3yjgwE3yF8qdI4LdU4OIBgBI9Rjetz9czU0lWA
fAr0434MVGgSXZGH/LFBW98i3aD7h5nR9NRxefocXwosed5YVudsTbg9tZqq
6j9d7pctc9GWl2w5ifyPNkVuX4fHqiN7PFPpmvTzeY54TqspOqsgSVOc0df7
PbUM7yzHq5kIVlJmJEJe+EL/YhCLYSup1SVI8Omf1CG6RqAv6bloI+8Gf98j
Rwu/h0n1mg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQozScqX01C8r7rckxvVm4Y0UCRif1QuvmitGV07nqN3LWtB1tGNuQFzGjaa8HNhH92XU/22JOWU8TFDv1i6OMjBz8kcxwOnG/qvtoDmtTT+S/y4nwnZlYpg9EzofmvQxx+xbDV7rep3xV3Lvp8Gj1nitvfsyvj2f1F/kCM8K76e0Yk0vCf/MUsMQXxysS+4CXmLvyyuZHKTZfJur4ba9n+L9+Kq22hS1CrMr8jxrQe+2DBUEPIufnOwXKiJZEEG+7n2ig2zt1iistr+MQdla9UhzIkHHQVfalfjPP5wfTHVOjNrZ3kSfe6WvBP1jeK73qg0pujAO237X5tHvUKrAPKyDa8ienAFMUDlerzjrdQZLdWl1Nxdf3NM9asX8e6Cg6zq8CaIrL1kKCfo7lf2Oi6nE85GBotdBvidYHsHEko39rVY6mM/rJeE83ZDst9XW+aN1zAVhBgoLGoEomSDV18560gDRr+OLvK4F9TpLdu9XOI5kTs/f3kBQQ0lOV4lF/MIEnUysVEj6mUDJye6e+OH3DkcgG4ieMT/tNdKcRrDDwCJR7K0xJJh5aPTyF5ZBoH4wXt4jxPFhjwW9lv8n9QX+NBXrS0NCBx1nFZ0KMZ6va4+NV8sRIA7TJESlPEe4iBvPmOk1ckAGHXYvLVjnEiVzYA9A98rxoXVsjYL2LqFs2zAgobUHWS5WSn5vSyGazXp7XJt4ptvhi8Mmky0bthiPocowghs3n3yLkFCIFW6fns23WeUT25CwL3F4Ok5/6NiHTldd0ZlkBR1DmLHSX7kZ"
`endif