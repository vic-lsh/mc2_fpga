// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GoO8mb5iP0Bmh5qHSVAiQB7amo23NcEqREYkovXPOzA735MjK0cH5wAo5ucT
7jnVzVelqPIlFPJLTrVgM7CLwSHvMAsX4EDbI0CasH0NfWEpO6G+mBmSopG9
wTvhJzRSjbow0+5wNeEebVbbYwdTMeSkliXA7paO4kY58BIPeeEZ3k+rcpXj
bHr+cjUFpj7BXKSf3WupQdIswg+WUrhdIGiJQnRptdd5/L2z4WDZuegw+rdV
zojodECjmO90hv5LVFVaHmlhAGqWYAqw+P905ZCtAaSPtCy/po/L4GbTyi81
FijD08LupWy2jmWilkVpdzqFADLVxRi1tWu5YyfpzQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QbcyMMV7Q3y2SSxSHbw8hESOqYEiGDzhNFlmWJPvpD+ErfTWmim83/FnTyVZ
u2u175wzJYqz48Tww7DGH7z0ip7CAKgxlYrd29Rlk74NkYZEd3sKBRYC6YIi
WiiOUjpgw+KgslPhWEGhIvzSRzbtCvvO7w8pg9LUWCTi3SqgnWLgLj7/xBIX
vtcGKxXSd+Ss77jypDAeDAel0E/j7iJgPJO0/TYjJkKFWjyS5z6HbKito0pM
o1KfxMUkFQ1nBzqtEce1NAEQvgps9MdDjYr6Bc/sm36NWgyHUxbIWgRoTVU6
7XVPbjXU2kXpiorGNUnbegGBj2tkB8+/Oe0jbHV3rQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rt6oEi9ampadGA6skjp+4RPmXjIdmKsI50iAeQqXmamhWu4/0Id59/4L9U2X
ZX3VKJ2qNNsIq9whnnAiCj32UQcXII72PC+Cw7CQCalhh16Um9pV20F/Ub+7
8kUpQh0L1rR1yn91cAc5CJTM23DXsOo3xEWcX710D9wpzjY1GcYWSyUs/MOE
59x9C9Hq5YDgKFbuml8t/MW7AxH8w2P8DLUj7FHsEgmiS1kZsY8cv/KDrFTu
7zWg+bt+/qEQZSishNidPvd0VuSLTHeH/AdRmaBF/PuOFPiWHOPCCJz/nRFt
IP4+oWsv4/yYUXWMPjO/0OQ8Oc92NFh18OSTx9DhtQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
X7CHV6rm8BnvMIntZPLZDQ/b6KtcuVegnzLB6rlSUzppVGBm72t2a6UNWdQp
iqQi8vEnrG8C6hTIS8KMMacz7mFjCKUWouJsb8OrYiTRlbLibDyKj8zcgLVn
Wgclb1mSWpmyz0jNJDeQx6dfRJpHIzg/CvceCNgv/Zw0Dqd6dhWbBaETAWtA
9+c+3l5KT+GwrxO6ppCM+fgIadHtQXafyCnSQoHJ+x2D8Fc4Vc+Dy5fOTLUe
Rd7GcOdtfcyRcQDm9CbSPJha6VJJ+S4dy3Iem7mHqwKT3RGgHWKSjKfXtUsF
DS2pJP6GSs5UaxVNhk4lrP19TA/KhAxlO8NQpdWFaA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WHnjCPpfNHOX+8lfmSE+IcHKAoMfJzzfJQgZYH1GrqZiScPYVAMj6J4GH3QQ
6QTx92gI0OFHHrrA/tQCl+TKdNUoQJkztM69TEhVZGfCQsQvjSa15yeMZNbg
f+/7XL/5Kik12KToO3hioObVuwm3yfu+XkYXMKkGY5KBEAd1LSo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
UKtzhn/EmGfwtU5FkoffK2tWUfGCTMGjOGBF1cav1DCjkyFh4p+O0LTMIR+f
ihrqbMO1QgjyREJz3nejJxHWs1n0qyC3xUrumLI0g7S90nFXKcPxGlwmMMl/
/JU2qqyi6XoDeNI5xup3yWmSYeGKi6dNDchu0lg8EJsY1gH0Y1HcPxYFb7/x
RLtD6iJg7OmaXJflRIfVOvoMs3rnpOmb4SKDYGz2n73WbasnhSjfAQkBKN3H
+aL1c1FXxggdzkbxNU0gNMNrG9TnR3kueMIYB2NrHBDcBC/pTgFfIHpSguGD
ea/lmpbGAg/y0TmjTkMB60IaQ30qIDNRxoVxpJm3RlmbBanLsJB03rpQh7A9
6N7SD7y1UYLDMl5CejggJNJ6hjxkPSGpB0HDaPAeU2ZDKP1r4EF/0Y4Bn5yi
BiVifTfmlG5o2YHC4djx7OXK80Xn+4l/ZzbXQ8to3u8zUwY3Nav3VKsOTgdy
bX4FRA3uFL6TWAKLM7mO5UxWG0BMFSye


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sWgUkGoSEXw9MmJZiOGWa6wuDumfc8XJpOKnAoO20j/yLoJniGhAhRS1mKGp
PJ0CagqLjekkhhnbe01EqC8yV+lEGjFBe1N5mF4o1S9yjds/11vRNY4e50v/
JnMaSM9pr/PBpR18L0N0yzNjLIUK4mS5lTBK/0EBBzWeJ7DF44k=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qdNk/QNcgao9fM37cPbgZrgO+dIZ2uw8nQtp2uokOHME4QzwH4J1fXYgITMo
6JISAjr3fXvGndhoTDD30AD24Xqc1Azho7mUG2BSav/7BM02ccafBUijJMKx
d1Utn67RDKblF1A9EaVtj3SuDdQGKD92yO2Ig8weR+OANtfUrJQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4304)
`pragma protect data_block
mlpeHV+zNRNdMS0nMbCJ8DBondNFm2ZH1lqrjML/PpSFY97z8R5FbRSdHoQa
Ay/Op9J8P8dHKHVoRwoJgPrhmMFtiPwIozoQR2TdgmnnMuPv17Z+afMBq64l
20ED/dYLSwzmHliijugpdbioHkCaigG2kXRtigJyhANJ7dNITcEBgVtaRxSu
CgNB5l7j3NcTOKqheRKA6iMvgze8IbR//aDgbzWLExEF8J36mpy//Clh01Us
jiM6OLFMpDZ1mTdSa/+j8YhTAeA0MYXzPfLlWeJUZGVUQW4LncE5bGD01DMn
bvwTNstgcqLfy9bV4tImTJqCmBgHGJLY0JDAucTlOvg5Wnf8KX0iyUwyj9+o
DRJu04ABCx15jchpOYReJ3opW/Yo55Zs+iFrDMwMFe4WHQLYYYTzgEpt4d3Y
6IWdWjkigHHry9KuVwQEHq65Vp/ItOo74c/UjMT3b/djR+mBKov4EOj2IU1M
ix7oNRUI+TcxzX3JK9GuGKGvSqoxmaQ5DLrLjvapQFOD8cDpdIHfZMY0JGqf
jvOwGw2vEIegARd9rvGBNl7DdRV1K/hRWcy5LsuY0IScQznHvMNOqdgqm7nP
AudLUUQPsoZFIA11eRWmF56FxjnAa9sAnD4JYgR3z5/TkJf+AzufaqGEvloz
SyML0DrF2XVgWIIZ+YKbXv826/2vKR3thnRe91IYo4m/xjmbULNWZaB2Ve+/
0cYe5EQV3srNSq6xLhkClRfZrYz2HKL/wBQ6A7o7y1YEzLyUwvOkdFkOd/1i
oQezzDobkHZMtAVLuQYF+4cwXwTo+KpRg5KLNqzePcqS9SrSIpON1IGbns9v
mr2POTiXeHKpwp+Sw/r/VoDTU/4wAjkpwh6KoVnjXkkfNEuc0KsvYGagOIO/
uhYuINywLMFwCPsLbCk39e+JNOlQ954btQgA1gnLTLaht6U4hDNqglPpWFDU
1fZpWARkHJ0B36GbLjKIOwKkEqRIZvAoSxHz4yLr068uPtufLsmxpW65e9U+
Rk1cgQl0j4qef6Cd6i9OrO8DPuMWT4mh51p+lrjfKeIRBTjh3MVotmSlLp4u
YSenr4t5pgmTFuUYsJFvJNUe+inUxi7My0K9wPNnHsoGWcZX4c/jXVxUDH+t
B/SCixmPmcgkEwqzK2Ax+G1/ldaSHWWh6q2KmXHxp7uBnu+8Y8yjR+n6NgA9
Umc+dSEPjtm/+5HqM+KMoO/kR3lbpvYLpkcv6KIyPBAuZUrLaplapKfxQFl/
HoOCRq8DAvo2pYJOW5R0jxByOi2zstHpfu5u4uAcmYk0q0Bhww/3hldbegKU
fdYlm8Phu5fG6umcREMuhqmtDgj1HU+V6PA8hZHu7hR/2wwuisJxitbYTSUr
94j+AjqL0d8EjkrOFrdEDy7b1bscGoVHTeNhCry3QRRZCxuUYGUjd3rSDxtZ
HWoBbCbwW05WUtPbHIkpPe3IyJQRu4JokwIHrqoP/58JyZxyHtrTMEkPxS58
DYuCMHmbT6MUO/IxSKV2q3nhlukLITrwpwoAu9IwpO44qzOB8cwjh3rQDMXV
OToY3M3rCiv34dABbwm88QZ05Cw0qFsA1w8MnhelNj29v+TmugKAcsm5fdlR
BIowszW4faNViil/xIeF1VGWnU6Z9qihzOgrL+6bfCJ+T7KKmUgCP+vtI6rf
V7FO7vvRednLs1P0EscgZdWPXYEZZQ/L0ns3SW5TFwGv8VXrDT3eaq1QudFt
ftCSby3gKozlrndZ2ojyg1k/klMxqwyN8bNOLmERCFeaKetYymQromRqrsKQ
9hQv51Ik5k1Xb0NLN71VU2rFn4NTetmjRlbWgwZqwmNGz1ERK8KU8/33Dbge
RpWDw2octcW9eH2FjimV+FNGvJ4KPv8G8DybV1LPER8l9GyZMfkBMczlNO35
5FD/Es6/QvLtDul0OuDkcYNdh8BOXejI6/XhrqtiN0r4yyyeKgEt0xRfv84y
pZNJYZC21+sjqVe1BhhrFOC3gbl2ISVzJZ6r1Iv7MQuMCCThX1lxoCOBmUTI
bJWCcTTWtEe/DnrQJ376gnH2lhz+nPAO6R4riy5CqVhOvhJH/xvX9I7Az3//
4kvWvQklJqoiFH1tqECIfMPwLbpTcn6cFvfREwoCeiEZFfPbcNLSEnYjz02i
Gq/x57TBzXCUS0CFsHxDKi44+U/3zuFtCrc7loVuy+EXoJspFXTi4G6GHkHt
UdWgBc/oKaItxH9+IN3gOC7F7NaIx/E2lu341ZzreNV60pH7XQqtO2WyFhtk
ZQyMkdGYVIDpVZNaYb0EsSZjH/uAp/lbRXdaU4SitH6ndIL6k6+ffXD1roo5
Z2fdUIkMooCKGR+EZfLYeBhZUCREW4JjNlRtK9fAm6VCA9qSj1kSNn60h+GP
7F39nc3Bqs4dHfa1weWO/+01aqHrpjJr+mUso7ItT+FIVd+RClYTrp9Z2RaZ
l4CWKAJijiR9+ZyWNh5N/gWFihiVS3kVSbLQDA692ByMIHKHluhDyEVKWkA3
LY2n4n04+Cb5flXFAUhlPyiV8kUuOkMFDANxM3hNx+Npzm9ETC8DhYl04wB2
TleG6i5jRbR2l0zqNPjoCD27VpbNHtOoAe/jdvEmcixu3Rkpj+gjzDMtrelx
PCoWUM+iuHokZmrwew8yDQ4XCOPxjuRY0EFv+6UTUBTHTj/v4xLeXwGKF7Fe
Evm7blNvw+vx98aiUqa/ShHc19ruI63+c0n8zSkxx2JNtknWWUWOri5aWb91
jERLuIPpbMIBF9wmx/jNs9YTi/xHoZa+G1FLVYQg3n0YvH9SBoPs8Ad6ZgfQ
pcyGk93HPo91JUmb732ywucwRImdI66oD1vNp02ElusB+pHXPkUKEWFhDAq3
/wHKKxOEp/xVlju8jYHqYzdk3zJKOvQ1yrt7HSmE58+qrrewmUMz/L0z9grV
wdoQ8O5cMTgJbSsPxdgQTTq+Def7+tR9PVZPtn5kfhlJAfban3VLySj4CCuo
wX44AoQwuL/QRZ7LQFkXNsxQj9dYGMIvBReKIiqQ6Ip/pGOOeDTLosITME6e
i5+S36HmuGUK4twkYyQibQFlAmAYG8NWARE5iz5Fy5kD5+epkXDpVR8ra8/I
4ctXwakUtAc3GsK7OGOhLRLWKm5vMAEPqkRXjGa3PssWM9a8hI62zXwvjWYq
Q9f4w+4ltahnHOtpmxdfEbs9CaAPlN2lvOsEZWGlcSlCC0fFZ/ZlPeCtFSsU
9qYAnjl66bXJHF9c+ZDPCHzE+I2gbFTBd55iyzqB/Rqrqeu3PpZH/rB6MjK/
v5TH0eZvlyXSykrM5IkXJMFJb7YaO1sMlJDQt2JeiwGFj7hYzypULoA6HdBB
pVOIgBf93QCFq2orQQ0dL9LwCr0cZ7fxZ3jtTJI+dBMSeyZs/Rfo/9cOVe49
8LswzpR7ji4xoyuc/HI917td/uJe5BuBGWKrh6jd6xiA3XLzkzIbeY5bF41D
hLOagfb9MVnIg/xsrsqiDvnCkwCxPkvpWx5dnerhs50nQMwIg1C05IOGaNnz
A7OwTE8UyVQWkh6hNkDMo1A4cCZ/L6pQtRCe2WvQnfSjV/wDBnCtJ30/XMfo
FxdfZXwEu47y0JiL85fcF38QBipIe+inq6d87hx9c9Db4x0RlpnaN0tC/Ws4
v82Pge2aJUxeUq37KFFWrAZGmNnew0bysgFlaX6uiom2hO89qPkCq6o5modT
e8qHCr7J58UBZuqwRKdPSQT9PuUtgFqoXId1tIF7+qfEVmy+m4ktWDzMvLPM
ZWqaFN5lgY8JrOKD+8iooMML7nXfD7sd7AuB3BNC11iZBr8PZQEAU5EG29/0
mSkY8c7QWKceLl49u/soQFSbG4Na4rQ/WMxkF5NmMSme4NZnvKn2rgFMcBj3
m/MG9Abd88Ma4htaSkJiPNoqTym0JKeyuRY5XUhl7cHTGE/ztWJd5YmTrg19
4BW9k1RfaAp9l3ze8n1g4OmHO1/SVfIFQWd/GiTxKSV4bOOB/aqFWNgAP3xI
m4cUngXqvUBw5Pv2ktMVxmUzFnO6749MkdKlF92YhTyYOq+wPxPZI1mZbDGQ
3fxO/9c//hJfCcDWHBdluHK8GcbPzwjKJZtI6Ds4kxuFUD23ksMjmn7shOxz
loV8EnBfUEl8SetuI+Q/Lb2mU8wn2KK0jfxGiuf6V4So4hqBTC9EFcqxp/7Y
c3C39gsd1Pzxw64y4oM+LAcg8GTeVaBTmu70nOv8WB2r/TTnhmKJvMKeQuAp
MX791p8U1OjbGBSooJ1kEf7HGw9EyprCeq6L5X1vy6EnjE7a98OjcE0uC3Pf
97qxLiMB3qXKVABkSttzpqwUpFHcZ1gLKkHxdI8oGPu+13xOELXdHIyK2QvS
/6aGspb+gHpVYg885Wq85Xq8yVoaOLBa92jfWNLOofhNL0jmmKUTTd6UftCq
8AM0KYG1gv3IGugyRNSrAziAWVMeahtWnvrmQ57sNjR9PovqwH8nq3wgLROS
rc1IbPDRoq2ecoyOR4mGFi0qJivJhWTec+Cx5MZE8FsPhJK11N/CdmLevW81
lcs8Q+nM0T6/8S6g0xv4DBJOkovLztEOClgvHwMZOsf6xYShk2u+KMU98zjY
wVlwv+Y99CIMKcSICFoitk6IcPWqRgRJsvDcjbpZL0whd23W69GGhUDu4cCf
dMxB6AHqlQ2+B1+BJf9Sue3deAM8/YnTNUKGEpCkr3Of4eIXtMmkhyMFl0Ph
tc875rqz2H3l6VKN7/gjHEg96rBvN8bXzgJIRsa8ZwpzLnF/9cts89xjS+Cc
psb6BmYbX0hesDfMpfrJulBs6MAE8raUtjR6FCplOOqppsL80qx7v38GQC75
p/N8FSubmt/zO21pLLE2DFQWT558OGssnS6yKMHeqoy1ujv67IhUPIZUrxVL
LzRmGR2bb8vTA2xrNDqma/g2CWtKjopcdf6X2D/lXp8Dyk3VL50A3BTumRcI
AK5BwRjvJrDYskv2Q5WdT0RaWdUp9q+iQOZ8wEjW1NBcS0HTGXsDirlSxB6o
ItVo+nuLBni3soGnvYHI9djdmmvAji5M+htkgH3Dr4Oa/coR1IgrqDCL2txs
tDqU1+WT9Zfk39TD0Efg0jV3k+a/fuldtigf89T16llWrXTEEp7nY5UgzGhm
eq/zXAJGoiZsNkZxb6zVV5BY0jEzvzcPX8VSI5GeErVno0sTZDBh+YedJ4d3
mELUL/nF1bif14uuPyf3Ty7FmLOEr355ogDaUcKjVuTrLedYp9xkdzu90HQl
hhLVHFMbTP5kZXAXUUSfXyfEtzpQHBUX1h6hLr8mdnaX2XWxPvGyNhzGfn4N
+x/xXyMuTCYwdS5OqDt9wl7Lq3sjBy4XWgCHWnldZxt7kUtTK/CcOx83uBWn
yEWZXxIl8yO4SW3YN/+oXnS50ePCB2sMnIlQdvCSmYjRk/JoEgKLF24OXhMg
+VPE06jrh4G9eBq4uMMR5zyOiqO7JG0ZKN/WK6qSmI3QLOahFBzT5Q9rjLYC
ImZ8DlprHZHC82ACTNW37x58NYSHH70BDGUE5B6tl8PX79h6mILIw8IJX5+3
iFrxIT9yFX66qleaAW5POX5I2skFaudfQzk1ZpkP0IccpZgPtcAvuaBeUYGh
QZO94E5Pqoew+i2C41OPXt1HMhNWOlYzZhyYcESBksQjEalw5o53ox1O8kPc
kQCzUF5DABoTFM8yXhgPDFqBH8sSvMP7OAuaZdk=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "NwPt+Pgys2qG1idMcWv8Fn/297svhiG+0npDp+FwFsxSj2TABYEu74N3vkvrkU0VEe8n9svI1xYDwBf2JdHDR2Xk8uQfGlxUyZotzZFIL1qqzn5tz4d+vaxhnnX3wa47rFkby4BNmPYN7i+N470jAsZuxqIybK6HzK9na+1SravU1ZtvDCvP+0zlhBs3liCFGF2TfnRM1qRxSrpw1P5NDga8XELxExSCN3NlfsvRmyKEGi9FZwIUiRzyWgF5X/7LZx0BXYzTb9Y9Z63RoplM9zo29DrGQCIAoZPZqzH0Tvhkr6xLHranck0xUYJnsEicTTrRy18oxF6oCw9EBDeKWatC5y3BVJ9LpiN8Gq6+UqBZEsQohoILvhB+GHFal3GgJAKH6zjAtNaDod7486bYsipygmvgZdrkkYp1CGqCNo5Qdo9HKhdiQepFAejIORtW+rdiPyJZTTIV2AVeMtfz7XJbreELBfE19/i+d9RZEJKgmiQrubQoAFGb6PywyE5V6lpY+QFdrCfzkbOiZzZF+cd1HxNpi7QRpbBD8pgEU/1/uxZpQC4EDjzwT8b/Vo+KgxES9dcr2/XItlI1c3Cn3RE16hHGOKZIRQpg8sSSO2Ix5E8oBLRWoc7iif3E7rvFhvRfNDbDWmr3sUIUr4yjozxmsnslGyVcDImMOClxhhVCxzUPYbaeU1w6RDVUCrCipfDcy3+2k9KPqxlcR4/h+tehQTgQR/H/VicvdZ/q+bBFqJLBbXU1Gf+VI4hKW2h7xw8Z/Rx7Tap78OJrne8xO5H3OVjEYCo+2qJrEI3evzUXXSLu04HYrRQ5W9rkBOGtcWVuEubL5eKqLTFPT4Q22PBUSMqpHbbXCWO0QCLnXjxYX4R/ZdL7HzZgRWdpZffglJVbGFRRtOxW5zQWS6KcBd7a84YTU9Jcz1dzMc68UnAeF62QZ1PRFeLzEnAKYiIdBaMPbxiKxie/+KaLP48AEnvJDeD45eViQoaUl845bgtelQe+G0Rb1J8wI/X7dX06"
`endif