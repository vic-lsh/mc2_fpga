// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YX5iiDNKEtKy7ACAsbLepKN0awpyIxC/dU7IHQwEQ4x8ED+oLvrjsDFLMWtC
XnpCDfnUYRh7rf3kJKXp5We5+NohYSpsc7ilb0RXr7WgO9156H1fnA8OeZ2r
YHeilBoL7eHUu2d6hty6f9sf/Yj5UIxJPBncZl5pTEFxtZ2WD4CtikyFQgF5
CYqkl/eUfr+5hQM7uM6X3DGD5PAiHJ9bNeP30sGd/dBTpNu4qJfgAeS1DSd9
EXSfeVcJIF3KrKPiRNJOxteDIqpto1buFrziYjtXcuc2Asut/ZAnckj+JrRE
v1XXsAUKmGeJTo5Os3xxsetTzu/RyEKmDRSUQlMrkQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
L1bkm0E7lmP/lWPoRf2v6TuE6K9ofmJkHmLM7/5FnRRs/7HpG6qDRbERqIaj
xB/aB9Dbinn69SgFyZTKcwoBphvZSjn+elG9qVR1JEKBJO6ZiZRigKVCqbUC
z2xEZwqlKDLFJdWukpy+2YPq+d5pEdPalsHQlNsq+jbEAZB9Vrx3t48A526e
4vegxFINDo8lDL9SUoeRAYiMnvaLsnz54WEgO3B3f0vVYD1NIxlP1DxgVRjI
lt7T12vQKotioQR4tPPwFYeph6mM9Dl6hxrWTrpFxoqguTWWnTObjxC4dRPA
M8ctXeCSRQktQ0Hpfk5GPKHqe+GSM9ZDWWBrVTZaHg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
H+K0vD+H//WTwE9aa7B/OBz6qFC1v68zkfIBVk25cMbExsQTgZ+pcOowoao4
8i1yw5zYS5rvAXXUfT0U48jpHmym2sm982o8y6/hxRY+FaX/IQksAVrhGPUr
SFxt/KkhHH8kweV2u1mKOabIqweYRQwLCKPmfn9CSTS9SR4zkWwH/GpzlxPb
E78MbUsj2WIM17t2hOVpooDUk7PZcU7PVcqlSoTdjZKRyxu76zlqlrY7VNU5
Mg6OsgfTAOje/u3FTKwL5ZPLpaJQumG/nTnFMZhDb8D/eh4YVA1s5Xvja8CS
02OjFEQu+4ax+eM9B3sALl5HQ4eZFmYQashd2jMqCw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LBJldx7tFCXnv215tVwsft6ViXKXS5Tbk0uDABRKHUqygggpwaKj2+aJ3ku1
f4ssYgnZkZbYEubt/6kDAgX+zDJof6NfRXnVxXbryMUwQb5eNxCJb09x7Xa5
xF3eZUWzqjt5Cq7ahj6+xh0GWGQl9iYbEqQB3rXR6rbdbv0gvGLcmttmdw80
XdLOYIPI52f+u0AITQM67QIPr6uiCsiY0bypXBydgdOzpKTjbOPQW9afLGNk
8+VPKE10T4ZwmpYp5sFVUN+Bq2U8iRc/0E4zgm48XJrqwkolhJ8x8zj1bx0L
/dt2FXQbOTOl+T6sH8ObaHurIUZ3e5pqgIidc90JiA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Dncmev/FMjqN4DIn2rwYD1nCEXKCNVyhTWRrQ+HfnU/E1ZO3P+gUHvQtA4L4
lY6PIeBpx4gNpWPQRq1JCeEaKQR72Up93u1S0FQRMsHmfXlgctYYIE4zLUqV
aJdJoCSntOfbZvEh2gLYiCeUvdyRh+ANyTYlXX5nTga0++ZWs+U=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
TZBQ79AuYRu0NDa7C6+OilMBLTmBK7nNZfbA+aoIpmK/9G15j7C8O0Gqr1cL
RVTsbbmDOSMJBEWl8PEQJPmkiLrbukUrshB/QtWeWbV0+N+pqqxi210hBhvI
Ganu0TOV1gKFOEeHmvwuOK6y3zMSFacr/ilx9v8CclE+xiKV3O8nJ5GOE+cM
lK+IxA676ORLatxK17ROhTbIQ3bcZry0fS392PLvJspyvsgese0VQy9AqWxR
5ePZhYQ3RLgg8v9IDarOyMAglqmrDaak/hG/9RMtpmlF72SxBaDZ28doNPSL
ak+J4nkwvR/TLQgXb/K/cY9r0OYe7145jUVRPKVCS32QjoO1+QpstFbipNFU
phiVCTQema0aT5YB39mBG2MPOEV8DW14LGlN6CfMGztv84pleAwKD5rWXUIY
3q3FI+3ivISms2tpPmGZKlQ5CuWdVQLO6vBVlG5dmhBFKYF5hW5BN8WOjnmR
68dg7plySFRHcNIX2u5reraG6KlzBHzh


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qA1EpjeUYj/X5bJJEIgssdQv+8VtUDFsu1vdwSHK4rIC2LRDxVzBhifZK/uR
NC2LZMYl8dji928G3fcKEbwiYEUNnWmyuEWeafUihHhjne1MeSJbqXWpnXRu
aO+Ywnx33pJXlgr2yNpsa20ZqDd3M9+AixBgACgGNSDUzwoLFXc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XsjAZ8HZ8+RNm7lN174mnREn1LPWvv8isJrDWaSEU2a9Ei39+ytnRLf82bcK
yX7QfWBsyZaTaUTEB7KO8BwaO3DDXwKW+l5hzPHXTJbxrvgz0cAJmETPw561
4aN+bizeLLTrF5gdyd3ri/PMo9eFCh8enH4YAZgg1xQPdDz8sKo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2464)
`pragma protect data_block
cbwfgv08ceBVHFDEVHw68yfJZruc3NNRxCcmEUqdZe6NfCBVYenGgFfu/8Cr
MCNp1v3lpbRRmselBa0q+Wtov2TdMlvigcRpIa9OgYoUEEFH5OepR/RZ6wWb
YdP6Q+pkVkHbqJcKtegOUtmSe2Mw/RXNh2XsKEATe0GIdMYrkCCRy5dM1E32
mJW7L3O/yJ83xM3B489SkqEhEKcN/umGgFCq2nsLpglo8VX4Drl6cdO6pcKq
xgWl1uVFmkCfCNXM5rzSix7ovXDMTFQZtwOjItKQGfwW6k8dxeSIHEzSoeP2
YoE67q/WYGbsEBhxwEZdpGdXe9sJVDNQsVv3b/xDjAJ/3fbzhx/fOtdohzuo
boPUq2CNx3l6kDk1cAYqvdISU+R2EfpvMypxuYNfzx31wlKRZujmXixfiG1V
DCmJ4VatQrYi1kvNxCPNhfui+wedFJdhvvKMBCucpq+B3Xwip8q2NMKnSCgF
NERgEKEndlnS/psPfZoauSF7qD1hbMP7n8X4ANIszEhIwD+maIh2CEU4GyF5
xJJdoAag01hQTCqqomP8L1XdbQnd3ak3wTPisVoYpPaKifXNfIl2eBamm096
ksUdt3BKIkAZoKeUeGZgA0zQ8lgx3DRXhuaQ2oqsCW9UB7CyzAAJ5yTgyCMG
PC6O3dKhCxqHEYqkQZ3QXSuknGb/LebU9IX9YiWq0swbcTVZfAO0v+hJ3nWe
vZf1DcbXvShcK1gSOYdD+37aOnLfbEbZO8uRS3uLYxdsAsYpR5B9HtbYI36q
wPxR5XuldEy9hQZEMn7+qyDRN2h74gWUkRPdMPnvZHVARfikXNYzh/3G68xJ
3oFU77qIOQGHV+ZoUL0WBz5r0SCX92R6/wbzmnFNhVcaRD7bu5aStF/DNg7F
P/RLEoLhTIqqRmZY5xyMCKoxcvzBGWvogzG0OwLTtizyDXk+QBA9E8iXf4R8
C2I3lV+IuuB4W4F0FGDtDMr1p8eC5mznP6V/dtFlivcu1IHZikBe2efR/zTU
h+jBoi0ymOT4ZL6g30JQV9muugXMaLh8j72QTWQwztTIoe1FmXP30HY193hB
nQZwllFjWhnMejMyLSJ/fSzcLWnP99dn8Xs1LQUT1zLSGhS/LFAW4XnIecug
NyPNZXlZm905dqb//99f0Wnd4hkzLtQUDJ6KeVrKJXRRrbF3Aa9SVQHREjWN
gx9gps/S4we/H8Y039RtwTGu6KvrHbV4yZ6HIw/EAmQpwfNIrSxkTZZc+GLl
/U/F1H0zmkw/Hm2VrEs3FHUFOCSNSjmFYji+kFkcdBobJEs4MqewMPcT0fzM
4Htpd1azSEEdx/+UJIRmoaUBTUSBpyVz9fmnrdvv6dsN33H5nb1uzcE9cEcG
RnJlm+WMCnzMiErjIf40Sj1VX6AIv6VQeoftNZ+OUDgSHz2Nm12He/Aj8VOS
r7yF/hfe3sy1QU+J4mCFtKAVVhJT1UXlrpTZpNrjCX4zjwASKO1ZtaGwLlJ9
WoQB5ZjVVBPqvgOc96mQBmI/WFAzaZ3P9Dbd6ItVXH7wzSM92CWAxXApg2Mb
H0GHYJTHRzNOLFl/lhHAHx9aDlvgBhV9y0az5fRj4YdqMJilJYf2EWQ1hVb5
nGSd20Y1ZUUp+uZxC97uVWhCkyKyAYaEi+47jDxr7y9PnBKcWdFgvHnVl1ws
dFFWykFv5OVI7vVLWtPYXmO4+9JAsTooCJPslcIBnKsX+kRQI+MU4qyHxG9U
A5Xrg5yMOaLFQSma6VcuPrF4/owkktwjhbBpY74BCNEp8pQF+WftOFgrLKJz
LLdC+O65Im9skiYxAlHjGqsZc63FK1z4Sjk1BVwGxg636izI+txRexMujkO1
D5eXWuTb6OI4i4OENm4CKLPSjctNyEqtw3VhFkRD/5LHGaGCir72PvGjflRF
d/6pJo8kGaM0E5tW/9PFhLZOrQXzBbumxtYOAmi/nmIrDqBsSc/C6BKRwwtx
xuVl3fwAukOT8SI01iNuQfVz44iPmb8VawU22IsyaYUO9WP/d79Qc4KNkWkd
IvoLaEM1G6iaP6QRaxbuy+tKolMpz/RjARs/qDmscXKIyZpGKVYNoS1P9pNC
V80Dpl59eegJa60cWUS0viP37Dcsgx5wjPmzl2vWxXsX7T7s5gHC9BEmtINE
tHNTq9SIkQelxTLoIu1/AU/26/NKmO8o3JPvB90i6/Z7ejQclKlb7VE3QyQR
d+gmqt02GN5AVNwpGYNJpTYwY7szw8RPFEmAIak1uSo6DAeUvTIO8YAqGFob
GUrem6+q7mnOUdhZ09Ocpq4N+T2YpwPV7OoyieCK+MgnS5uYyuMuG8XHVNgj
JmkR5i4b/xfVvkucQ05GDtQq9YUQPmkcLp51SsZMaK2GnjcFhMxXYH3F5PRN
KVsX7ZQ4wvcMEYQh+qEovNd+o4q0vTJ4jr6IsAwmezCjQXIxXhiKWDVKyoV8
9WtduHIZ2IHstj5nB/46eoro5mkK7cF2HScY5OEM+FqawSbU7D32wQEL0RJW
ZIs0vMoiwLd0rLAewANX0l4ly8+j4BH3DdRC+HoaY8vYMmseBO/FTWy3TLqD
j7KTQ6TphZx3z+Ue1d5RIxgzi913MD+XpTaB/SK6K0Q4LRVgQo4NWlVmL8Ho
MckuR2y9tt1qD3y7nbuywMUxWj+NxLV49FCLywS+Bvtm8fZu7kwDPFlG5qhy
d0nXwwuY9X+VCd0AZCseZ/oRTi1PdmrKM7eaqZStrhIH/DvuLR/c+DALKeSR
qQRXu3IO+93jxK4yh6J8fCEgnSy4w1YeRCdEDIZFIvkv6PvClyKtuvFgy3Td
Sr2kEI23KW5sXdNrvhyQvyRB0KeYvj1yq68OdlhKk6xdpdxEMo4pLGSBnZu3
BJsN+t71R8M7O5HKFTsPXsOvNoIdBHZWCCcbVeSLxm59/9VzEzBci4/ww9lz
gptVBL7MGZyreiyGWZQdhBl/3pbVqFACnNBLBZOK6hymDnlSm6pnrBgAttp5
EoiRR6FAsxmer4bEmEjcQ1lNVr0qVXVYfjxR+Nt1q7F6Y/+uiMvSoNCz5eGH
0NfUHsmibc/MskmOXLv/zxWG8VWewRSUuzdar2eNmtRXCQq0cjLMAPLedNaM
/mAA94QuXg28g1m0Wt/iA3XfSa5sdIUKCTCTfqzUDNZjpdt5nI95WmX0Hd79
QjiCotZ7YlIpNVL8l5PHVmQe4kXJIHEFB2SSnK1Ee/7PfhoOhnNA4jucW96U
1J5xacTdNmohMzn9EnWdAq61Mn2HNsFN4bXcZrSnhIbuOw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "lK4MM9NDeLrdcSiRM+VIuNgpOLUAzWAt6nzBJ3Vw5tvBogzjtStM5gMJjD6PMmMyupOFzYouKIpJuOZh/11WnQBMmqEc6gvbtnHqfGmxFaxYyOv1rddc1B279ac1WEgUgi2BHG6DRj+tHk4+Vv2VvppW/Z9gUZ9e40aCxOYZZHwEVb/SJ8ximgD4Fihl81LOgt6U1JRoR0S/yAHMZXIkaoJ6FVEBkPAD3J3ew7MX9EwhFbdl70pvCwcwc5G4mfn0cwY56QDk9AVFBh2o7DxSDdOWh2VNnLSJQjZiPi/S4j6b9WjSHNmXGW/c/E5WpGm3vjve177Uvo+0OpYzhyDSAxfdHnKCC4x6EdOPmmbgzjw82JgQTPIaQHAzI3OltLxjJO8VrEmjagAOMOxm4Kz58cpP8GS/wCyW8XXiGMNh9Wja6g8bOi1/oWjAjgVXJ3bPGZ4hZ5e8vK6pwYeFqmxYBJEj4XEWkNJMxjoEj8ayKXwrSLByhstqzUSe8M4cwxrGn+WwdtVkQ6K98ySKGwjPM8LkUVdOjK5gYTf/MxM7wLoVTExI+tLABrPevWQVEFJ+eGUmHnEmI+v2hS9DFH42z2npLu6clEH/+b1IQQFcL6E2xrW78WvjpcC4AqHERkKWsBx3z42tnSm7mA3pzlvpc33xryB8AMGLDqWTHjxNdx0Yiy/ugnui62csCjrzWTK+jKPySlD4ofolaJTDlZ95a4MLxbL987gevX4UQapGNQkb929ABOF/djh3t2InhU5bWAvLzIlm2bMbqdeu1ZFFiVhJSec1O8Q3JQ6S7/wu0Sp6NENcRQQ6xs30CXOD4mPj/tde55deiSCZnOepSLz582aSZ4YnKSfmgAnqweEr9b1lw22jJAFqxvfwoFn2kJtUr+4R2ws+SYA7b1MSNnk5AKuHeBKKnG9vwkMef/zNQ7MONax5WtLG/yHARjxCCnCxL+OYhDkij/oLDMVoInlLijMpVCTTrT5nf43yUrPMd+qS5pcTTIw032+3Oz6VQ+xp"
`endif