// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TzbPxLVzQzYYADrxHpdMiOdL1/CwnQi8iKneOJWbsj+WP82UhBCctBAue7g4
VjreuJrlYV1yoBShGFO2Xh/RzJozBQwxzO5l3mAy+dN91AW8sKucmtPdHeDz
RVfiA5DI0FWtfBIExE4ByBu6GUdgyqbK5BIOy2TgqadO+aGRh3WrE5gQa2I9
Az3hGZtYJe0HBjMfv5VlSpO9TkaNbl4PiXym9glJ5UdKet26Q3YGkFipMtTr
BR0EkdX8GGwm7gcGBgUt8RJ9hyGMWEwxy6qUYF/AMVtLS1va2oAqHOjPvxq0
SdeXzT0uahrzONcBaq/JvF5DW83vSmJtu+68XHy2MA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fNPertCYbr1q1ltQHKjcUCb2IFCcu/7wGrZvp7kVsI40jo2lYTJh7W3KKKsc
CcmJ7nNC7C4ptuYM8Coj5dXELMuPVsdDQVWMzMUxbhcxoTBEWYHKdxbaw6bs
J6umyItkslqyqAEiM+76Q8ggp9JP8nuYoir85qL1E31fyqBa4JvEq0OsoDS1
AnAQ0HMTSxCBgtaxDYxA7gBuXdo0JDD6CFhKWjUAk4icli1vd10P6Ur/AoHt
o2u9eHqLNhAXm6cdD1icVYRZ6QtQlQgY8YG6NLDA0Q3ImXvhR3HtmP61ywYY
b/vxZ/CaNscQ2czYoOUd/mf5/qoF0HqkjF6drX08ug==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
g0BfaZ7EOQBk/5UhrvJZxgpRJcIXMjmzJzn+cBHFZFVDd1eN4lm0k4HF2JwJ
iP2XHt6DtvgQdaVR+v24hOqpGCdjNgOwTfhCXv/q7ZzbrLBk3DHOw+pYo8ob
tqqT1vk7f47D6Q04AsCJBGcVQjARSl9yf1elbe8BGw5JiBQzX16K4Baa8hZl
lHm/yUQIC0dEyjCEJeD/fgWf9tSYssTV3aNMYLcRkxv3gePVvwqKv/34rq09
9FIgEbEJf4m07Li38oMv00uhWadAStmND4bm3qXqohfuGuZw20MSyhjAQg3i
1GtnQlu6nsvfD9smSQZoIKbaJRAM9ik7okmC9Ba1HQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
b5iZAcKHwJQcxliG8jSug9shcFwLkrnqh3e4dfKbuITEXs5xBUnfIHkCf+GU
NTltbvoSLowaKfzXXU7711ojRfrzPYqIxprjEyPG5rcRPV9FMWhWQMJZy2bc
M03aRfWmmbQ8YT8fFPqcze0DI1fEky2IpZ08X7AO5kwewlKJvrWpZkx9Ql4O
K32dBfJNe+bQCNW2gBgyRWBCAOmB4KehTccMGLgNOvrRj9y3KzN1YJtLe435
BDig3DikcDUOAHqMna3FDegfrlXqlQXJvOdek+0Rrp7QSxHUSNWuAkiEL5up
jrwIM7T6yEHkELzuWt5dAOUcDZxBS6kbrjvASzzY5g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
L35oJTuIn4uMborvs48jAWFNY/E5/mRRG4TKvwIyXJm10fEXH4ta9YCeb7vr
2C3S+DXcxfiNSypRijTDqWvy2bypfrF25v1CVNLCAyksa6KdVIvkgN/IWVKd
D7mAhPKGoC+gjNtEkTdpmdn0ayxVWixdjN+oAZ+RJix1uE+kmn8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
xYHbOV2gxLJ1YeKlv787zYX//4dnJ+byKsLX0qna6x8lOq0N3GaB/TuayxnV
TSouo1Bd1eL8YuXlTSUPXkojV2MnNNclBMflM47CrCUy6FogScSX9sYBBcpv
+0vY1Nz0zSPjNtMZKRlLx9J1wyy2ZVdCwYPvfzimabb3Yb/w3Ka8tjhKx3wD
8RatmhumCtxZN649zUJeyMTUxqcdXD9GdQ/KFTn5Lgig4hSsO+dEome4t0+n
BoDB/zF6Bsg2Aca5+vThjZhrit6irvCwic25oFyjuvFi2hphu7oIaZW42auQ
FGETXH26EvwXzZz8vaAxtoBwa5ZmwZkAOYpXaDkgrajYMVv/iiWM0+rageYJ
AnqbhuUCtpnXSq4qU3MWacU+OyVMMfGCYyDRTZI+bVBE96iggMEIJQOAyJE9
eojgKrc8+GKTnzxpkVIFnqiFT7WUq7BS4mrjwgFegyzQqgsoDMlvyZCLCNLh
ojPlj+MyuzayE+wdN71h6ModQe/etMQb


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rikK4fNYV9irBA7BL/Z73W4cy8Ku37sVdrZlMafOW0VoJWunVv0D/zLtY0yf
eKnqF/wUnp3+mQ/+XxzPapDPZk2+PoTZuL0FqetL1e3NUThsRMiiYwI6mUOQ
cQ0+AFtl6BzpbmFxI377DWuUjpsLtC5pJPHSOmXFxSqV8OmNKVE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MOlq0ufE7/Nf1Qy3NwV58tPJvHoGCbw9dur2AcGJOCBaZGmH2fIvtEV1dTZM
Gbld6ec+A1feINj5l2USxXQxsWlPqEoVJ6hlFaDb5jXt85/uYu7rX42Zo3yv
0pulTV2cqp+RAXIMFeF/BtaKvUPDr/27arSYkJtl3vg7q1KgRWU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2112)
`pragma protect data_block
W7aOqja869QsLmJKRIoDNPuq7YY3ooSkaDyn7EQSXuRtZJdKiS/utE+Jq4A0
ubuQKk5v1RTAeMbhzC2l7tMHsA+gBL+IBNNdXl1KS7PwIjgp7uu1Vrg0exce
djArmlai5C+yEcH+k5ysl5EaOMLCVIF18thYfHdwv7dOE/W97KvS1NnDeoFc
CqlCJGiWMg8v5c2kNSMKx2704FGUXBo+V4gVA9YGrnNZv0ziqtXg4qU0Sw9Y
RwZcPYTmhb2T/kWfxjXHlMpYJ/4BLpMj733AHeJ+Vd+ZcjA6QueT1OZBlzoM
F+aql8CVSq5w2/CSsaBcXYLvK2q2vwYW266d+5nsYIHnDaGmd5sKTmR45q2J
7yXlgkvTutZTnwPB2TvMmaC9Eyijja9SP3aQr56Krt6+e11N8b2zUAH5IMnE
Up1Gjo3cbg1QiPfb2w48lEaquVK+GWk8omAPOiclID0J+DcIBUFZ+O70g/HD
5x4thdSgJJ+5NxsjUMyORFInj320OuvqZwyrJflQE7U1nQhLUNot79SKzHtJ
lC6ulOM4RgSiPQV+vpWGTd4Za4Vek5uK/HM9KE+iE2g2RGLYt8orWeXp/91k
HE5Hc5tx7JznmRIVdGawHCY1J/syOdDtdT64+WC5jrea5cm5SDi46FgpIsrU
T45OFyY/78jKd5c7gNVxdOyi0ShBmM3sU9S91nBcLoUN/J5U9NurJkBuA4PR
Y3JGTsS3zF1bEcoEdZJqGzKgQfMJliDytP25zrW8HghgQ6X5UsvtV53DiNRB
NIdR+7kCwu9TtQ0jAqeDzrfTRCtGDKvMiHdx6If8So6RnZXftAck/of0PoXw
DfFervICyZyGsMIfZKvIqfnzNy71/hNNn09PnvOqPO/jtWfbFmgh83A/I6lQ
27OmyBQTqixQT4DMU3q5uhZKyI5U+psRKHKof4jflcrrSfzFwoUyDOCfJg8t
CBiIcViSikgjnAhmJI2kQlqsKhEUAZaG/8Jo7IJBsV639x3yEhKaQXH6u3og
oQwfiHQuYfGP3rn25CRJvUX6XnZGbnwAKuhaZG+KCUCOiIRN4dAqODiaNHYt
SjfNGrpXz6ZGuhDKTL9R0gTTtcvlG/bcpIXgbsHWAxynlHtky2uDq8JyFpl+
P8DZQYEn6adlcB+fLxKf+Zhc3OLXJBdyektISjzH5NZtCXmYEB69Cq97V2DT
42tmgYEX8AmMpZ2fPYdgd9ABcIUKC9iFboja/fqTa/stC6rLujnyBQAl5vue
VP7m29/Edyun9Vv+sRByLkJFVGoJyInauFoAJ9BicDNr5WwlU6FQbWvTQhqf
Ke+fpxekf8nzAnLQBdZqUltrh+IXd6FJ+BZSaQSGM2Sk6TTJ1SGQGoIqoJ1W
kHeXTNlJ1us8Xin3ZRCmJ9rdFMfHNcmhGrByX0lLPZlL5PV+N3KDjhh36jJX
8PoLZ0L45lvZ8Gkri8YYVMXy4UE3LbD2+kKanQBh3ugBsfOK30VqBj/tPcjO
fxsTta+dXurH69Ps2RJ/r5ozYtEA2aFFZC5yjEhX/htBh0f1UWXQd+jndSya
h1pNvg/pZTEvzxX68w42PXmgoPu5Wu1ySVD2x961aIQD/+m8QL/yrI+9bdbV
IMpNWZEOcwebjzCl1dnwAed1cn9AbYedrHqsFvly9jcNxwWiPqMMV05a1T7w
YaOU/tADfcnwcULB5Yt1cw7EUqXwtVCga6lCBXacaAQBbrl2nROYJM7uX43d
O9cPix+LwDfKaDy+5VvUvAp0zhJtpGOKINr9IWbXxwJK1zRn+V32DORdOAS9
ivY6LG2VjEhthmL+TuMhm6PXVrpPUDmfWJULvS76TQwAQ8s7V9ZMOrKFKrI0
rpxGutlTjk2Aprk3TmccwM+xunn6z1WbNJFMDafm8u6UuqF7JTj0S93MANLF
eLEMAdCgMsfq//5aRdhsd60Yq85jjo13TBt3w2n7dthb6y7rUexy+1j+RTI5
/ZucG45YrA2Z9czQl+glHMTJ2CrzyMd3FfLN+QsfDwaWNElS00kuknw/862h
gN9vhdOPd1J0hwowR61zBciPi2gXs6Yuhj2F072dF2hpuf00UWuXxjjyMMbo
0s4jHe0v7UfouA5ek208v7UfSln1zxweDdGSHW3BRONjAGhdstSkxxt0yr44
82J4GjmK0/a1z2E2pKlnp97RMbxvWyQ/jCxrnnkITJnwaQAuaUnvpa2iIBkR
Et+g7A/SzUzjnl0c1VeZOxSJ9rPTfhU3SQgiZvcK2QgChHK2K75G3IJC8Hsl
oKcw/hxjk2KrgDYnM0bb4Bg7Kqk1gXLUKTa+CWSrKF2rAsRzJmGPK4IPrW2u
qOvfGZ5DZ1ROGODlMdmV/b1JWg/sHbeME+HPH6n0eCxl+rMXG6MbTHhDtoW2
E9ghWVJl1c5m9eTEfwCUbgbxgqKJ2LorCwstnKmRiUHvOMtmOpQAy/hLx36d
fDM7MKvbrOAeWUpkOY1qWuFE2H9DLPBSqNlUdP+BnR1LxQEI+l+WiUxVAAZC
7wbsYDznAHKbWbPmPb2kV6CSz2r7Nyc/E0mgKrEPdjVZYzbGzqbOCzHBpJ7T
E7HBb7GdqsQPSKKfMN5MRY7lDnGBWj8C7VTe6qDFvYrflLwydkfWR9rg64pC
KpeyNjnhUldCTorppJ9yVY4t8PfsKCgucz5qjC9KHwLzZhUqKPdLV/Z8P4Ww
xltmuCPfjGXZs7HCMvO7lQZ1rOvU2r39sDZC9OHIhCVEKVp5nu2kp6uDjQQu
/3CUBRoWUsfBaymTP7HNl5p1EHaARm6R2ORwku+Lfu1rZ5oEp5sSgjKk

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1JAtVEO/2Y0IFFNfLdnPv2W/qjul8yY9dC5OyDzPQdSJSzZXxh3eCM0q/R1JeQURcafOTYaIsqdrkYHXW3s20uvm1yZm1hOv69RXMbWeOP3BRO/w1wxm7rFqwgUQON5wkXE11Vr0tJJ5glOpFoRhC33NWFfVL076ZyGKq00xTgxPH52cW5Yvo5z5qmftZciGiPRHm+ifuEwVpAdblr9l3KrIam8p18PKFhCDDLU0RAn9I/V0ng7+3y7jQu3nLzDJ3qDovpoqjsvDfLJ2W2b5A7G5s23XdmbmF9wSgvhq1q7UBsXe7w8W/MgsdPGNRPaoHL6HtrINHibrSpBR2XczddcSiPsKUAhV3Sdf3gWEitTlDIz9O0KADPQU66r917xx7wYMBfX9YSFHl+BXnqo2zyodkMZ06byFh/0adkYQ+UpnfgGZtaEZnGL+YIw8ageUE0KxK4AW1SVmuwAQpQPmd5PdTRrVtF0eagZypzgp4O81Yuthyncy8/aMoZAlpfyxrhmpuprGyoZ0gF2mp+Xmfty1NvBIShBtolI/6SyRH6eosQ0zKG0u/FjSWOLLUhmAFRvofnZ7bVb0C5LVCZtLb2DDzMH3aRCyRqRGN/icn5ACyyYB7nXR9A9Qj4lQW9uxa5Pdrpf6thAiO+XGwmdFE+QyS41AuR7NPBddH9LDuYwiWypZP3CydMJDqJ/W+epJuJRpkWiYxg/PjrI3YQZuMR/ZynbrazbDFLpGDQmGuXN46U9/Uv+whGAgdRiiLLl07n7tOZ5m3BvA5YG43pUUcLh"
`endif