// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FSw+mVbh1uVFG0CRK6Q5XDr4jttu3MGUeEO9Rq2YnyhZnrUXq1G2nXGPWeZT
2R40erOu4kC23PzpC+tbLVO4rKUS+9jBUkX407dSuw2DmR2u2xJzLvWNcEdS
L18vI+SKkKF2yd1iz9OGNicr8Oy/gZdVSvf3Npfl2eRZtZ6KqGT/DDW/OBIT
bJF5LDX9Iyf4z1IlhPdF4BXkME5OK3IdVF5RNVx/TDLFpDnrWVWP1hOl2NSw
fr+AVMMZ/uV1gWrTkLYvr+rD5oBCN+6LM9InAGk7xH1jlvQ/2a6J5O5jrWKi
iNb6MDh55dqIj1wTovykGp4hS/qkbDt4u6dUNRk02g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gT7lSsq5iSEONNE/0PUDSTKgd7R8mjCSG3YqC/LN2OQxEUd6ov7wV2JLZLCh
kQPKHfsT+wGiKY41yLSI+aWrzjHLnJyEz5EEE+for2FuFfuk8dEtFKiwGyGJ
P3urKy/ArZRgVJXMhgk9sthDhDPZuwDTp07sT5LotKV/tEsz3uuaMQNnOqHu
HmyQi4RjacCpqNyk2JPrwXZ4CeBlehgYeGxgdejcCxUjP5gF3yUQXUtCcbQ+
5OgX4Itbyi7/nPLM9hdtaZ9gdyyy1UhUZ2bUkvbjcl+qDuopk1o75sCQo4yo
wBoF++EMFdFoYhyNqeCLLL7FSaUVuj8VjrdSVH+KWA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZWDE4/HQL0f5W0Q+fZVzEClMg4UQtWty6o0UJZXT1xJs5MkFCd3HYkuPcyZX
FoHRNgNH7faz94cEE1LwfhjKAjlDiSrH16QIRRJ/IIDkgIvtMYSyv5Mvb5DG
oIMgHYd7/OjLoBY+cMP3ahQkGtWHLfJfdeuxfSc4Xe+OT2OG+OdwcNUHsOHe
FVdurr/VNbbH7CDj2nuZh/aUZaQGIJjOfliMvVcRuXupgB9w/8wrj3CGMSfJ
W3dPqEhrGMFogf4Dx0L5KICjX2K6uE1XKQvePX44mBuV0Z1Ts6/GsdPDXA53
cepBdVafxSl8syqE1INgkFzRcwlrUOjXW+y7MTxhMQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NFbSCBHNYSqkJPSLFR4ALkw2Gl+f7XV090pYvBptIXyaDK0gSzvbxd8AqqNr
iKTkYMyKmjBWFA4xqZtX08Dsp1fiCZbBZfI50orpsva40Xfpq4ugjXoupNy1
eTT7UIB7MxkNdPNJCI3zm8znD6wbxm/I+TsRjhfIo4pVTbVnEqmg3VbYfXwx
oioh603QtlWmsG+3VbJllKp70JdJ2ESPRFsrcCOH42zyJVFmLTds/AEt0Hyj
Hf8Ya7gdutfvatlGBSHG6mfnAFJW+KhVZn+rjSjXdYIC33clFWvyob8dEZzj
oCK45r+pTp8nnzwr4todxLuL9TyzIsP/3/q3yRfvtw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cpcmDgEZeNSGp0lZK67afDWYiHrGD5w/TSvO8fw98VfxPEX9rVPTu7tc/byf
CU7uc5PDglo5ibjL7b1zl5kcLq/i3da8xJK4ripYf/1UsotGotjqjq5O5Vw/
gmBzUohxPNKypzOY+QVdNfzVtjOEaqIzoJpfh66VGhQOiOyP6fk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
yOEIvm4ueb0OpxTBhcZhwzHTD2vdTi7WL8T9ELkT4nKTvuWjL/W19x/u3Qxf
Y3zudLx8LtymCVJ1sAIyg48O8StMZdqYJWGnd9VrbVt8rbiz3kqQwabmD4CY
oADw6CES0JV+OcnCQUwdwunCnSTTd0dJMI7kkil86vL6rovnSaLuIXV5721N
Wt2gdu7QCTdZBs/ryYK+cqX65OkGfzhaztCctGDlM03NtnjXfQnt8ZVunspY
yLfU2k2eM0QD4EI6SK1IPpE8iu0vcyw8vME6Ca77a2wuUD9UDdmPhWdoXNq+
KQFXNnZLTaqb9v0cWGPUqpKyysdYTQzZvsILMC25LK+zW3/SXC2YP/FV9n/g
S/KTbm1gr0LQGY+7Pb1BM//3HvdedyR9wU+ajjbj0O/K6EtyZK6cjA6hHCqx
JgMnQCm2wA/Yyw0NEADgEV8SPU7sjgmN/HkYwvlE8uKLNmRSbTblNI7E0KnG
kdyKdSpuzGilQxVp8i0dlrDvNfE3/gjt


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nAvqHYeenzTRdfb8POhlPjyP9k6AwQFKcqqw6YStL+wfDTjsKYJG2doLzXz/
mrlPSGBvR74FaCcG53g3u4pfm5yid4ePyu3VxtHIGd0gyt6Wi/cQDozDF2nX
oqyEgyAHa80QNZufF/GNfsKLgrCu2Ww/dCHOOk6hqKcxaWKBb78=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
G6LZMMPZ3gVak32Sbezw74NUYo0a4fFIweGZqpfE2PMoyrZxzhuaXURwfaT1
p+WfPbw9jM5ZWAECspSXXx9971A4J56mfDS0nTY93cQ89YSTti5HweabHWJD
9kRGIIhoMXQ5A2aPqzXwn13dQf02jWJhUVgoN3w0MHQV7fpB6PQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 11280)
`pragma protect data_block
VVdTf3PxEBqg4q3JmbchpWCKv74yFWrzRDlVOWFQok/mel1HW0YfNszD88kJ
YyuCtsZ+2EEQmNJ/CXw6Vej4P7V6IByK3Lkj2qYQ1j7ZczoY71t0MsrcBwcq
Q4qDJ3q6NM1X2v7MsIAhBH4Hcmdi9OyJ2UfCRR0uZ3Tds6CCftlbgKWlfbXu
XLVaX+yTYrEQc4qGEI6UPCmJsskPnYHk0OXCn4YfVkhrJdJcS7coyXZ+dtpp
NuLJD3fxP8wEs5nZdzFW0biTCE0gkEgUOz0W+7m2HFKE+RFMcsGnXieJkffY
8HdsbwHBKvldB8PXrE7jSfhspYCiGd0RPnkRh90/Aq0tJP7egyjmx5KER8tk
sJyOcA8Dztie9J/S9wLL0A5ZAB4PwhAL34uSqAfJSf8rv+tVts16EszKjmaj
MD2YzyI4YMwIJUdOg6GnwHzxcuhd/XdTdMzrHnYIa+16qvvYkw8T/5QAi7w9
zghfXjeZaAaawa3g+Tbbq0DhUeufaxIcwtIFxQbOdJctip6W+WMTuKdIrAZj
S/bi1lVTmPQTCdOpHjO85d76a6WByceaBamMnMRaRF9aUw8XKgdDtIaGAiMv
Y27KZRqR42QVord+kIKpJS5uXafK65+eP1tox2IfnJkd0M1DhPXMcHrGqf5m
/yRHsmRNd5sKOidn+/6CWydjtcQyiFmqgaLpdKJTaCVejMPrR5fmGWy3rTc8
tc5Z6VgnEBcSjjbb3QJg2+Bk+YPiaCHT1BvPJvWCX0XkB8rxLuk+GwlpcyiU
QvIdnckJnlV6xbjMZfyR5PHMWnEu9tgX71alQDLqflu32s37p5JwyvVIp4z2
NtuUg8FAn8TiyyXOkaeS2kSZVdaMcshgiI8wPzA2NBF6LsJcBmVMlBaFpphW
UCBK5M78S+j/WQ98p8Duq7deTzwt5CWj0HZy1bWQyq2tYng4nlzHlyRtP9th
oXEJSvUeumShiciXSvyc8e5PDkRVpy9H50Fbu87fOAxv2ICAlmi/vQC3lcLa
RzxZRvieFVrPHk+TyT/V9nan1NXxSOwV4mZvVFw6vLJNl1+Pyrts8jyB1KIo
R05z/HxD3LsszPR2C/Y3Fdm5Kghis/1Eb3y1FH+wMgnLHTJe0u9bZxGWnPEG
Znf2BrNS2J8Tef0arSvvfUVaEm6U6yJBeMh8HY8UZ4oGhqJfHVj3uczzsBYb
LEGfHiVpRzGTDFX+oifnL7ZB2exd/nVXi9exu1TaUbRp1Ur95Z3J638kk10r
Ptj2effHzw1cLQKq0nwGh8zetLiqoqswWdavAgpIrvVPiZprAheaav6pkcu2
w0cscR/N++q3tQ0kPZdVGcb8SPS+2mvpClRUx+38fLEtLiT0GGVu/Lmpg05e
sArg9qiDCN7/AKaiIKE0dLhoUWoyI8Sj3JWlu7q7MQoPGxVRWeQcwqcMAC8m
LffF1RuW74XHeALiAZvXGFxfRIo39mGh67HewwQHSXylxpxzzY8DIu+/NIXg
9pYv1UQg/BF+9yjmzVIoGny3K2dAuki9Ix9cHn71MP3vWkDx5/aC2spj1+Or
ZYmabPPagLxFLYVoqrtgmGZRmy77EZVorUdFxBseJTUWnY/Qnr9kRutylvz+
NAYnq6jJFD4pOaYMLM+s9+BFpkbbDaa5EoMy41rHploxvTKMxYOtZ1qBLWlg
dDG+MoejOcm0lt30zXbltvnAOSgj8jmV6BBBH8qOb9+tgkH6Xsw3NYY7/T2/
2bCLIfDGDm2UN3RoGlF7dDJpZzDFC5AhtE0bSoZALsvpVClEmMAZGJfYMQ8d
8I7WiNSNiGMPanUDjSc/haAepo/fzlfdIWEG8uYLuMYPB7ZF0aSfxdyJXCXt
nllX7r4EsTQbwz0RK+3VNMHeNrKnNy+FLzeyxzFG5J7ilpEAid6FjvUpc/6a
iSh5FstsWMtr0dz9dg6Zr/6qFMgCbCrBkPsPPwUkoyEjPMvfGneGpM/C2BKP
cYktmrOTjqyp1qCA0LKhk9bHd7DXzHQ910omAdvNK/Rz5xFEpnvvFrPUYFdA
pDiti4VBUSbDlyyItEg2O+2c+qAE/I+EaVsHBkEiWi0c+ks98b4iVFyCq2Oc
8dI11Ol2dFZ8mg0aMa5WmSw6v36vvMhgV7kui9LTA7OsgMrveRPOvn+yH7BI
GaA3/uuJ3U1wn0llkb3tQTL98RJ2HHFpeJfaMfYeep2rbXshdKxev6Rpy4jm
Bbu3Kktm7Vfmd7OngRBiZ6cu4FoCxDShbf0+eX4ltdSwmreE0DfHWq4yDtH1
pJpL33HhjJb+5/hab6WtoHvhLeNMb/5iIMf4WgVUTVq+g/F5ilRdxE0JYbR7
namruAUMw+vfJLte58eiaZ9JJmILPyItUdxqo2NaU5z+sVlB8Dytxgopbbo7
PwxC4hPc0cM2iRTgZ1a+rV4oVotNOeh9AXusp5+RwqC0b1LhprBPF5xSUuAn
13etWE3ZB1y2z1iD6D37R7Fk+CTWpa/UgPhCTMoBYVyuoIee75UROzMvSU2/
gZh15ubbgxDN8NxZMeDU653KcZz73189a3bHH2YGG2aonyjxjzhkCi2UDkX8
Q9qPxNFXKG1aqS4PKJvcRc/Jjq29Bmy/USqY/x/YTkyW5B//I3cBq78Kj0M3
B2by4l6IyU55/Fac0DumO9v7dRMzODHe9fUdBJ5ip+4XaMBotVM6WZGZnTmx
ttgDHICQ0LJUx+/U5Ff/EnNFfcYjsSr6DrY59gdlz7DKUq66V6moSFt9lgFs
U9YdyxHvqheT27WBxtp+9RQB0NooQECP6dp4Zq453t7oPNtSlXnG/ZtHUOOU
ek6R4m2//KAE/8nYX5gwl49PvvVHaTA7ngI2un6Z9lJsdUr8CcgFJ0WOSfP/
40jeqr+jCNvtTYhK74cgcL1IXqih/P2qJcf10RrNJXzZ/f1U8mtrBEkv84cs
jz1llYUhQVf48tml/w/tEfezwCQClt7GyGKtmFlFG/WCmVcQbCTdJXmJo3t+
8q+MDjV8ILZQekeab4lVgGahdC1qbpsGtK7t6REsnm8LNZaZY8uqgEJXkQgv
iioF6Ohp+J7mF2Yy+PmqUJRcfwdvlqvFob0JHAKPFuOuTXG5aFEA95UxX7qc
8zKu9oLa2bOoKNwDVeUtaKrotffS+jh6XKauFLy2dJWzKUO18m7UW7N0JSbF
gtVqTj4YWw1GvudH0hurA83mUfX7rKi2nCvAt33sSopK/NiQg77itXG4Ch/1
yYXs5k5rWK0D+9AaVC3Yc4EQh3MS58rlH9wR4UvpVC+zYyd9XALj5ZlSla1s
PHLt9UtGhOXDNEY8bU/9MmJ180F1ZObkHIMExLGsipCKQPKwarPNWBveAI40
PotQjk40z6d2YxKcyY3ggzEZQcLWiNMFIKIht5m+JF0xaN7JkyeegHyY08q4
fWvdwMdae5PS8tVWzk9zODQ2mTVsEGeHBdjKxYYQeQgbyA/MpVuzCMVEsSjB
XVw3qaSIZQ6Vf6l2q5kZfox2D+zOfkELRF0a9rVvEu2xIs2aJ5gwLkGCHliW
OOecHSa5/ffeeJinWuonRQayQTHncLPr+NvyFPfnRdeSX4YdjCU5gcAe4DxR
vZ7K4hPKUrMm5Zmqfgqko4Rxz6QWgC8gPB/4k3otiA3hlX9OsRAi6GHy1OoM
U/7046tthZIlMoBaN52jq9HQWqOTZ/XHRXGAsglbxm2FWFcOB9R5ZhukzJqO
QY2q8rhgyzMq5uRQ2vI+sFLAZyVpcLLCFteceiSpYziibbhLc2aPSyxhnxvF
o6ygeLk1vQHF2M8MlRJX0uxPqoa8whqSz+3dhaVh7vLxw1IuiWhAT8hz2zsr
pHNDLlo7+mMK/mcOv9mzVmOeWLnOFfzvMDdlDXynUYssLWuV/A/oR3Fg9H/T
NEkFkG1f0ZYlx2e9FUW+BmuDc5/prTwfl0zgCKMt+DcKLMs+5ocJ58sQqodq
D+CZrF3tO+IZC/e/dFVnslQO6HJxELbtAwEW010bp6IwcX+g+iV0suzheozu
JoVDKkwyiuwjZP3hMsht3rMOWZfwdAgOhVLPyV8Rx+9fK0eaGEf02K+tHzE6
i+grdQGtzCy0cuQO0LnKoqhYlDS6imdmreNRlSvU2dqLsuWFGQonDJYMPQk1
FyUddxqOWbc5+/dorYHjAnqmxNgk1Bj4gj6cqPRIwuk0gKKtprVxV8olvrJj
uGKQz9IAU+QtRM1VqaijilkDFPBW9hGL5pImZc2MWTFSA/2V0T2pGs+eQhMP
uXfyHXdWg0U3bvFZrhR+xUOTQ8dy0Bor8goAUe9Yw/YmdyEf3G1CxG3rY1KI
R0OSCWPa8Zfg5iMouXFzOwgNFFS+Mz4rOj2xgpbgtCwJhWrAAjP13/mLyMYI
H3lPjnk6/5gLOz75EZvDa4akaYiMn2g8sKkKJdXaKkYfjWuolrr45oOJmq+L
Zi8PXlj/ZoLBKtXZBj14+QqlTDFwL/GH8JCWM5jXpcVXENZnUK55ryWnuiiS
OtGpEUy/FU9SSHUqUl8UCUXereaPb2nkX/hJot686o40w0mi2sTLuXvjj+UF
gJaHfj6Jhzn44rbMObjCCiR9ACWyFMAmZkEicFP+CyXNHml2k4N0BehEzLwz
ihqT1UDY/6dPrXEMXjcV11aTwGeaAojVflymBEJD3ANAsvJqhYp8y0Y6gWOg
cyigm9x0bvlETBZHJSW5TiLIr8zG63yyaWg5eorNHKEAd77SURB4VQ483sM6
6tUPvLkdzcxY8psW5dzKZglP8N427fr0xdKuggYBwRk6mMRYjkDaqqhlqYap
jJ0T2q/xVx+23BTtxzhPHa7QneIDhK+UnQOY6H2numN/393ger6JflzE41wW
jIuYMrBvRZJtYlBEJ7sexixIDVkhH73nDS90el8JFHZdf39yLrt+e6tvldOO
5rdkCmr+A/hS9kLN6vGECCHD8dDg7RJ4dfTcJbwsTkvNXiAsvaAq9ZRoDql5
XLqoMmr0x4JsK36NtGhQUyirYdePYom2L0BE3g4Hi/D+n63ciYNRMGLSc0gd
59nm66Cv4IlR+iqbEwlpXM8gobJODfaOFbToAG7k2xQlgJI50fWcMIbkKjSs
zVwrNN8XpLQF8689NHYgxgnOG6TeFagS2Mv9V8szayrUfnfDh7RvaeNK1A/X
qoMsYfwWyglUfZWcXkCKsdx/F2jTHPwatRceID5MLE/3QLBvAb1p184ql4ls
RibSwTPAt+XeCo78QWIpoOukBPeUC3Zk790tBKZlTZuDRBVc2LhTqcaaxSwG
CEpDmwNBSZwlzCuNqRhj4Y5B0tBvENSbMzipjOQzaIQll81eh+j1IkTs5tie
Z3Ladt7E5zDR0t+aEGrXPEo3d9gEPkTBtZeGCJdEWXxSKVG8Q0KNtASQQNtk
37soQLfRVGj3MKSow2GQJiOmDq2jASDHyf69t0tUHGfVwDxamuTqTa/Qj8T+
oTjfOfwZz9VUX8wSnViY7abX2zzGfz0SKVLDzOk2C8DfQZmtyQR0m66Pw9AH
x3xwxePey/lLU97SM3GvQlPIoS01Ioq5NwbJCmxAtIh+QzBkY19ncRFGzI4U
NtqTpIwI5IFsRK+/aJ/vv06XJjRB067/JmT7ezEESQGgpZBfKugAC2G70LXv
FJNJdzMJeWJAWJbhCmSy44lTXFVE4p4SGfcMnmN5mj+sWYMJQZMK1AQ3HZ0i
Fu3i3ttEbf5JXi6ZtgKokIPXQ5CF8+IoOFIOw5MvSn4ZdceQF/693FN2fI8c
eHsmRj4snnnrkHs2PkUdXZqEak1T1nWhNYu616gADYtGMlgPyrcjcX6R7YwS
UBEvTGj3TMnM4C1bnNEo6Dn1Kjr6JfsESmCI6/mjOzhW8slLkktnwfmeelA3
pggYWVoN/Snk821n7BrzW4YpFv5FC81hb+FXpHX/KPD+Ukzb/i8uxKok6J+0
PSJ40dt5dq9TYfxT7nVOXQ6o+s4mOm4iO/fBs0eZhr5IGOCjSQ24SpNv4Gme
pCsXIaDl75ed9bKar901S4fIximqPhYR6/gsd+zU45s85kR6jKscp7jtuzYv
/ym0BIyYYvCXMItRYp88FYwZ61S8S5+WZw12u+x2jUnxV9Qx6xoGJGscgqQx
6Yogxpa30jt8PsBTGY0gbEYvYX8qpERBNrNemFe6D32qPwloi/xiUVkWsg8A
BFMAwLjSHKV7bNqdEoLF2+6vhiuK0JHxnlJomZgKTFZsj+zInD1VZXNU+q1k
BX9D1/z4ngZRD6kMH/hOc7ugw94QGw2qe4ymq/CLCmVKNPeHyBD+NSTYUuSA
A0QHg/p+tVToXhQz6yltDZp5NjdMaC7pc+KvMb219izbqXzKLdRMpXoK3r75
cfJ4DuozEfr3J0+pXollOp/db/kzoSo+XT5Az31M6rvTdZZpJc8wxyXt31pO
IXkvoYPfWsN1kC+jYiDuAIn02e4TM2/p7s/Fw8oo+inkw2fRSs7hxLn5x/DS
jzGK1RLroeWCmELYvGyitJInA8ewcdwA4UM1ivxhMncjQhFlIaJAK9d0VZlL
cH9cynPKAwYmK1QLCr56pN4kq6QCw1s2/DDKrwww5hhMo8ueng69ZjStuCAM
i90u5AE+e2rLXi3TMlbZxt9h6J/zFfPudwhFNpSFdf9TcX7m/z4gYceCDW+U
6EohLhEg//yVdj9llQ1ukJSMDQHSxvNdCNxtQUuvmp1hKRNx7JhTm6qPw62m
ITGett1tjcvK9wiLC3Eth/51ZvKsg0tDXzXzYnCq7Ej48AgSoSBv/SpY9wOa
fWq7rzRup+l/IAaVqKgV4VNKW6Mf+bAbvv84KJUHWzQ3yayWrtX9n8TTOpGY
AcGozsnF7Mdn0uehPvGsy5q7PrhyHYUKy7tThgYHHlADRxPK2UZaUKWUEwkJ
22Sfo6H5IDdFUOgPvEi0fMfnMudPcqo96CMXuErF45+XVXoe+jmquT8GwdIh
kgzTEY931D2bhLiVQHrRtJdPpKYgnyclkVyX56Gcixb4uz+v4o9voQpu14Ks
F4FcZIQlX2ncNDA4t5mbVRUrxaEMNFcyZAs7TI2Izc+8Cwgmx5n3U1RlkcQJ
r88hMg3EyQvmWepGXlZ09UG+uYbQ+oWJm0z03QbvPu+O8INznYT41BAduRNL
VdpyW/UJGc2bg7g5pzy9syXlwbd1PvrvUMN1LQkc3e8rLplfVmR2dunLOwO8
fSPk1KiaCQzie79wQY7nXB3xV5+ngNwGFSkOZBys8XQFt3Nd2fuvbM/3yaKf
9iPfHzipRSFfy2GoV6V/CzRP3syp9gXGWveU31XcI/0gTkRZ0mayLEC2BXk/
Jkw5yMluo9MVbJ7y/piXUIH90SdFctYeHKdi4viOtIX1WXa6c4GSFpNyQE1J
1p2L6RHAiKhIu8hLHbpKOJ1YMN2MLPhcsGTrnJ5/PDdS3M+qrcYS039r4Onf
CJQEzOGNn7gpLeo+pD4KhjfYg8zF7c6U3KrTBXg2eQHbtjBMb3HukKXxxnhj
F9p+dI/c99HjLkDwMVHoEQRVBx1ukHHLod1UVK3V2CTLoSbCXc7I9QeJ7uNO
h04L3l3JAy/LB+BtcyQHccqhoXvp7SPeRH9a7PHz7Rf/mIgQGVBfQUFA9Cnc
g2BdgHC3n8l9XOk/hQqBe88Pps95ufPZZiyRZV6n5dyFS/8BOAGpRNjn7F5n
zJ/4NbWZaRSxzut62SxYsAGVgmL+O3yuSK0WQ0mQRxuvpSX/NKdC1N9MsdbC
bExEoXFbdgoztdLZn0PYbNMFsy27WQUrGk1hjTamDIO4dL49EcoxFXS+lO+/
dPZ+XB9Khqf5M4OfaM5eN7KzTJg7H4vdudDtjQ3iXQDeAsJlm7ePtzozpLmR
knb4AMfZfMlqYTVEil446Y0WNpCYwE3XDs0r3C3edQ3NYcs6vYAdCehZ8RSf
qREaQ3JLVrOWBkLPaAD5cKz/9T0vjU2oh5lRSNkQuqQKwLL7kVAWQOFlEmr0
AS2X6ruYu4RlEkJX6ws8gHM3arbsBp+NZGQ0uMyOd6ACmhizfbmejCSUtdf9
q/hI/MftqAK61du7CZed4KXj8GLBjmFnZ1EmsJ8kI0Z5wg4oHM8gZnksamqn
a6346+pIQW3dMYuwgdvv6Rp4ZxdmHm0BiWEY4EP36NWJUUjpqx3HKYefyjR8
L8ub1Z07/YPwUCF+aNyR9x9FRXDqB+od4pgNc5IHEM0PbESL8xFKMr40x06z
d1gkEg54VRtjOzdG+XwP0ctzXRBJbiIzCk3B1+efWdCNHqRWHhes0OQtyGMA
P+IG8DSEoahv3dqIVyu6EGLe9Wy9bzwdF9N3R1M5wowp3qrUu3sjA6tLPg7x
gk6hFI4ihJpYoOzSlqRnl6TZriziuh2XhRtHGBWS8A4ym1gIK8pIEoAZf+d/
P5hiq23Ir50zlsboblTUTSLtB4mllY8k4fDBxu6OOkO6ZCjxxGXtu5wUdkEJ
qo8jcdHalTIRZelHBTKcHk+u0AyfdjTcnZlk+dwGWigN6V8/aDTdWyuvaniw
vYBfLuR8xV+LHrgOAorD9NhG7WPcghKEHv41C8d/McZNoEhVQ/elY459FnaD
5XPIamcvGQ6Vij4aN71u+qv5/2hnpuZCrq7jJzKLL2T+5CogMzA0R+L90I3n
UtW/Sa0+JTvRHQPAPUvdecoIHX69AT7BgVEVDyUhFo+b+3LWiRrz79/RREwT
aWkbfXtNjnD0V8SgdlAzwqynzIZDgyaPfHVHDZTvYTrIg1BupyW3hZHT72pv
nFbcIT9T2AoFh8XctjB/BcDFlIez+o27q2Whrk+uUXiEissa7kMOjblNbWGl
XLggeButMd/lSbYdGuiW7fjLIfLTgwxL+IB/SWFsJzVdXVBovk343r2XQDlC
ddRd/DDDN+1/X3VOaD1zLsYC6g5yfOI9q+gzR118G5C49Ec0ozlQcp/R0fRJ
ZJkjc5FRWipo5Y3fCKdtsd9CbTVvwlirnTFzF9sdNm1dqsoszv81I4mwBX8c
ymH4cEbw4YZeXgUj+dBhe9AD18GTJAFHDCrY86Q30AdjEnd/gMwmOBV+6u5K
uLAy6ykDNO4IXJ1QFhWZvzt4lUsjQxLXd0DnhIbVSS4KtkD1cjnlzVNpzGz/
yKd05JIUXBjIw+BUY2nNQqoHSX1crZybVYfzl5hW4Zl8ACUrR2ZRlBgVz18T
yaVsWWa1fxhwTLeqQi8kBHHpO0liXzPCQwczQvXAeq/x7HvJ31qHfu4jhe6/
O/1XqmtOp9jR2SmMJbO+1WieYqRxenv2lQ62j1ROsXV7rXFnDOqJPBq5h1We
m32y7AzIl1EJ/b+/so8nYgNtvXjih729cjmKUOtcBr89vlGBF6w4gIqsSLMU
jvw60Y2DiziWmuBJ8Eu1/z3E4Cjmu4hlei26WvxbaT8Nairc7nwI7EZ/ibFX
QKMKUbOf/5h1n+lxdD18Co4XQyliiK6xc0TNR+jrUgpQd1Jpe2KWFQuMF0oI
8ABG7DxZNW7PDOQ8pnGMjxQ8kAl+OWKcpzo+WAiGnQm18phHKe+15nmv4E9m
GqKWTMGoExE8LJNXbrL0LojthyF+udBnhP11bgaPkID4v8TFLVXUbgEvqrAJ
DE80IZABLxhtHpRzj6tg6vSPFQI+jSyIwk9JHbgoX6Ax9wyiz406j4OQEC8p
MTd4hOALKPwGrkNEacJJGrpU1ATrifg/m57R6EHW0DI2Do6NQJp1FjFPT8Wr
P2LF8MiscOPROI9a1Jw4CuEUbQ8V8g/xVdjLKxVOINVsBONEBbAP2y4qAeVe
ZHqpO0d6yvLVva9ezvzclxmg3U0rkuknHya+V3nqHrq2TP05pPxcBK0jbFj/
ktUw+d+XL/wODdc2oXSM5elDOmCVNzcmmbsdZ1v6lRWjPstCm61dv32UKWfD
fUfS2G61x/1oYLIdeW97rQSUznlDIiDn/mQHA/tMTOcV8vDzw1nuAv36Lqsk
z2SMpsYQkInoXvW47KAUFvydKx4W12EGpEJw+zhZGS6XNxvNjKW3hjaMaMHq
r2f8zdzVXyUBvIyP8LR1x6Czmac60/Dw7nXS1bp0P9IIXMaMdAJw03Y0oHsa
s+kZRVnZhYHDWu6oi84Man1IBXNp4uE0rog4cb8NT8/GHcjCi0110Lbwe+zl
gT833yDmrqw4IcE4UmVKT/pECAi9mc7+DdTciXG/9oto5U3x5NMSKMixzHWb
W8S8NjFg0+DFpA+5COPA81Lc2E+kPz8Y6twgknTu2sHW6T38KjLsdSlYTPXd
MBhddJfoSwl2Vsx9aKCxv8G5w9SaTzEr9qSrPUZXk9dNVKIWSR1KHa940bdz
C6juCaRoexsFY78fkNTfDCcpOO4hcHEM+vsobBaKODZNmlYquLJFsT5z6w0T
psyHfRGAjai1yIF5ZxZbYhAhPALXsS4ZVuY90W2wPKWtlyk84J9tbC1yY9ql
aZAMV6VJlV8Q4GedjXGgt5IR6X7VAxggl1DYorVDCuNtnaJjNT8eJPxnrQ3S
rs4BCQY/FgBpklb7uf6TQ1+sLvGD7ZHaTC8TYBPeRSxThIC57sVZHfBsDhPD
ojRc7icXCD+7M5pqn+Go5RAciYnIa870XsiHoaSfkdDvqH00UmWHXE5q+EGQ
HyUH75wQI9yFdaXnE60KZfvDVC4H25ToimHuCsN7echNRnruJlgadewUhtfN
osJuE+gM6R555umsU6seDVcCRE1QCg9yqrSwvBHiIujzAc0tNZ0brxaiLDof
8wS29b+opwisRRGCvIsDJS3Et954uK/+Y5uSLALs/pHYRJmKTa8Gf57dvzbv
zQP1sSIKqsLvZMd/EGL7whyOP5EqLzskDV/UQe26p6sXP4m5ZPxSIR7opIaW
HRik3dMUT1oVeF6V2RwhlwF9Mkn3CTiVcujpRX8il4E28j1dX/Qw8E/9X6OJ
jo3klwjXgN2JZW1Tlde0OvXaL06lgtyNuKBKEUuYEo9Vb1CtSl7grCZy4J2z
OnmNE2roVZpCN/jbxEN2QF9IS9UBS5C0YztAjKCmij7HasJi5oPyb6DokVJK
re/b3H99I5fIV0Tde38ikT0yWULIYGmfkdcrDhlxNgJ2NcTOdTIiJuUFEVU/
Yrnq8dDv5NsCfOoCkii5NgdiycAyAtLd/kff86DNhz6pxzhpxsy1TCA7Wpgb
/ngoszxtuJXfLQR2qICVqtcm5RtKMLTEll99lBjaAG3uTIynd9jpbYpICIyZ
kUk5s5y2s16BllBDTUxV1aGyMrgeevWtTgCEoLS44wB8MB/GLus3gWkwy3l/
k7KCUulqaR1hbxqesl+Y+bKR+xY/EeDhXx/UR8mfrKr7nNc83/HIVDrL2pFx
kc8okC7V/+Opj9WBm/ZndvyvlIE4SLViSV7SFumhGWN+53olQ3kK4L6ekhCG
i9WFPrphSwrBdbAoOFOkHq4XkCzqRsHSCK5rNb6CPr8Tzr1/WUmlcicltKRn
ZmSZoItgzrY/gD+fQJYDRIsh8JYaaCtLIdON57tFKgSkqbJ1np1vC7RWyPuW
XKNu651roAjxuAvSG9AwSQ5ZXEKYbRM+s6mXLxyGhAvH2PgMWhwAbuuVA/5S
DYGO4yTePfvI6D84WbyzBwvCnzkXcK0j3jvbkGD+4PqAnIfWp+vuW7isZ9nv
BkNV+8qwsEDZcCgmiHnIdJ/rQWHIXxBTCveSmikbgeFrkuDrc10gM1sVSPnZ
o4ihAvNo8e/rVHa3kb3l9WKOkWBRK5rFi33w55hDvHO0SCALLrtLTCEBn69A
lvumyVWQyJZdCgpfSIkg038rQZBHsjZKIddbc8TY2uKVj3YH6VmnuVTOiRc4
VAvCJPjzMl+0Zyw96mgMPIOMetpBch90W4tsmg2rI8kUo02ZrflDOXpO5cZA
QTwyps/vGwNKCbqFhR5TeK2JMtGBrXl+eWhE0NTI7DM9v88OwEeGeL1H3r6k
JQxb/Bjxie0vCkcjEMgoPywBCoVsgCDELbAJH+Ym3cN8GlSKbqweT3TDWE5l
63iCqpm40ErWAaCzJivu9Akxk0dadftDy3GTdSrYqy6EDwxvHeXTuUuYqDEe
Z1PIyAV88N0+o57g5F9BW6pCNzDdZxIVFzCUSdBLy0Wsnf71x7K+YZ1MSFSF
je9h6vyTMI1ThWeMz31JUXJSCZ6tdXRt7kBkwbqph43rv6vdGUAQc35jm7ZH
8+mIyX5UMTCgxDc7ndqp9MTDxCd06xHPMMCNalBQEqyFKVirxytHWMEXXEkI
WK9KiZmZr8IDKPyzkjgeT7khAtRuyKiZKv3vrCD1C5ytdS5MWS8ouk4itaAJ
yXwdtsOcxgUvDtNCpcP9VabGjRXGqB2d3buBfAdmyyvVL3IvujNLUiKZQDLA
aeDzVNScSIVVl2IKbKGRr2+rzuD5eUnney3QcyAPECl1VSN3L7kTqqSGXQMx
Z5rAtGq2kj5o8swQRIigtcRL2J4E97ncfS+xV5158gb0A+4KiBpfW1+20Iqt
UEbu1d1G+tRWHgT4iASrN6xh13FLPUx/zCoBCivpeHABMDEm4fchzOZs/MJx
zvEdZEFAjBD40i8TC9gL2fczkXaY0M2aa7BvCz9PS9Wez4SeJRpASNXOPgES
1k+Z7XftAPd6l9qExbduRuI9etm2qAHwAZ0hWqIrB6NCGZ6PhuhOiw/pKsjH
wTAfAUITUhYDwJkpNSjuCRyLA3ucjS7eIFZj/Mm+GbZvYL5O397wUx3qpY1X
6KtVq6ysbObcE976zueg/ZBY/eyBGDloeyb7PFFWjr85FY8QMHWy9lHisd8O
QBSCJyFhQ6axitBRbvdVcIe4nWhZ/IO0u56lE41P8dVlf+F8gnVxIueVEwVb
MjAGhL2xSWRGDmmHhnYt3Q31VXvkXQr/0uSmydI8DJwP9tWhFnpA5GMIX5Ne
lmcUiySLmhnrjEAOfKGE1e/BT0AJ+RU9XnOYrZMKNh/NqJMalcVNgfUaH35E
ZpGZ1tpIsOmrexQJeN5T/VTvrJmHLzEDxPKzDoO6rQ7DzIqtQ2BBaFwnhzw5
EpMMcShzLl/ewqxzRUOuj41/7R0nWu+qexh4RbCfVuhSzS4mWc9+aw/p5rfq
JA/pSgHLzkYCF3yhzr1Y1Esr6sJ7nGnjk0oTvpBZHZkHZesXRdmUP2WBykmC
ZJjW1SfXGTg8o4sSfgpY2z0WPwuGGbnvs1L5GuUdP7xkLqtmilOw20OtGZAO
wpARvodemmT8Gz5lpJWQMFOHMRLVOuAKyqJfqbAhlcmO6RGeeOxrL1ttPZ1t
hrzrG8s9non43LYFJd7I493sCu1k4N3KkUO4HnhUzSRiZ4O50G2pj1bcBPG/
rVXq0K7sMMHFIPK1Alp/f8By7OUtuZ5bRCD4nxMojf+yX5WH3rmIPPSghycM
7AqCNdOEz//eVl4uPsNwlVpzxNCh9kpRU2j4OT62FlsnqwdbkEfmzqEb/OfU
hXMEOaAoxhLCD+Tb/o7nPGPXbpUuB4nEaVF3Ze9J/6NtLyrcH1OE/LVL7hd3
yTkQOyuZgfm/w/jsWAP3PECxylKgErIOSovtANbd81Xm/lWiSeC3q2Apfhwg
U6otBswa/VDCltwULqIJg8ns2GeU80wjkj4U+UD6M5CvstOntXgaSIua5wMm
OIhv3iKQIiiZEvJN8RlikQYqFqFjd573uZGX2bgi/KBVdXeSRwKtoSpHHEt+
OGs7YZBSgcXF+U2U/7OLHIwdYYLvnDSityvMylVU1fnxglKq7OV3WWC/2rlG
/Q+n28UiZSrRWivvjEKNDc/7l4bCVKUOUFFf27O58k/PNrMbpbSKWuXVc0AF
VBOstDmfKsbSLqj3ikkEq8KAxFF7cp+NeVHqs40Lhuz9iZ/xvlTcGpA1D7CU
Dsw5v0nV4o7RLv50G1KM1UQWlBza9rHJW6UZAiTl5o4/nv7ZC7haOcYUzbhb
UaCK7fO22HYQq50fO7imyrSxkQYuZ3JwMi3jRWb/qWk7x+2pgxJ3+MJ1X23F
/urOV57t6MoeHwZNcbdd+piJrFYLhjqKpLeMS5KRyd3i+DZeefXZhiDxiSln
Z7u5jWq6hzQZIzZVKdR7mKnxiU8qFRpZp4WGSR3o+fw0qxSSlF1WF8AFNwI/
LMjBK2VCqor6L8it9inWdvbX7vDAvax4VNyoFsgu2hTGZB8ZwqW+OD2oWiBM
4DRdfC+LBJ7DSyBDXYwT9OoKOQJMqBzyWRV3HT9wQpXVWfLkL730BEwaH9nN
OotApDw3+9hK8mpAY2qAaVEF9x3c8aS0VH3qtZqw/VwzOwoIOIiKC50uzfvP
xB8uk6IEussg7DvV9Fi8UqrT9WeiE7J6UQnPUkC8zCv2NSYmSyhGjnKugeHK
KsNO2e7zDUqa/VeC6viSR8zfWnKuATAthWWXpidGTQtSi6LbLmEgeun+mA7m
gk+KjhOQbW/PgQ3DQcJnbqq0uX+uoKvCir6hFrE00/EnORrLXlOiNsVKrk9V
aTwsl/+dA0oE01Kppt+CGy2x0nOPKFEW78A+jWGxbUCfec5GNMuLLz6RIGhw
+iGPDpHUprHgJKHGQ/CPXl/efpCb0VHlitql8jjQFeWQCrV1WALnbkjX0d+8
Bx+I6ynOHRlya4+uX+Nlsl0EwY1lrEusljCqm3Owr5nwdQgKHhz5TKKx96Me
x61FcBc+cOgOllXRAMOQaOqvloAHx94OnrU7YNKa4g+LdltN5Qi6XRPyePYy
V4spOCpZ5gt075By/cpTy/1VgatXAWEH4+VAd72bj6gS/rXGb1thzyy4cssR
tarGLRseCRYTm3RafCHWBmAOsI36PyBC5sc2zjW9O+5DGj3qZPNx10OZ0Usz
zgLNYoUn7Qs8QqbZlNtzPotVhDh1v56AY46uAM4KgKQHjcAa6iPQVdMzBGO5
3NE1pOUOfpSKFeFb0Z7Sn3kVpTj+TIbtK4laz1/oz/s7XBDsYQUOmWOpeoZS
Up0nx+4zkLtE01tTscrqQy6R6apxBZliJ+BvZLueAHsoZLUMCBynEa5tUSv3
ls7bvAToCq0Acomd6023L8IG+5JhKSVYqRCixYSC

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzf5SIu73GzJPk9rxU99CIS3AOJi2747jg4LRhFWntS9Y1GkqDpGQIdekdp4xLW49lgfhGPxe451iXZJsBme+vda8FTQqBxq/4WJSyNBoPpEaPEgdeFjM0JpnNMFKgXSrT3Si1hfM77zOpoydwZFQT0qBLq0BrbfuQvK/gPmSlqO+udM1I6asKMA0V8tq083ESGAhfOQmAqzsSSJNVK44XhPH5Xxv7GZHtxrsePFg4cfKUaZR1qRlDulQEoH5ytXmbKcQqmB26Ya2ghy0spdxbthozB3FMFfamj6Q8Kn+lqjZaiFnilk4v5lJHX+Fm0CmF99NSypZzv9eg9FId57eGfNXoXdBEh7AfrOPLRFDXhn4EnZ1mjSJ4T5F2zKzYXCWaSZ3BJX+cxKN78etsyYhGwNPy2kkmpW2a/a1RzRzwmMFA22PqYdni6cj3aArqSa0R5JQbAbte8Op0+qtNsLkWv+rK8xmc21oEU71ITxMZQxMyxOGcYeVX7SOT6zJv8aDu7NLmqvQzX0WCAH+Y2gnluEoe77VcPltpxaCrS5FS8+T/QQ7l5qjaShdfC0xOG+pcOdQDSdXU28wCcEHjS2cl1efBl61bL/Tc9bv39VpsoF6ZZGSgV4m+dGlOJH1KQqRqRsBC5fpzrZQX8fJNfk/TbAWCkR/BMRbuJptJpiEIqOuAgRS1ffRE87HKghmBZNpboVVjpzECr+4wI1WsLl17Pq1n4Bvg37rJKLd3m1zULkWKAP6H7z4Mx+C0S8JurkfJXpokRt0HSMYvPW75YjK8hd"
`endif