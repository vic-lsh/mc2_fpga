// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bYssQWV73t3cWngkW5ZwSDK6XOurtHtUoHNpDY49f2fgoReUMzvmnXLRyhYN
CqQUyx5M4w1m1FHxFfh3eozBYBXCox7SkhVxtOzPCO28O9BgiA36AhMrRo6a
NdLZ3wHQI74MpXicZo06q0WWhvuOxV6kCIam/psu6XcQcHUCgX+8RYMJIZme
OgyLZ2LX6uWeHCluABA1HJ2faGGNY/0ChJWLggCl4/sjEXE06L8qgwRSpJCA
eH6JzzU6HgAPA60N0jpOtKsS+pK6ZDAKEWB/68QV7TRrN5HHHHNQ7WIwB9dp
HTQdZVdv2nPT896D7/Pv7hwooa46zZGlTvFSoovEaw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SgNXcc9QlgnjmvConk1vNHTKiBLk+hpT2rrZbj+vkHiYkStDaKVsRCfHa2IO
a0EtXKUZHkvbuk8bsw2K8PAoKleC3CkM9xCOdKeNZ9Zl3df44UGhEZlPpxOs
OXt0q71wPHSQGcGZrtGzALuKYWrScqMNpwk30AH4mobBd//Ng5ZZ7P66qN+F
WJoahQyUVzj4F+MDq7JQBzPGyEV7fRcQneaHvecYMtzdDAour9b7RlffohJ3
5Xm7PD9dX5oN1B99qiPBqecKBMPbrQb7xJFwOPAJ3vAsPH4eMoD7tcZSgqmD
RqGLKpQlXlQM/2gf4rCbVCDuyErVS+fQ51l5c+HOdg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mzBus5SHyGXwZTqiBE5QrOLcsQzEtg/Ab2n7Nbh+NDpCnxEaDa9e0uvoBc3P
0MexOdMWxcDQxyANCmyLAUT1bHF9zdZPL9ND0C+QlDFnbgsANprHCB9Rs8CJ
P/ra6mJHeqKaKmqfcQ3+JNHWT0OgrNazMis4BvN2OG8M4fHK1kONMXEKpIwv
teQlSd6CNST4Myu4oTkM6t6P89mgjkqmpXAu+2WfI8cWemxhKdZ0AahohMKW
NhtaYIMQJ4h8TjRUJFuChNHsqQnGKpNbsmfdd1R4H5EvLNNQ9ueOtHSDm3s/
xDZP/LfPKW0M41z0BMSkKOKXcQ2lvl334Oa95OWdpg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cNv1ft1lgs7Og/urtzEo15uVlzGHFZPPujo6Px92V2SiJcv4wuiW0uL7MsjP
Ljb7LxZKDwH5Q98rSk0EvQeEF1HiGJnJDL9JQ63BssOcqtDA2cxSuGTDPzQK
oHxolPQbQGfPeyabqU/uo6vxNyfwCnyoywaEIq/4kkAtSv5dJCB6BpyhbtrK
S7DGnq05Uty3wkIMR78r7r4zGcWwJAyoZcEtcrvC4N+0NPuAlsE7TGDuU9la
5b9r1jqg2v+oIND0/1LAMIT4Wx1f4KZHbo16gTDkunh3kSBcMrSsnF++fyAN
llmXs0FCDIJH2nIRYEBdOw6Pcvmdj0KRY7rpqZAE9w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hq6QuGj2OyJHA7wWwFM0gCxlVntwqKREApECD8JO4FeUbrRGbtO+nAglrbcZ
Y3Wd0THgT0/xxW1X6lCE50Ic/bthza0rgoaiNnYigOgTsCdzhVhqlAoQJToK
M+Ygezk8JKwahIEij6frfqJJyseF7snyMl3mfqmenlSmTudA8hA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
o3/+pg7Ex7xlptCezWGByFCgf18henyALZgfQpo7VNvXBMcTbFQOq/XOJoNA
aj22tlV7PUFQvqYHkR+YsXCipjHno8hNBbHzDOYBHgh5gyAryZAeVSdia6kJ
gejeG/4Jx8LphLqlNMCMv7YKEuc/wzOS/svWrm9ujZXE4423XBu/Xcc6egVQ
tdR8OLWAOc9QSDnnkHzlsM09k4ItDIY2U7lN8OI2ffnJwRJYa1tu+fradfdy
Zq7PFKmEmTCHMdFpR2nnSYv7cg/7L3RP0D+WS2wSkFzbpZbIOvor342G9i9g
HXYG1XbM+7XbeXVfFltSBK6apqKlaQG+xDPQCogX/9O0wTbnCJoukcStv3K7
55WEBZo0grZ8bpBxHTmiaS48ivr7FSVCyyQHU4vFyUZ06xPN9pFAUJmDbp+1
coMVm5C8smuLXvGeBqhcuroGOY3wc3j741vuJG1Ptiwt7mDtEI+dNOprNrBy
S7jtDBrcQZPMaudILkyGc1uuASEVyhCc


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LuDwp2+ljEguwvfXcae5zPzbHUssTjXZLl1CO/aE1bfHClrayOjH09Jb9Uav
lNI1iM/Vx4cJcd3gWnFurGW2U+e6pIEhVUWcj1bDJFk9MGJfPEQCZ1SkTpG6
XRtR9ZAOurwrn+J6x3HcSPyPZKaoCxEx/G0DreK18RyG3Vt0GvE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PGHer3m6pr4U5sCxdmpEYhukIrPB1Yt41Zz96fntzoU50ezijW2zSDhyWd6u
YBgk+uBG+twcusAwyK5peyqBJNSMIzrF+2+gV0tg4r30jkx6QF/QXCmWJBgu
Hi/X5sd322Gm0XoOwbItgkVne2syZMonem2CfDIzvICUjOuADOU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1360)
`pragma protect data_block
VDEpf+XppMXQrR58F+8Q/reZgI9JvMsCo4hzfKL27AncDKVh24A0aKRzAdbz
rBWtzjIq+M2RjOf/MRAI+sA0zKpysOOJyOrWXpP2OuaCR7mq/bhIlDXw4J0l
KsVkmIPhrz0n72mXfqaFw7UcMWVI2By9ZdiCfj9bZCVTlREg33KBrPQmB8/e
BYs8P1bYRBIpphGgZZ3mlgFt147OjD+LSP8NiU5nnq6DBAF34oJ22ewdue3V
azCxa5iPhe0h4S49TQAZQq8QIMQPLJwa9IhXbgyceYXLcxnRTUx/Nbg9Patc
9uTtS3k0VLvS76/rxR+hm4bJOX+9FVy9S7/i6pp4e7QhZtiLNmPcC1OT3Csa
5u7H9r33ihVo6s+U7pvtlRduL5q/gbihyLYoPzw039VcKKrfoC+vCExISeTc
Im4RLcSQFSLaJKHRpVgJfUU8y/C9lp6RuS0SwPuoc7RETJ+NpQd9c4VkYQKU
7TQ9gHHbLnMXoo7J0nxcrRmQFq38HwmYtzf+UGGrnvNwVx0lnWebw09Jb0w0
DrOL7BgCsQEIydbgaZ3bS+PyIIc5dKi6etQD4ocnq77iXSdgXm/PBU0cNoIY
8dC2p6W4tJ9IwtZBenTIvR4aTUKqiiD8aIC0kY1lQ/f39GZ2LZBY2ai4k4JE
LmlAzMWHWRbV2Pc0jOK80G8dy39SBJwrUxRn/2fzNWpWVVu1LVttjLRfsOcU
N4XFlKvt2YbW+0YIWl0Q9rXUV5zNy5BOWFesVmDq0KN+K2pZjBam7Z/rLZ7d
KUVvW53FD9D/f+ULl8dlCi3vPYiplfCYViPqDGGQEIQc+Ql5Z1X7To9F5ETz
P8eOZYwnO2Qps/UOAut2sNu08yOMdsbCcKaou+0YJoqYlhtTB+Hec9oZeOur
5shitl2Zq/h64pdYgH+mvgnvxvIWe0IvGaNgCjfzv6CxF7BtQxvCWLFw+YYo
rx7RM1mO5TIpEmlOytoXX6iHbOf8PRbzXRqP5qzSa0ysCBwuaGRaV+fuWLSs
HodObbVQ3L/D2tS4ZQ238Bc8goySZKuFgnGkhWv2BbVmnafFG++ynd6G0eQu
rX51MpE23+4r5u+BD5Cq5vrCfoSWHZaL8L6vLQViyvv0fvKbpxAhHbnJ3g84
qAv+DRTMP1/WzQrzfR9XMy1tMPdJjICGY1NDwNifIHrnbPaGzBjgh1WHj4u4
ypc9yY29ewMCAv9XLbsmWp4i02AwEOQWkvtSHKVad5l0iZ9z0fIUibwmnorz
IcoFb00Kko4AYdLPj8PZXkt9R81/Ff9Mm0/mlVf8eHmt8JW//mgrB834oDZY
/moBoSZLCvdkUK/N2bjWDn+DnonI4gc6iU4co6PEUUAhus1mHS5Fan+1e/11
Y13qthmxXWAsbawFmgRaMBcgpqSLGgClxtg4R3Y2Dq4qOEocpeFcqR/TqBpk
fTwEDad7D90Go3cGgubkOjLxRrr85tBXwVxPnKYNNHi3Dwc08UTWcTZpiQdP
xFRmkAo9aXcBTDctwuG8xZJcbX5+Q6pUGn1XdV491lA6OqBtCf/5fwPqCQDL
TFwIFqhzfGunKtCqdvXlKVXxtFlqxL9InnZTKrOtwftCF3QlkeC2hzt9YHqC
5if1rz1/bHViHoIbgwRJxyknR1c1FKePxpjfXO27AKx4eBsT5tmJI5WEdKa6
ET0zS7hN7165zz4iJesCcGMqynuW6sEPTWRz3nBKi5ozJI6ap2rudRGDHho5
cMVthzNH0pl3mFwOiZFA6cI3DaqAt3mebA9wlDquNedhe0VP5yzD6blIbvPv
oI3k5gncXuIgbA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "w5NDXoZOaZRMdd2LPWz838Uah5+hph+707bnMl+8KalRunv8rE9KGYraslwVSg02L6MgFyy9XCf7XW317iZv7r9DC2kgtnBhiiiNS2vCH/1OQJblkj0K3o63eplhr6TIBGBecvN68UxWVwAzgHvN4JjUslBrlDNoTH83tAUUypf2szYr3Wfc+sMGBU1N2bNoPMyTXef7D1emgYN8UxG+YqtHmdpkJzpcwojxETAcVqfFsbAwQEFRwydwq09UwOV899dYdiR696nVSso7rKZnYbCT+o+//yKSGWZK6fXg9Sd9Seplp7VmYAWodSZJWOvhW8zAY8ZJGD61o8BPyxHej4KkzEUqvFahYbZXtnNr76AJ138L8B7oi4WEqlwZiLKJOVukFJ5JKGtP3sWxL124MmHQ7uVmHDdw0hv9YWl8ZmLobCl/ghLuChkXD0NXvjetPUbSXsAPNzvHuY/1IobXeFlBxHJieKgfHPzQxIb2wLgtJO5iGBa+lZruibTTzM9T178AQKkIoFe056LyF8kAkDxgR6B0wDCd04FccnCufdi1d7RZxOPBA6yjgmB6i1T6oh8JmJbqO1bdMWsczFkPV9+ntcnrfTYl3gpKXo9/18A1dmzFE4lI0+6FL1GK9ohCya4Fd45lRJQRT+5J4qwdosXJYxyzUjJ+dYhrDaAbmkCCcrYXTUwuhvY3BCWST6uJNl1GDt8oyeAfcRlRy5wFVuWvM9ZwS4BV/uzbMszMgKIOSAkHvvg5IsVBFWkzXRxZP/t8ZUXvOcSNMWXHN5LAYi8ZGp0C3CNV9RDFCvroMfex99VZLXFzePHqSLE2oGqR/T1OGkp5jQkgDmW+binz+HbplW9CCF1kFC3b8oe0F2OKRzH3hpY2JyTr1I6PgMK90EcCUjHCW+HXbv7PnqIyYhBtM8VMQkBpXvb554go5C3vCmqNELvIj/bV6Wotxf7zRDfd6CMoJY0TN6MgX0EaWuFP2F6IPLy61PlQxv9UseNnLmdJeEbrdBubiJtBTHT6"
`endif