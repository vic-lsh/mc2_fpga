// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TxFYyuZx9K2ppTfZRVNOGX+wFxijJKtWPujr9iDSte5QK5a5/EAlUVxY8EtA
IlaEqB6kGSpYJEx3iuwYiI1++JFzRpILBGn4RyrJDnIRSwAbXuet9IBywNZC
YOPaa+RIhIytUwtRsremQM85GXuzUm5ev6lZlEQQ2EFcLTcGGDYxWFsOqaro
jmhxhSRdSA6pVZIUR8mXvwX6cMxsEJPXGAydkH7xgWV9Suc7JmhrEyQ2MLC8
Z1rRCkVkfWbYkuBsoXiNVi5oFgCmS3xW0mhwOT7T5aVfuVrW0C+CmAlDO687
tffDVG3sKTEHky5+hWAovhWTl2KCKQJ0gIMQzwjGeg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eJNj8mwDKYmNUwvsenhLgvdNZiZCO1/0IVJAaIMfUrdnyed31OD9EO6YF0lN
dc6Av2Xzzs7X8cyufV+L1veryXmcj88rnN4nJKo20xi8ZE7AfH1MrzsrK5mX
T0Uu6llPXcmavxzUQ7KJxplUxkO3dP1p4qUUR+sltCw38rAG1kIy3D+v68ly
wgKXsIJAF5CGep3/99EgiUNBB+EbbEw4NWGfY8rTBmvD9SkXKjyQROiltVvz
our7niDDxeveMSlMFzBN1Qg0Vs0EEOB8CmuOYyZEty4jh7CS06ps47mp5Vo9
FSHfqVzH00Neq+ltHaCyh4rwBG1GBzV/t09FMZrTxg==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hawte3mbLbEUxJcIgKkV4DdxoU0SW4ZK2DSFd2jI5MJOqi4mRPehzfhq3/Aj
8uT0J+DNF5ozRtvLqyJfaC2utzYq/av9eC/kid+hDy2E7ozwLHV1OTyM8ZlX
S66MH8Nrom+ar/JJSI0XdB04B+euX+OLh9S2He2YfVyUCgvV4zsu54twWteF
cKIMtboTkeuz8pZxLVcJfI/2ANukAGXEd7TzpMiWenzErOopjfm9BBwjW6cp
BLnNF9pjFQx83Dy0icRMlo2mb4xZ7KeFLZLwB3U7mAV46LioqBjjs+0dKn3E
Wf6+SlXMKPvgyUGqVh7PxYfDwizPdbu/LktKlCeM2w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rhtUL0u6aLFV1XrVFu78SEcNrmc5W6OTatmRhLSOTS3qV6kOnIriS+Zy/Yod
G/Q5VV9gKIyUxo8WfSQSCH4N9Q60Q2cfjb2WMWOts1ONmdq+wYUZTdXFgoU5
r1ZypzT2EkfRy6pqeALoCys9GQpNqa5V253/kcf2vcRmy45XbTjfhm0vefLM
9fQOvhyGwkt5R4QnTr7pHB2dJsRgJu+qa6/tEpkp57qpTL7gYtl0DfHFCv9C
aeJ6pyeBeSV1JvaiKuaVpRuMeN/JHN+BmUXkoIe71wTwUrQUfOzjBINuV5PZ
ZKwySTx5Z7F5Y/gA6jkzXGVURsHcdxs9OSb6BmWlgQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ncaZGCV5evAyozKp83fpwRwQX0rtbLhzjuE7gUiMIFBvgdfyqwS2Wps4q0wA
UIiu0wvnjA3I5LsssaJ9/p4O3HDiBl/CWMHLooWglL0uWUruFirYatsGko/u
K+RNwAPlpN5za40m9QHN0zwEFSpEFI6lnCtppdadlLU17A5ehZc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
stJd9yG8pqF4Zq+PJ9bEpeXaIoG2/a3xOnweMOMX7FQV+ZqP9cMn/1/elTnX
LX6J9i/MBVD/uOSUkwzGVU6PUfah9R/oAHcjhdFy9j0/mcR1kx7JdR/bd1sD
NG69zeuFgAO2D1BpyGdtxIJ+cNjJ6IgCqSSx054qlN6kdbEvLlHet4jSGYRd
x5ORycBcXGz4nGO8FnjeYoNhdWbwFoGvyTKlDg8P6gxSRKVW5aOvV8zoyhos
bliKZGcvXNq8rvcDtwntQBauZfhAURXY4tBe+DsTwok4RyVR75WMitjx1Udt
cV/k+mOoev55Mak7OI9G9NBvH0t4g8YiBLPqZkaInS9UkmKfvYnNG29ODD+7
8WiYCGtfXp4090nddwS6wgbvJ79ajq+4Vuzqa/LU0B2Qqo4csvkbRIc6faGa
NEhD1lBr5xQycEZTylw/WgLa7DS4DGwfGYnReK2czsc3PLLJKTablcKM2/H0
9BNj0GRb2bJrkY0Fc3JKcSGFK66sikrc


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kawyZyiymwCsjP3Qw78AuoYh/qefwmkuj6uQUakZ6G6G39ICh/BOiGJv8qlp
kbigocAdEBqROgFOOUcxPlXTEEXML0C5gXEOxedzn8zIyCLOMjQRzTScWiM9
GQe34s+Df8/WvDXa7UpobZJUyZL3yNTOWvu/N54kMPrYhuDmOdE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jgExAyRtFsZo8mb77qprrwfUHlryZp3C/tADVRO7P2ZbYuEsUp/1VkwepPGe
b/bYubAGhWqS3qcqAuuHeTySBWbnJkTAlo+qz+pgB5RX3jcgInCrJE+1A8Mc
rtX4otjowNm5GR5wX0IyfJCGsgrJt5Z+fDCaqCiLZLSF/jTSjhY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1040)
`pragma protect data_block
y9cSeGdlzzZhENPeB8vNstbLBVqFv/o/U1BFWB6gucWzM7N+tGvOq4oYZtOI
vYltiNo+GtA+ROTBx4N0gQuO2glk+t9Zz73L+oAilXr5hTWmfozXvpBfwJHm
VaZn9WH4C2gGAmtOTXV6AlIXF1X8KyJgtycW17kXJH2qzmqkAGg2DvnQ9QuO
zAZ4mTgx66KnvscOXQ3mpfVjuktmd+ZmB6ULCQbHS0ltl+fX2nAAz5s3hR5o
ntIlZME5SQu9tQ3UYPSwtI77k8yYDiWrnzG9dAlRHkOlM3xqPKfD7x2MVNAk
1guam3j4l8rcnx0b2gKH79kuoaCHVQnE3czj/K8aeXDG414uZikvRSE9KrSS
ElUIOhDlLRU+wXiHO3F9m/B01UQTnae3Uh6lnIAjVC9gbp1hdy9422FFxC3e
iabXs0rJPdvwccvu3OlQJcN89y68d7infrFTCDo6U5qijDU7SJFNXELXNHnR
LfvcnMfNjVLkqZYAeeqP7tnodTyctKOR663nrUZMvpI+jvrDVgK6m0cjevYo
RPoDzsRqL3xcSUsOkszQcOXEOSmyszqEGJnvIUuDIMrXNtHnpJIeAtQw0KM8
64vTgzgMBol2SlZoIXysd5VjwBC37uKn8c8qIEJCdrs6mpVRM0JkjYuPGb41
mlA6j3ym+pfVQcIF5qooZo4NYTNinwD7PGjg3GUTZa53Y3eSCzAHcGvxaZsB
dAJCSEjdIogButWuqXCzqtJ1hpzORGq9dHLTAkVE064lgkgUqLrxRw+Ml2cg
YF2aRE0I9qS2Ii2AL9I3/D5QF8OKWVgJ8oc/jSbGD0GtJFosWOqDJy/QW288
PS9qSyIMsuFuQSyeLraqLNG/DIoCJaZoOf8aj8AEzsaBj/od3t3/5w19v25w
t4MzIkm0rvj2gO/NuhUIAnV68QTU/ZjuIUc2aOfxWLovedm7BYLRudqOVZzD
1mgNzIIeKt/bexnn3hs5fjf8bjMeCbyO/A0VQRV5hWaA2k7ZZ/Svxe1PtTC6
IvJ9eXEOy/Qcbs7exkSKcdb8e+31neDUQCuHXGAkXQ/XpOEAkZoJuFkVMa1p
d2Qq44WE4QVZ/LZXaPVyAqLLtNI22P5hpzJ8O98RqkSWTu8sW7VwpA6Goe6J
E5y7mnaVyRX6o9PUHhnD2Y/HAuRBtDubWsEw8xwnFQjZkABn2aL7oNrOLyMX
VdUX3gLiMS0Vl9LwrVdoo4ZOoOtmTe3kPrPO9etDk+AzUV6fxr+Ba0CuqXtq
oS946UDo5EyP/6iC9arxb1EpJMJ8NeTUVkmuLXGz9mgA9AfoSywwRZRDIupF
A7i/JR2J0i09TM60GcvHnBbjEQzDr11b2KRHVTrn/vVvDkCChtzxBN0YcOWO
CRqSIVE=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQoxF3kgpWfVy/zTk2XTFFGFYBqcFf9woMESopIumACBTzkIvtIvYdAE7hN5yVWoC+EGCiY+jeo1wPeTmrBpHtfMEyPF2BFaYuEE0cLSuxBKTnso9O/6gvPOO5REvZo4T+E/dkhAD+MzLBxtxcDNu/hWstvtnquVIn1a3otlnTCc71bTdpHXAu9+w+T92Amx/1XwlXG/nfps56iWEQzrdFBvVE+ZdUCWXe7bDzgmUlis/PTW5y1DP0E8Pz2DlCQNsmtukun7sM4V0m7xb75nKvqKcrR3MN+87t6cn7ow3Jtmys++RdsGI42z6cHLBfTh4wcKOmTDvpNR3TvvRzTWBrG9WXgGRQuePI6qAIJ16mS6pjMZqfoD0jFdvIJ3U/AYLf3Y1bUzcealVur/0m6lsoX1cZoQ9fTRHQ8v9sglDCQ8bIspUp1RNQMEcG4SNDgX80BiGgrlMPiVjprdeLe9Uijz/Pj15hvZ9SLMyWSCGf2+7vvfNi2ubd4ZNmNCZZOfIIu4FldVPguu8dhVoJQwe9ZzUAX5sJjzPjVIODnXX3gqnWBsOQvtO6zNaHaIz3khx4u82hzPSf93ZH/t3gQhj/gdS5ybtMUQhSz6a3TqelxW47WjOrI/pOP+1OSE0TH6MVBBtXPlvMQjFFJtu3Vs7uUIVKRc5haRirCVJ8wW22XxthK4LZPTQTHrhzlaak3aUMvo5m9lLPD84AJ2kDdP0VqHi80leif+90lVuWeCJhiLPup8bMc+6hvvXC0BcOrdK9C7M7EHXjZoa91zYVbB2qmJI"
`endif