// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HFI3nsOoOf3cMY2pCpI2BhmkvWydMJLakveb6a/aBM6hV2vaEMSCbfeb3rVj
4emIphYW18xWx6wcCG/S1CBALNyR1IvnhHwcBKM/+dQ26sj/eamrY5fq/Miz
z/EqKSIievHfN5UBrHTalwO/BK88XxIDoA8hQjb/wgCSMn+b3Rb2LSISRssb
1fpbECbPbt+9saaURQVFD6W53BlhW5C9jhXHtCg0Tqat/LUCh6kgyU6ETgDA
5uQv9O1RlojKoG+HebHLVSFbtDEkyWQ0le4dC58seGtIF9yjqHJURNHO1Bas
/9c431L+m1KoeyejDj7tHbwvapfpSX10/gbE5XYsmg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PY+kLfZqwXOxizFqRq9p024LDDAwTb5H3bG6rsKl7P/QGD2rCmpPEGpJVZJI
PpRqUaVKXTfkypktmI/P0luMbecIf4+Tinvaim4+hCtDqUPuTmSjf8vnDuwL
yR0l5xOEjEMtM1zhfxnf6uW/2FRNsO1s1jrNoXciexXaMzaCBHaWL++LwMBt
GIXxwQzAILv1bHheM8w7Dh5s8D73O016aiPXYpnJaW/7cPKBvbHw7+bfj3Gi
I+k19ug1FjsO5yWzD8XWpJ3wExR54Rxj/6AwqihDn3iSi1SyTxkMayOdUjje
Tth65VNzrjSVa0hw+agA0AuQOp38Vz9QbBQF/bblTA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZFkDiM0IEU14/OstPdQX+uKfZek0r51NmecISCuSA8F75kqOw9J2EqhTFuLm
6tBGpMzoxSulTYzuijijqoteOR7UD7oxZhaBkFTSJul8G9NRKcK0/hs8luKd
RKnLYklA/IkeCamkUYJLTYpEAa4mSelAEyULXWbWYKQMo6MH1rsdExA3bkPS
Rm7DKMxeMcXsFVfyoXjzOs8jNJXCywj3g9m22W/1jlJ1PBhWZM4cIh8PSt/P
Bsvqo3merBY3LAP+thmFABxwbp7isK+F2JhJHtZwprnMqu6uaP2XwKVI31gj
tqwvVrAb0cFrVgGXNoL9Hj8HoyxodrmBH2iPlQlF1A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GIRquyKWCDomg5aQ/lioHdYRJyvMWh9XrqdS771wjdPTDw148SwnA6uPWvxw
brG+GRkPjQMVU1hkymtWSrbhUzQ4FHLtlB1Dx6PzkMQWBAriiJ6OF2gQhpK5
cDTauJ55KSu5WYOLYpj4pix6w3qyiUpCHlQXiUiUDoMQaYmDTqU/xZ5tuSdo
0V3OlU3XYpRe+IpbPgfXwvnytCr0WA3Y6R7E3rlg4f2qiOJj2ZWCDjd8dEQf
CEG1TJiQMFfg5JJdAN1VytYWrRMsVP2gSuud3GlHpLPBqlqzBKanWGjvvFeX
VHjsxXqY99yVDNqwOHCEKxJhC7G/Ul4nd73QzyrNmw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MXCk/PDX7l2IMkvDBbrMa+V3WGZUzHU5F2rCmsLN11g9uWdTBByJRzGzI1Ce
N9Pb7ujaiaRoYZzle6xPpJB61FskKDa1wcMb7H0AuK2kGSuNT5oK7mOarFcA
uJ0rcAJ6bFnipUEutCVjuYRe5bRiEdhNyPBfgEb+8j+/Rz9MWCs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ke4H5ReKSjvq+wVCdXGUEwGXcFKEvCMlHFEfejWNm0JJc9SLFsYdR99A86wn
bWvD4rz0v9KljEIWlYnWBz+PsciX2S2DUr5QbizfU+3z//vt4EaubwoDLnXs
Ol7DsYZSCeXGuBDSypJ2br24utiEjm5usmsvY12EOESmajocA2R6rAu1yc6W
gPXz1m1cTh5f04stQe3rD+hn2/cX+M/DJuMb77piJHndHFg24wAuXBt7HP60
wXOfGiiXjNX9uAV7fcjztnMQ093BlXUoQ25XzBL7hXKBFx3U4gAF5+wf6DkK
I5Hx+6ad2i7T6GdrJPsa6OXPIIvr1gZdh3MfJkkydk1EGfrVimdqtyoFhkOM
cjoHMEYhnsQecEVoZoONdVsFRVOifl7OUdfxzJFcvj2Z7RrMQNF/f6tfaO21
W6oGV8ObZyt/69gt0o8nmzYvI1hfxx9hnBU9QlQ+h+vUnafSZ3DVFnixJkbD
4St5YIV4MJfOorRaTam91WDxz8buIZDS


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EyKSNUqVNaIuI/XO3PMFLu2XrO7wH2sZBqA06XbeAybH8Wq2/OD58Khg2eCm
O8ieq9Me+wGij3ftpvqQ4C0hTVlwkHr18BbAJ3seJsAo/W1UHPhbsKaM8bia
Nf4Xlox4TDe1cr1kx6jfASV5/73sI1eDkRziI0Cu+5dOof7Zoj0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XNsp4tbfJ9jgE+J9n4MqVknCwxxG50q0613wQyNi/Rfoq4XYjKizDFUg9H9v
gSVxLKZz6uVhHn6Mw58h/jij1GkyN8LHusIt4mNE3vf1NldLtOnwhqfUTyMp
bJve0+5lGr6+3lmH5y7tqwASfFiwMWFsEpWmKl+YGq3IcFXHCvI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2320)
`pragma protect data_block
cIKqU1AudZdj0OvBE/s1UUjigDmn8sJP1LUNhkWtaEPp37Zo67ASO2xzD6T/
CtDSu8a3u2Ed85Dh3SuY7aIEfNz0xzFgcTd/TvkG5lf8vjWkV5+tQvlyFph/
kvXJ9XRNLfV+pz+VsYs6JoRWvkqM9zxJKZQrrGel5FZVmNfzG4zL5+RSbY5H
yMIm/divy5lNewDB+Ou1xqp8Vor8GXx618hSXNzYmyd3t8Ov0KLYLfub2CHk
9prhUk8z/3lDjh+hCl5ilGokGzouk2O3fE7egGaGW18qe28rFJVhWa9EjRcd
KA0PknbKcwh0xQlY10vg7yjoePSbtWtJ91a0pjZcRHBJWLLnD+/+rjur+Oo+
DcZo+zZ8F6zV1T7q8L0CYH8tuFuUD2ABQ/clWWHGUSAuQWral7gvpNAapUPX
wFfytsayj6zlDqG0OEeZ68FCQ4zJ2xdu3zMywYbAHCYBgg+BbM7t/LpNUwd+
yK7rUP+fEV+bo/OpOQeNU4DJqTdodtc3sdREtzH9HQU/V8eX8sA3clw4iuI0
de6gjsj40wWcYWSa0eNcgHJ4H83Q5V69mMAPHWKKnJKFXs0pxDhDloZWyvod
HoXAlGbJXOHr8zrxQmI6N8e6HHrqUrPjoLXZRfW3MRwNjeafrDOc3NiPijDy
u20U9h7T+PCWEOwusP2breUWpdvJvsjR4UuHMavXtTRImQH0zHpN5MmROvUt
tgNz05qw50h+wf+KH3ncyoFKP1C8FU9tRs+U0LuSqFcbwbTAvcujsfSPfrBN
4piJEIgrbGH1GPVrQ7X1B34l0bjUHGf8XA6PwXRYtcbM3glMAlCdyxY4HwOB
PjaazZ6gHPV0Nz5gIUlCc/Di7BX6XXFvijs0L0Kq9V6F11UjJwVjrhZ3CIZh
a2v1ORk3kJnsoiH77tNESylVGinUtUC4hFikY0D5W+ScWwNng3r7I9cPaYC4
lZJRAMYh9jB3Rs5hcogzul6rFyTz0oDbYEyeR7nlCW7A1GL2DJfSmu3W/G71
ofpyW3tektEbE7qdl8rWcAZFbc+/+7E3VxuoK6nhdqvI8EPp5WaW0+UBdckw
bToNpGNMRQKaj2T+0ZM1l7mAChWJY0yiLRD5PBrhhVDkYk+lcOvx6cRQW3pU
xpmcmnG9h6BimsN7OTPo/B/H/Ahau1dqsRBx+lJjAM8fuvXOtpeThVCxDxta
HYVjxPqNLRRLhqemtcWtEwqqVAAb0Joyk1Q4YAhHXFpayO1SV0BIVGKbaKis
m+EL12RGlvmtRkIVWJJecFQmoYGQYm4c3PaEy0xzLof7d3ZSJjB5Fw1SmUwH
q/7diHKGbf8bNc1Y16qCr9O+LyI0oYxqHPKHE5+0iSSBGEPq0k4QmX686CH9
RYRFGqCpf6t2eCWHm5yf8lNPu2IiGmXy7ZOleZ96lXBOFo8GV+tqjX2cKaz7
awCiXibu8sluTmDH0O7PF40c2OaWrtAYme1A7JFnR4ghEcwETx/n/P9aaw8Q
UxmeJq/J4hmkdBLotrNam8W/hoain1NFmaPDeEMa0KwUjMRXv7tQA7tWDCU6
ucOsXePyI2ROaYlVxscqueGwyhUXpPgWy7Q7KLEpTIYV4XBIrKZvsnXYdDRR
852SS/UbNDBG8hSOukHyYau0yV7QbaAicHB4v30sZgNrBTYlThq62rRNt/db
s1425FU+F6Q3hVidVDgc3c1aMuVyIr1A2PtOxy8ueCPhUqgAiFwCFzr8halp
VnlAA5FoDS3gDIf8dwqt9IkQ5XlZkfLn53oZFIXhJj1QXAtFO/OhsyQORodh
nu8yDhEe0q1HK9f881KlR9mF59gVB5Mq9BdL/beGK17ujasY/QsU8pfAWLHk
Y4mqNRKbcXuwNkyOMk8akE6pgE36EYXvqFtJ0Owq6wjm8TiW6a/uFStG+VLP
2Na3CAUPS3S+xzojiCCNvW61jlcJymJCm1/j+COqFfsdYRPdhr/fvO7/rAzW
XWyriTvXHWZ8gr97XE09gS/3ROvhFkqkYCu5rop8r0CK+ry5/080hD9o2SIb
kKSyGgrBF0QxkgteTkD3cGIC63z/mi05+Jcszu4uXt172IXf67wIDO4Wz83k
Z03UBrvu6n9sxWceH7Y1IFA0nK1YRShUjzx/6gL3qc7dejNjQRN+YI+fweeM
MRY2pg0CLH05e5oMokqduZdCSNmgaYSEIoIG3opnRYJXaUDrUi/qQ2XLDEcY
iUBw50ViVREflZhJ/7rbnDHXq+Ug8to6LLe4n05RKl/JcJLyaVhy0YVZw7dw
D+b50KkKM9IDU/NyTeU2qTjGUSNt5FmoEdcxA4F/Ts5rjK3TXR/jFNLbR+fN
8w39X3pxYiFMfMAQgEJ3mdVIBJ5ikBbkOIM9tqzmevYxH9F00eaBG6ewVAgf
WYeuZORASyMaTh8CTvv6DBgq7zmxTF/FYh1ebQAK92gsR+wNpZCoI0+jzqjW
9DMFspjFufP0+Xvf9HCu+ab4jiuzt7XuqvpYUJr586GJ29zjQfm83zMkTM0n
vSY2dnFByoeeT7jNwJ3p3i9wYaajQdEpp/c8inhukrPNDgmD6+p1Husmesar
l1RqdtLpSgEsAnZJglfNhNxDZgPPreTf580KATzZB44hc2kGj6o1Lti2bGrt
G8gZdlJGPt5E69vtk0iOqdeW4GIGIwbsxx6R5W/br/lpFkah3tZUTP/bF/iK
OOQoy//3xV7Ld+zWrFM/2k8O/GGDwsTRrsTcNJOYC7iGaIRctKmu+3Sg7JxR
kPxjV3rwkKLiHtNaaU4sEXYUKbdLO2QLuabf24ulby6izolmsabgFLZI1mqH
xkGvi5G3DxHYLG1k6kkRaGIiQmw9P5lEe39AD2RrMOq9oBez8kNNR+VmJUMF
GnGu8R6O8+7AHnelm+a7FLJ7fROBfufgTdRpmP03ndIeTi79Vz4mmhY38yNX
eqkifJKCa6gnndFjVTRYRpxKwhU9uIzjp2f7qI4odtRkIYpzNkWgu7qxGfvg
FSxo3Gi4gQ+NIUn4dcr3CroCRjJv0bbIJVMiM+FbTc8wzeTlSF7j0srUL3iC
FSwlzKYacxtuO6t4PziihxiW0B8hro0U9A==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "otez0kW9mi7Zi12YAMkjasgIAsBmZ2uUssuHYIkyqYZwNXTfDS0Pzy9DPD4Tah/RXM3x7fzV3iKBSrws9MOStn7kJ8z8r+VUJlSSbSROvX90gAb3JzJzvIlHHyfYW0HDlSmULJ7AB2pabuItYvXEDzTkfhmdj0/BIPNDjGSSGUegQQ9keL9s0N7tOw+fx3HphhJzjKsOTbe4+r7joyDxoO8ldNXcNRzcMdj/Lihc+EpUPFiZOIggZ+qSZRxbn35taNK5RPv1kUBe7x2duYOBwReBEDKSbd3ukG8Ot04xpFgz+ODDqC8mASrH9PXSprK5kivIm27t2I8l3yp/6dP//dxsf+VWvJEb/OLWV3LlUhw+zAi5/WJe4AbO8PEoeBUq+s/i8eFRc2NnLoAaquCTetUIBEHAvVR/VM/z17ui7+xAxhvi6aHXKLme/ERxWjh2xsnQl1Y416joTFPobFaDS6i4aluT8WxP5Sjbj42A0HyVwSNOu3MqfnoPoGbRSaiQ5BqUflcVS8g80yCSK4p1qKH/dxJWkRurjeOKgba4S1pfeuaZf3QpuedFLSQ3+xWIfp38hY73axwwyHRW2x0fhA5+1xLYc4jF79QsTdhJAS5oRYT4l4y6rSBPfwLvOnbBVGhgnLydLLgFBd+4BFOE+WzBy08B8/Jhj1LE9sUiqlx+SiAXxGNLsKrBEaAAgutPqWqpq4gtE0+JjhzAj5D/47e2km6teWoMsm3yL8S3oIiNJX5evgnKXcrBPjRb/bi/mpV/xkQwj0t2JFTHmQauX2/6tUy+fJrS3fsmoAdyXOtkEMUz/w93F0gGhsuh+MLC66yORTlbrAgqmtKTGp2fbfRft4o6aGYoNpgbPk3FFfcnJnaUWup/Ois3armwyMJpzhgpIpzrxwOQFiWE+wgnQTyU7KcOntwlDoBybxvvN/BRVyr7DRgk3pD/3/c7EiURXCMVOgnhkY5CAlsKFcbwHBGCGK06qd9I+mDMYAZYiA6mbcXlZKkJPGU6dEZAijff"
`endif