// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mQuTsN5gK1HLZqfp1GHu1aTCn6w0/yW+hnoh8P6c6CA+c3ynUhE/Lvi2kNMB
povJE7KC70joejo+E/WYN/KkA4qInArz7ebiFGOzDQ2WzKv5ll90VtGcATE7
tjWwGKkJOSBg8862mgVTZjZ318fZDJGqkuP2t3qMjrkPeTVBMElCnJSKh8eW
N43FfasUc7x6DO2+f8e1ugoMEgM6byWRzrdrdmFLd36o/zLgMHt/LlaUHrZK
f1SqXnkdfY7AeHYXCYWFzem796L/nn6jUJ+jSLj8LLFgTjDVXCwDZVnuy+yv
crWcH5WOVmWmQB1YP+rysYrH1+/GX1Eddk7RLOU70Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VRNpWCFuP7ITKoqSSW668RoyIT0zMk1y9lcoZK/XRU3qvco8zPE0Dh+4v9PT
npkoohV+0/muU7xQu4Wsbm5+NYKtj/gOG5J4bQSe3XTTd7pAr2Or8bZ1kW+R
YXudfO3GuBgpXLmUW5+XwCbOTRSHee3Ygd/QE5yaB1YwnxI8yPHktdg0q0qL
2XNxFqej4rdBLZyTQYwzlHKWd/0fsCfta/h1Hmn/RBNXnAnMESfkcIxBqNsF
tEizfvblL7MmKGE0jJw0q/lAXMrx05LdsnDhE5xAaRzLGRXLi050F+hLKFlQ
9hl1v3b+h508lyKh7ZUyROlHgsNIT4Q+MXjH91plGA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bmZXg+SNbDZabxfB3uwWJ/4/y6++rgW9ra6QoomemhzvgrLVy2yj41WaUVmY
8FXmAQ/HFdnBcVAvm8y9N4pqPap+P7ORb45FCI52sGsDJjig7StqarIUhs17
Bd8bLu2D+cxCVaSy1LmyKIMDT1sq+1rSJWoNrbdYvI93wcR3PgDU2r/hVxih
oVpZYE6KV5HPA+ON17xwCWzFV5rvIgtjrzj03jfsLTVG1/q3++Gxur7ssT1X
wpPdTf76SqnUz4evi/LzZFaSzWTR2UmotBkz4y9s9Y0XldSWKIxt7bAwFmCv
/Pk2z2qhma9ujZDM7E6jDxyIM5yuNKpT3GPnzLdHpA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Hl8HsL9BghP+vXQrxUVcufWy7HlNJ6jFY1BeHFTzVrnuXArCciY4Nm3piK6+
D4Wt0o/4JjRUew5W4IVy1IlUunLN9kSUyrXqPCxgWnJ+y7O6/iXSGaIZ5171
tdSoZeIGDROsJPui44p3GGwjun1MvS454V8qtIfcTQcxoiOrGrNyoZbr2HgC
VoLmjVIrM4D2Evesfn9OumWbqWykPeO2lZ57pE1FPvLZWbmA70n0jpYL0GLj
DDd5CC4TvNEHPci2nU2Aqx4WWvyHTmxGd4fEXcwDjb5HxaQylh+AqBdJkguL
jgTUZ/KahoJhen5NHI3BGs6wfOxSDYoINYqxaycJDA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ElKznQIOmomoHVAs1znVrMAi52eaktRR59+bMZW7ChNfx0i5TR1HlvNTvoTD
oOib0ZbmTfsWIsPh0nodBE/Iti/LqvIjnzIxAlbMLi38dPTLWV3WOYEqclcz
T03s9KtHT0fw3tDUSKqy5dqNVLmQiRZIrGyoSJmWerVTFEJCwy0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ybkIWMND/RrApCeNHncMM480aNJXm/a84jDCP5dcdw63gDcisDNG6LIWtcYf
hWpYNRx0O3aNUjhgIeabgzkQHmaQAlNfgL5PsEmFqDX0vxxnAy92yTCfZO4E
wuo3fDKke0rE6vBTu39kaQlVyTSIbYzlbVpOzwUXzsNSK74e6LLp2thZA4cT
vWY4Pwm69+A/UeMiwf9QCpL1B8hMZlERPBugFd/Mpg8T5+iqBoiSTaeJkWN6
82RorPFc4O3TEEXyD3isCBQhogSgp9Zbq6KD/QBDt2mfCgI+byDSHfJHtw95
1zPnzZdvhHvxoz+xOYWfRdlHadzXcA7U3tIeA1X6wotI56TtPuU09ZdGLDhG
pHMDVP9gYy1PZuHX8aLDkLeZU8j3PnFxagwCDk7UHmvnK0w5AjaCOiR7RxPs
L7z5f0/M5eMmEwpEEZvkNrbaSMd9yiX7RUEwsM+OUM0be9wmw1Q6OtQk3t8t
ASKI+D5EgFUkgdZRz0kreRAxvJpQ13fX


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
h1bQpsc56R7IrQWL1jk62nsFo0h4d9cyU8v/+oaBAgOAcey0ZFcGwBTgl/+R
jKAhYfpuf9quAko8EwqQK2k/Zo89Inp0fXmTqKSGNb5F5BLRtX4F1NxkA67g
kDmPHxbfClZ4IzPqGLbrfPPB1L/jK7UXjlpWlnJEejLvLe3pHww=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kaLINBzbJwMdGpmUwLZYj1f+DTndsOvqa7MiizC8pld6MjAe1BSEbeIoaKqz
PTPyCeT5vuarAWuC9cydOgw0XPXAJQUi1Bqy2BhXYoiwqiyAWPH285yfDWdG
cnFnZ4HLOeAV5GxRl+RwOPrXa3oG0K6kUtQpGAF97Wur6fCGqHU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1312)
`pragma protect data_block
cJv2DDjBvIcnfYxwHnvSujSUPcSJecdzlOtik3rkDZPZHzxX7uAAeLpmnYIA
4hx/hfYksPDAasq7pvvg0wqCHEfdFqJBGhqc8/S8zU8XUNXiNJoABW5wH2mP
0KBxTIhN7b3Xrn0Vve6VzwAgP1NyVPDK6MU1tj1QYNIpW4mQate7gSIL9sqj
QITx5eWiPzLW/GI6ZD/cllUAEmf4elOzE+fH792EIINfULUa72QC0B3yf0Hg
rQNLKD/gb/8Wrv1F4vdfjeORTvLtqSRstWEiUwQI1K1+ADSoYARYDcmfikIF
xU/Hs6CwjeGOvhjOEXohEHat0DQRfXCZng2rLRAPNw7B+E2n4I1V5wbslWL1
4Ps7rQzxzMGoRHI55yZAhCGFXMCKK4AWZBEhpLXpC8Yrzh5xfuFmsh7R4HCY
ZeVLOe+FQh5I7yxdnSpkcR67KzYiXxUxfx8WKwebSWiTUxX5uJUG0+w86rg5
y5ToiSaxnMiJ39ShLmVPVE8xEb7w99/oUTjJysM2eK6BSYliZa8ke8XtNIMx
7otJuvIO/VPBdCvGiDE9pw6Fq7VKP2aPCgipjNMBAK2B8oXLffO1kxjyJ5Z7
4+1ekOg++VXuY2N1HNhDh97rURbNx6ZwiwRQDrpQyJxv7YjLBVWDu5r2wt2b
oMIxCDPAzYF7H9ZhSHXnI1+RBOcv+WhLT1ptSC7zF+4ixIPJA0jz918auuBU
1mYpf8ijW5GJpwb6jY+Z8imeALs6cA9C9aZFydGRl2xa9cS7/XSR3Ar66UBp
R6snCBwNylemPo75rXCeUejxaDvRBOtpHe0VZnwsczk4zbKc4FPCeimsD8C/
Fx7YYTbuvvClWqXLJi7jt/DGeukZwkAOWm6+yugu3D3VvpMomKnZma6MEzJh
iDl4BLYO8xOveuXeghYNElTGTU4Af8K8wkG76IPbJJNvksthu97r08wU3mmc
ebMDJCbRFVGQPWzuq672zQHKA0nvUs7GJKO6qsaXJdXl593Mx2y67sTZjJSa
xODnVbvtiATqeL/OHoGkSYyljqaBXnJBSjQ8IIP4voDhFnWYtHNT/rnZB6Rd
ZVkHsBhbKMIUJeEjayAQnYNJ193ZsLsxoV9GYM0u8cydNWxQYq288rjH7kJQ
JMAtj0xWBjql0AIMAyQ+SuyP58RxDMf4WUNuvtss6vhvr5kfgCayE4mkghQR
JmsdCpYD8cJ7nSYTUoKKMcle3XPLKf0Q595OjW31GkrWfWsGvhngxLR7CUhx
DmJjArdFCZihak2C7BjczVakqJF1xJ3VO/miY+hiNEemAwlBq98vInavUr/P
JNDdFmhYNjU/90sMaNjgwSDHS6RMvpZIW8Hr+LRFkgIauNGnKXuQ9d/FHpG7
FjxuFkICPMt4tqS+tQa1GAqGbILLZXXuJzzhB8HFTAO4jOFWZsoQb914Sz/C
1BTyvm3VAAHXcyYipxUlqKuN3N2nJsKIN0jGfr9I6AZ5PAa1m5jW22XAVrzY
KbqCzA5yPuq6TjqS765popPzhTfb+L7yV/9E4a2Hin/CbhqCAuEE0sSDpJPY
tzLXuKl+qE+nqSq0+nFzCPDeCo/adwZRrCFlPYzEgMkta1rFI4jYC8Txmi1v
PrzF8uOCwNfeV/rhauwFeaQ7LTSwnReN/lbca3ACCJcJObpLnYiIVgBKgTg4
OG6H3xyzBeNjdi2kGq7XofDlVXV4RhOIZmYMjU025xqlClwJ1ZFa4NwsmcQQ
g0lg9+SXOQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fidd1oyAhusLLJ6+7Y4fW+UxvqV+8TisWbzB76p8J7jCbedVkgTXiBKrUzNVBIRDckfBwS/gk4qyrpXnk44TsazVN20DO3TdF1x8MmH2pGcTjxrJqgYV/z3UJLaYPiY1WrKUNRPOAuHkyYvfI5GoAsKohhmpB04sGLV6+cGIymx/RXK+eIUgAROf9S5AOXsk1U/Lqv4gR7i2yfj3c/IhJWMX+Ld3X1LJ1lp+Ly9OQowrepytmThE583kmRsWwT/WTEkS+gnmNoQh2zbr7NKlG2X/ZKeJUNw/+rRaY0aDGUdZdYcEELfRjEQlzjehhHD4nWTF2x8riNBRcqYbkH3CajdGHu/nk0M81JluX1vxHfEF+LO998ExegJOZYODLRt+jfs3CoI7yKxj42crGo9Wp17PuDJyv7iWZLRHYCYsN5EbmGg/m387fDM9UYj1zJe8Wv/b2qEfFCdQ06omZRQ/O3K6Ki0gxCCK5BIttNDZj8c8nKWaKiO0Ndmfe0YZPV+FToMR3OEItt8ckF+EVd/x6BokbwQk5Gte8nfmEIop6SrweloljDc+g3L1cY7kzmbdRdOo6m8wuWFx+Hu4iodnAaiA9sPw/Qlneq4Vw6kJNbLMqlYoVuocIl03kcIOdyu8JvRVMlqCYCrOjlRCAG97mi4jqRf/MYejpthLwIrxjOG05GhDF7mbcjVlyN6GtzQipRimFD/RkiPnGeuCUoAzx0cG3p9tvpcov2LVik8wkjZkovrpannvywvG0A63O9j7OcbiNfiuQp5f5NMBPDuRbHqT4Bn17+gGwn3SYNv0moT9lJkuYbSoz3exxG0p680Ng3+1SEVMyW9oZkgmA7L0lMwLsZA2igRcJ4A2j2tNm+n2E7zqfWp5cIiIIJzIPmAGLub51WiZFCTKnz0qQpvv1eevBwth9uZ9vf27q4N+bmYLRWbSlBWI76AIuKCGrUfYgOjHzjbKHQFPuUQMExHTiXfF4xjtco4zLK9Mj5Q0UQPDbBgtCAKxl/22ZZ7e0TG2"
`endif