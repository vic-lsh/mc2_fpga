// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vo/jyxrCkqM+Z5EIqeT3WCf6GIPC14+RtjsrjphaM0847Jd3xWJkKKp/r/fb
1qrwjU8WNa/jvIWPyiR3iq+UvjMttQrnqVAFkyWT6zCoA1ZECpOKY5NoyHsz
FtlbvVpCJuLuEE3w7fe/wZjpbtoXUfDULcRRluloNEJR5y+KHI1s5UMTrQYq
/umNjGBPJ4JKHVhzJ2HFdu4bbx41PIT6cRgQOKJ8GbTkZiNiIOqLdQ88Fq/N
1CogReBjHT/MIEH55Ef6xbxSCMr0g+E2wqT1xGwkP0vzuh9gl8tBKysr9ehp
Dqc/1ts9ytFPunQQtoLxi/5FsJinZMfO+Ukb8zTkjA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EoKxMCVY5oCul3E35j0xPl9bo5XhtEhUuCQqUPasYdNN5wgtvI7v5dWWm9Y1
DpNyJnT7TyNB6L32S0xDe2DePNIvPDbRLnhPiDQSpFyv4LTzBgQRWsjsvHOD
NzGGrLl1UYLv+CC0ldWgOUdIaVwDvjif8lfZlY1b/hDW/jz29TzLmbi4jQ+I
DSGyg+UMESdQkpTlq722sEkH36NzjTgi+3/0HiYy7pA9MhUnDNXrGQoy/aUV
OWWH1cU4dYOxpWTypmOtFzgvJHvRcCYyC4/Ipr/hkQzNjY0rUs/6/IJTIoHe
XL6O6YrFLqBMIiN9CQk5uwadXJjR5TVfG95jgsTJTw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eYYXNHKSKPQAsj5L88Iv0QQPD5GnAmu82+nWZNPAZcLeQE1uapPaqgeEN5ea
GAlHgUEwjrYv+BhyXBXAfo09MuuwJ+DkzVbO5iAwnOROX88hMhK33jC5QY0K
6lqCrV/mUTb8pA+lVpX58XqvZfbI4MsS1xt8yELLoZQPFzmWmYR9/3+vCXba
bcbdWUsDZHbKvRQxBeydLcrJE4wMgwyAnl6ekcbZT7JXe6b93mHVjZqsvrKA
g+5r+vx/A6KVytra3Ipq9539r18bYLYZLasrt6GYAsIU18+WM216Nfz3eZUt
nhFascd9epAYeBjFRulzVX5mypiHfVRBZeu11o/Lxw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iefVbIVAJB6+Q/dYmYmoZeJwtzCdk5jXE3T/atLdMbwm4BbPJsW5iA9tXos2
AcLR+4G75xWr04JauyxusenfygqS2QQyL4Nowodo70odZiDUdl+ZQ9CldKCJ
nGrs0jow8qGHgvli4eTqwxTEs9UqV+ZRPrcDVu53udtg/1TwCcxGp+sRvIPC
8lJJ63cDvDdAvcKFP9qicpNu2p3A9/8Qqhfj4WOsNr1eWiEyc8x7doiKba9Y
sQthfZY0DccHKdCrT93WiaiWGcRps8ca1OntSigd+AqstqgvZbYqda1MD3uO
RBQUwbnba2iXB1w87JPqEhdUvOJsUTNe0UujwGZAsw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KNDXRkNISCLu7mPfovFOeAYwWOyXg+jmd0lLLM1pYnyRPgl454oQZSdiJL+v
4/4adTrY3wjhno6neC/ghmK4iYf4WRmM0lSOpLbK1sClc92NAy8AzMDXRJUK
EU0menujfotT6uUblf5Cvxn2i9/0tbGhf18xLNck3eDmRHJFBOc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
lpOyDKBbiW2NIxgQaeCKLWh+5asXRNQTLpTCbt1Ub+GQC0hlBL40xUvIKxHi
Nbv8op3oc6HWOWB9H4oLwLpWUztql+mkWUYBdQrxlOzQTJkFEyE9cKi+39iE
F0kEVwriE7PwPOHV7Jd6P4LcJXi4iYQga1UDA8CI4LT2AQOHwPhCNvY2wwMp
gHLHlg+31B0VQFIlUkWNH4Bx/dvLeEmuA5rHdm7vf9ntHUsBYkmm41eMGPB6
aNu12Bf/sIxpwsq5KNHmDSewF59fzW+gFA7kQbX7xrKvIlCHn3wwbO/COSU3
SIAXHAaBjbV4ZdEL0DbJUGXlQqnafy64kyHslBr6NCghThhJkjr3CCDFVBpo
cGH1g+ZAbmKLU7NYSnLHYYLvI9DyOeeF7Ljp9nCv8nEiwVINBIFl+XQCNSXF
Nxp2XkoJNnBnbXO0s5A0wV4GwHBuMX1enMLluzpYJVjvcr4sShLBMc87Viq1
/a+5rkP6wAQvUw/8oohEg3T+FMsEnjyO


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sX35fYY0/vnxSNfmzF3/e0y6dQ1yXMJr/i7JIRLbChi/hHK7lHuVRy5hkUhF
iiCeUBWVSsbrkOTk7phqk26TaXPEa/YRTFxCfb7TPDnPanbmFYx/ZeWr9NkO
FP0Oodau1fPbCYIBkd4X3n14MQZmEAH4C06BXnr9bIizj8d0070=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
c6N+8aDzccXK1jQlqR934VQEB0mSi52xmDGiPHDdOF4buJUfx9OnfPzoQoy/
FB6Uom1EaXCuI3VAvq1u9VPJKJEfPxL/16DXy/kp9zVbLojg4vHaOunkxP4p
nizSG+aE/8EC+71gyYxT6IR4dFUe8ZSL24t2eI2P/pGVYJxhPQU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3184)
`pragma protect data_block
toQDDfhNf5TGWc0GJh9PU6JYDkp+LdFjN4JjwOU7V4zYAtb4I0GS+/qua/Bn
ux6sGDf+IRVk0d4YuFDEChWf4cvR68OEOVI9VpKXIe3HWXtBE58Ii4Vvp3lf
oX5j6XPHR2otU1ok5ULFv2wcBe3Xgzvt1qQTB8NLQLkHK6WVpYQJtMNgsYW3
4vfsShnVofL1rHCw/F6988/so9pvLPlQp217Qr1JfSa1/VBcH9oYul192ndU
m7lzAU7EdKMDGUmnoO/7Bc2fqZaGAk1cE4Fszdbr2jX49MOg/oYF5cnxVT6U
Y36+c3XEsD+cwP4Ri4bRj5UTYFhT5qeB1XKSpDcTMAFJ9BSey5jiodWTS0IU
EZdh3KVqU8BSXu2whCZuV8IlZ5reaG54dFgIlvINgdanxSyra2nG/zHchGjP
hJ0jNQwXKUHQ6GT2929yonnVVWcX2bxoVWICvdCricJ4mllHGCXJd4Y+wU8F
+ZCBOmG0l4e+4yL2rBN4Gmuaw2R/znTBNXYBUMdunJ3bMmHDblP/DoI1Sn9Q
KvsB/1LAZtZKoGPNPyrrMMjOZunGohvF1Uai1798lupDxY37MFEZ6XtgNIgh
xeBXh/t4GR/yHOtfPrDz7b9RGMmTVvNPqZnU8ABbgU+TqPKLcfZhPPh1HPe1
LPKWlnzv84WMdn406Rq+9gSNwEbJVP1PSJyXyBjnke5/VRTQKyxsUkvWiVG8
yNn9DQpC/WuMRdlU+kgF2VGvre/Xso7YodpFChJquIhPzJxnx0Gh1eL5595t
tdIO5Q/1FycUnoAe4dhpWPIOf7IDWCbcKv8Om1YKzd55yCOGfkgHsaHM+RkL
ZlzMS9QeHWICLlnLccEjrBAJYmD83ZlUKmk/g9Fq2LxeK3RIO4N6E5wVq1EX
0gY74SMlhYxye/ZJwwLH81/GATLIGC33I5sgBGPyhmpzH4mtlxNRWorBIh5j
ogfJqE+A5EAF+KQzhcywWWoYfUwZyGuZfqD5S/KsiApoEfkRAa5o4pZlwOPc
Q6FcUXQ0Vaah1y3o4iSuCHUQZ5y2PxGmogQbL1PTFeY9ns297fsWFLxZ3nP9
NTZKQi96TaOMiR7L9oxfpwfP86e4vCFXudoI645AZe6dfCDLbEixRhwWEKdQ
d6hubTESmji6VI65yZyRmJmlfqlW3wnnzgOnu50Sz4eAzN6deXcwTsbIsY1z
AO1e2VPdgHkuG1EuloGQRjVZgVwNP/pI0W4EdrlXDUgWu7N2VkVkSTSuFeVF
wlaE94jzMl/1iniSLiaxVnKtiFQ0tM1ADIYjAAXfSUMBDBjwdBrHCfTkhM5Z
q/M5gNplBxrQnR+k4zVC7MF0NqJ9fWEO9NU4W25Q2G6NhX+KQgaARX5jrZRC
hZbrZWBONvYLiX9jxg3tj7MAw4ej08AKPEZiGYV7N5t3dTKersNvSx8VSk5B
juvs7GqWK3NCeXtgogg5y8CbP2MR86gdSOc2fgirRk7DI0ZdKZ2dqpdUnNEw
yhRFYVc7+4jk4zXW8NmcHrYl0WrYUYL8jDl+rxiP8udzuudu11ES1ZGYNaZJ
WGlz01T99Vl1JQmVp3WSql1jb06I4fZjTHvojw69evp9fx+VHWmrh7PjrssW
nKM5+UoR/M+MXdO5DY2K5SskYCg+Ba8WVUMYXSXwfrenRfWARoDf7NwC5xbs
Sdp0m8EvGXFQNMYXmw3dCqKcHKReC3SDvRU0tXhwb7z5ga3fNnZg1We+bI7Y
9HosBYt9HoZqW4/4aYMBA0Mt78645Jzi2KU6gDNOZSlPK6LLwywDO4h2rd9T
TNQKFG3Hz0xTFIVK4p/XoLfEaY30e0OsEtNp/HXTCo/H2XgtgB7yRuQuCfUS
NSDFx5aNCNUZeZ1sjshBemXslP24AWJTj4Wdf9XT/qQoVvkMGZ1dfnpzQ1cZ
2HUS6E+LnGTHzm2gGmrxlqdHY60LQ/nLNms9GsADLGra+YjdLzKA6tBkaKpg
h4L2CUu0Km4+W2JBOZxrg2As18PpkgDk2SXGvCHkyiosYZUoSCigW8KK2S1s
ZcJx+QJkYARlidF8EEN/oq3xTJUGAOnj09GQLxFqbreokeEGx3S1gEF45uLp
VNJh0ZJh2rGgSPpDmD7A+DpfC245DK1KUlnGQ5mDFkilvYFaH6hAR5cvfTBz
Q1+i7xEVZwKDlvjOUyNWfW5meZ0uWpnDtX6Inpy2k3/3cAEdrADh7REWmLJE
EyzfYLwSqW2n0D05C+iLwgJPOsy5E0SYpUaG58P7Ysy4GvzCtAvVZOH6SllM
kPqd7gGjvO6qibdD2PFkqG3btfs6WpLSe9SehsWLhXk68RbWfWWe/vFBVJNZ
3k2Qfsp71qIQn0R0V9m7S+i3GIN4MD1/QCTrGa0UvDEzfgCrnvw1vt60Oprl
5EHl7/tEt0qL9E1pY+ZBkQqznt2vYJgNTFVPTYajm3mbZXoZvhA1Kh4WuEcE
aQ4zi1sB15wAWsL7wy9VBm+RNWWIeYKL6xW9GcH1vhnngX/ib3hIKK6iR2C9
psr4iA4ioBIxf+HGBAAiX40yNZT0liMs7KvtqEkbZUnQvFvF831VXKchZVi2
w4pkCBlBn1x0jKa0u8vppZnueo0LCSDAfL7/MQyuJacTugg8zsSJoGEugwqr
t4DS/AS/K52qEgUGFgeXvWGqMVO+dSyFQpuSG3rAzpFDxc4ZF/3edxvm90un
ISAg0Vpdo8oP/IYUSpPN1+ReUP771hZYhR6bZz2ZJnPJs8uN/LDRb8h2tZFO
Lhk6MTxpn9A4MLwop/lATVxFIEKwcB3hLhXgkGBgLn8mONQkCHz67W6smgY7
SWNAN7YRYCHiIy5B79sE6FJC1icS6D988MCrAnUaSwNJ688NiMZOFwhvlnde
BomOtTdLD5fbuwxsAIc7k8ZKJmekZU58/cHTVhCMmXhKWH5/YeghZXc5jWnb
TRkWpFlcw9BUUCvjNkVa4TT9UEFIu8IJVQ7mWkq89mLiY99lshgcARhyGKT0
11sgldpiEGMBIXE+ahvR5xKFd5sErLDDwOxXdYEtulAQe6zAKhtVkrE5mzTq
JD7RDOp9uYvwMLIXLbD1ONMtpFxSU3TJ4//QEclYeUva6+n4peXu3RlZj0qa
uPmOiMN2sTCYZcYGekH46v+XK2+6B8TdCXANXXwpdW0UIxPb1nC3UJasWc6d
YIchnNY7y5/lsaIgVqfyoFRVJGHHECOLZ68FquZjzgyKvkS+MifSFJZ/Ly/M
t0289EdeWsq6zYiPfgZOUFO+msC/lihsYSYo3A85j7lV7WQPVKpW35kLaszg
AIE0VtTng9ERN8ZkrCfHoSpvioYFn00MNSi5QX7GBS6FQL+5Zqlo0g3FRCs0
CRhAjxZdOR4cJU3efISG9EpdANME3CDzYjVouHob19eAzSGVnWz2xngX8XXj
foKhtSrI0Sj99/iWV5DDf3SdvMKKezoE5BWckzpwsPHcrWOz51+NbzjuyqhT
g3mEJQRxW5vCFhE9JleHt204BPhAOrzrDHFq45l9PXIhaeyEoXXUAwb3+Q2H
p90G41Ye2bdXk6En/jNZi3DM5eLUjact1YVkm4lP8HyQQ0oTB+DRqNuZywJT
O3WxlAk8YB1N/JimMUcQhTytYu4ohlM7RicNOuYvvSmArVVfT3ToU7bUDf7n
le2DXPLTNNDBp1E/El+2mb/i4KTbHbQePC1z/aq7LulY38C/MzZNkPsXScgA
iJWw6sGC6eLsBLj1/s4vlPAcOCfGzRWkIGnaCNOq3L5ml2MCuPn3HhflBDlQ
VeUlDMmVIvKHdCw2LnjsgdS2Q3R0jNIZ2EKo716xGc7tffQzs3FxkSoKqRBo
iRigIPEKFGxTFoaaFK6bxTkw7UTqKuqi7OixgkvQopDkgmC88GD4hnK8pGZG
9SOqhUzgRRQ5ZkDXL+w5T0Cc/I0nbuFO8V2LI5JTOFvBcBVjGYwdZpwJOcUx
H8ewf81ISb1lDzMsnXWZrwZacZgol9fr+S9r4HLxWkdQPKn8eV3fSklq8po7
7/93w/PvOMpKDydthUd+9Slnxua4zX3R2BJu7tVIiQIEg5SkBkFQYP+tlWnt
2EVnIOZhp6MpidHl7C8cjgiamDThsRRhBqH0CQXJhrBGdeJyKESsJgR/JF8Z
IQ4U4LE0BhRT9DEKr8+p0netl6fhA2eCk4UsrK6ByHO9RuBKK8w+gmzwkQlE
DAECFqhBAjzRSNL4A88C3GTCy/JSkCnNx/b34Xq+CPS0FQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "lK4MM9NDeLrdcSiRM+VIuNgpOLUAzWAt6nzBJ3Vw5tvBogzjtStM5gMJjD6PMmMyupOFzYouKIpJuOZh/11WnQBMmqEc6gvbtnHqfGmxFaxYyOv1rddc1B279ac1WEgUgi2BHG6DRj+tHk4+Vv2VvppW/Z9gUZ9e40aCxOYZZHwEVb/SJ8ximgD4Fihl81LOgt6U1JRoR0S/yAHMZXIkaoJ6FVEBkPAD3J3ew7MX9EyFzSOT4EA6RZvsJltvssSDItrXYXAoFKzgRQeSM0Yf1WqqG/a2yRt4aSBkpsO0vsisnQ/fmInSHlFF/wq52TrIXCUQG2d/PbuW+TY6sdsOvD9v9bJtgv71fD2Q6WZ+S2xOr9xeZ8H+NfuZdWyG8Pybe74yPh10LOgBFSSu5shzFCyy8wTK3T6djQ0wYSTBG/WxjG15qTZ5DDuhwzNJZeS4Bt77+DBqmZzLsCsE7950nWNpRD2m9cgu1sZq/fsleUsqqIQrnRq4awrHAK3ZQczIwUK3sOypPY+/sbSurgJkvqZyO9ASuKMbKgMXcT3ZnD46k+DZyqmIkOEqciAuMpBLWzgTENmecfSK2XY2mOZaMEuHlkwkitBprbaaBN6pi0YAiBp4UxNL/3qgel+iCgzlRShJDYyIB/yW82+Myi5EBoITVEPT+fVLTfIGJR61xQkwiFLQUkpvf6mQ37TQvCD98JHAhwZw+BrFlTJDkGaV9BfTw2FOdNiwyTPT2b7DWhhhoUKSvGgiii0t9yK3h2OivQiFnr8XEXbl2LNkVmpyMew6iMGbP3Zii/ayk5tkYqATz8uvPK/KdPL71wyHTFWuVZErAov/agS8QPxTeouBp6QzGiaYC0aPm2XY2Imge4MHVaYgIbyAHAgCvRrIUUwoVUBr+y8KiM5JksPq9Umk/CWTW7GJ8GiC48lDFL9zw9ejyMQELz54535q0utjfigmRFbWjEk6I+exAKw6gx6JLdEb2+mGI+XxB3zlzerp//3cDvhnJb0JlzWvV/vOp+tb"
`endif