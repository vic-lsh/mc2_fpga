// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mymf2OrOV2qkTFCIqliXMHe6baieXeaxuZsF7Oz2gQeFeCVd7wnxqZRAE/1Y
K/5vFrGYHH+GVH7ePVCFtowrMCqbqYLWN6/hD3XaGVcYS/37Mv3NYbCOiVfY
GYNl5gOlqdMEt5oO7JXoYjbat2IOz+8NqiqgPYLSf8FmIxxWuOiy+1n6IRcQ
H/nQEswoKyLu4mygdec4gClcltURfpK6e8cPxWBdn5S6cwtVIasIkOlUUcWX
3iMR9f9ZvRrzzG/O8Cm4aNwNOwZepMHKuoIIZLf7ue67U9e4asiT8GHhnmTF
Kqk4J1zhBmFOjaT4hCQ8bmcJEqihvZRA3VzW/2yKjg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ffqH41W9D+czMv9/Lu/r6w/3YfrtdypyqIi7XZlvNiBES0MNw+fcsxEL9PaZ
w2thnzI0u7v06vEjMRN25daih4ockIHe0o2LCbFTQof0Zk8saD7FBmFKKqN6
MEIoEDXj637cUClgugypdAfyOgAr3q8AjJm295uIZ6o711KARzZoQVq7Cb/T
YrwOCfNwV991SQSTu+mcAH4v6G+jk++cgi46b5zUj/Qs66c5F7K9zYR7CyLE
e5yXxKtuhmTQxYnxeujXVSWaaijYlr+sdcij751NKnWfhFI8DVjLeJmkSZSQ
98CIauXYv/l4Yr3CRDcG/GpGQgwklikgiVNRfhHKnQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XNinpY2xbs+fDue/EbU9BEwkJd3hbHafni7/9LUB0y2DewG/wkZWBkNS6XyT
5JURzZTxJPoXClCqwWCdc7PiP+vjCMEhLf2ccQNmleoNa7klE2id5+tukzXB
C06XnlZN66+db0YwIk4LP0Mzr8w0DfvaYWDrwQBUZzTZHMGqqhKc5nQ8u+Yg
O4nHwjiB3QGg+x2J/7X1kjgqMsZEng1CwKt/CgvSDQZHs2iP9NVqDWDddHX4
8FF4tL8FZdlHUPbSwx7adjyLOQQkYaVjs5MNAnU5T6JN4skyVI1hQGMXN/5u
XPAbVMGx1iF1riUvp+YNi2jms6jTRxktmG+sX0mckA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
laONAI3c84sCB1ZNM+4QKzxKx4syll8jDMEQtgyMcgAr/5+ZHYKUPu4m9pAm
yiFEnGbDejqrG20KKQtpkQr0T9lOzHENEDlT2v5m0gGW+lI8ugsUg32Gi93j
9Z3Ir4v12/7drIdkXvSUCKc0l5BmtwDn+UzGUdgodxcIDOgcsmR/xaG52kXU
5iPpxfZSjZ2CQgnHSCKFHlZwQay1B4SXHmBMUsz9zxSNOnJW+zcB+Jpy1NZr
KxGvWYJ24xA3B66xNKbN7G6UGc1Hy4+G6d3g3qnUewvBMWGxDzoF2vk4Oy9T
MIvHuxwopAAhSkeu6JwpjsV5u3Ml1NDdDVLIBdKCug==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hJ8Ux4wf6za/fx94MOuDqhOZxJLcqLzK+Dxl5cqKdSP8WVx0Jqc4zUGQ2Qga
NKpIJcFImNzZ5GuH5PgXnRIn/25F/StJ/22anEzl7wYE6nFMXsIduh8gDmu5
RhEgvffrUgEeKda7VTpCMAVZAokv4ht5H+DHey3NsXzx4FGh0VQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pbVYCrlnxrZyCvgRDUh1g7IzL1vS0SPdVxA0uqsf1pRlo4HnbWPWtTrVoCU9
nWeXNfLOStuRB6R3ERnGc1DUgieRl+t2yvfulETRUmPecvK5TNSKSAGalrUQ
1xtYAXk1xPu0DShCiupsFXjhy2FxfpQFMPp37RcWnLGHSCkA7QEnrIRwLlHA
q8DX3bludJ7qCcETZH/YHqBVu2qk/U5BKwE74CsYr1m6plcYesM+EB0pwaJW
JaDVM7QrxGkoi/No/fcrmH2AU8VOc4m8UhyPrXKgVNGvMQ0TND+cXEVlh2nI
3uAmyaWX+mTc1Pal4LMS2ybFXQYpqL+WpOK6807BfY0EuDStFlWgoTDm4LCw
Kunss34VTHRFTHMwtSX/rX4s3QB1FiKh10cD3GgraHp7YTafGGSIbJe1Pg2h
DiQjGck/nRIhJMc6fCHE2IRJFSN7ucDIOqFMb79aPny5RlKCAGcwGQbYSvy5
UxUD9up2jMlcAj0XbcwUg0saxr+CNArM


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GrG3ng+vXLdlW9urm53X4Y13VLcyTBfNVCTWpv73VKRjtIefvvbR/Qtmz+c6
TM5/P1me1B14UAqhqtozrlWIqHYmEnV16qJGNYTLsgyFhfz0+Ui/K9JT9NOu
EfHlFmNohFLg9i/Gv965wx2oiy1zkwAoOUNLMkHzxQsb6aABCDs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CzW46q+lkMlTc94UsbEicLQciJHLfY25iV4DVhKeVZp3ZuhraMDRiBlk/jLo
odn40/NQ0Krh5B0E1sf0EL4NEBkkzj2U84vp92ztOvhFoi7NA5P5YIqE37YA
NBzFWT4h5EOf/FsLYoY6Ffife4o27BHkTDY9X7w/9aNZhFqFOOk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10336)
`pragma protect data_block
QDu+UAeMdLyJ1ptleCI8/nKUVfqLi9NRdlxGIYuXOdiVYeJquDFdXDXb7+mn
ErVNFZAsnkIrUfBxtQGzQ/i+HYTvtY4aUozNeDD/5X2SD4kUL2alDOqEDVJw
SXbThuiHpZxsGlIadi8fX4FhY5szBq+07S88Six99ZxnkW/EWOn3Vuc6CKtY
u8tuGH/a8+TJEWmbDMvdq1UVYmFoJErL+0OkrtZWWAAJyMPnSgKo6OEOE278
bidjiR4wSTAR/u4Dfap7Tvi8ojA0Jqq1D9s3dbGQtSALm9WGZiGzIl6x+z9i
usGMTpVnZXWKI09yDBEXgcPXxVKCMdL7k8aRNpmeCKBbHE13H6HA1dUTURAC
riTfiXfSptJTW1uxqpayJUbVUR/rSap1W8Cz+iRmh1JQoKVUZxrHR2Plsg8X
zgBcEN4TNGJTNHVjrabej55OUBYJ17Fsyg7YAOKqDoBeTAA7I/wtT4Gk+UgM
M1pQNIAifKS6IJVZy/vKVNo+RD+SoMjs3WpaENx4z4h0FKBFjBsKXJjuVfe5
XdS8mlAyoa7E0ZA+zdxEJ38iBuPw/Qmxyh7lgLuLhPdOQf3sCNrrTiQoRNmd
6Sau2m2+/P4vcvpYNwuc9nJQwRFuqxGBCzBC8P7yeO3n+Cfc8EJssKTwOtrh
mq5NGQ8TD2KYD+Nmjeom17L44kGQ7w7cP7ZdpOp1/UdRY68HwQhBG3flGjKl
vUAlqALpw/QDTNSMxkiymiZq3M/G6H+/pgOEzpGMZDDKhmu+ZhTzw5oVSuVz
4IgVpHvz6OMD6JUlK7Tln4cASoBsXX0wNqlNEEIaGK+DBAWHCUcVbZY5LYvK
s58J9QtEDj2IJ3NRMR02pIuuL8d4W/8+OVznxBRErZW/Nl5PEtfSoOSbus+u
ZjGVSXctdaWfyGd+B9/LWojAYQCpun3diPwr2PyaOSW62esWn4+da1RPfxRt
IHRFkkvoJzPlGOv9vUNUWrQGlTAoFV8dq24H8451optNmZT9H7F2Yp+E1deS
EcOrwycua4eQtJJ4rezDReuRrYS4aEZHx7cu6E21xMDRk6xj5kFxZ0BDxFFE
+hkCWzFYXKV0IkJQ1+Aad0hgZ0CqQlIXMscwNJ+a+uRVjDh3ZabWje/AkKso
4wdvRMhzBH5qcp1MI9vLfX0RuCfY5a/9kzT+C60zJGWobQ99JwD7E/EFm7BW
UN1AP3DLTlNq/cJMjU9kiFfqv+tiQNfBcgFgEoEDmrLYJ7gHsBzEA5BebahW
rdEACvn5B2A+kNQvQL0Mm3FydsIHcRxjmSLnLfo9y2YxSUPyIIQpeHTK7xsi
Syv30UJ7r3Arfe0ag9SlgZqzznAcVsfNfEmZz3dj7yxkurXh7VtTW7GUm57Z
FZSgm0Pc7EnkhqjPWBPFwXs+QdN9p9CHAlA8a6R2kBpcf/f8xahwQBk5+YW2
cYygQX6woTVBs98CqDxRGNEAkaxjwxYPu47/Z7hsFTqnmhTvkGOtrO+JRi/5
DtiouGcJ4dcx7EzuTwD8JcjNbRDwkV20pfD9dnhmkV3WKSwNFHVIJ1oY8H2m
rXp8wzvl8Olkygd6MZqJYjo/Q0h7Y1jG3vJjjJkAXbx47gQMit8Uc00//Sw5
NN9OfHNILadtkCDRMcWkedBEF0/3VcQ3w5WTCM9QCUDA1uCY98VZ2JbOylEN
V/4hmBHUe45YNfB66NteYzmAFcApF9YQ3E9Aa8L+flVT1kFGvU3JK2nYo+Gq
B1ZLiHj64JdQhYo3VcZNZEcPA9OYNXXulITod7mewMMdnsDLBSvGfcD5QSLj
pn8wzfFwQPi5MqIpvoFP2X3LYueCaZl2XGlq8vUEas99D4g+SPPqGu6So+Fr
dBZ6IXA4PUhNh12NyzsZ0072sim/WugUb8LhvlLIwmL7xShbgfBZt00uxfHb
zVCjgoOqvjttmY1mrChPW9KnxreoeZDI//q0Bv/e5osJn655l3q0eGAd632v
susddVkHdnNwbNzEPXSdvqwtqS1KwpblhKmhgxwJ3HHeWkREF6sw/pmPaciz
ZVFmF0c8OynnCy81fK+uQtYo6YNgziKtdb26yrpAvVt7uSlporDCQYTABr9e
0fvd/2peGOBur/kg+GtBllCH7UOoLjcmOeXmP++kZuLDk03unbOVwB4lFuVd
Ip9KCwgqYCWltS1rucUrdwblDGzOUGvkiWtuo7oi6HLAYKSn4l1H3fWTntIf
RkaFPOZ0XoIWt33BxCyJQJrLqluJKl3Tfp3eWiBM4Iu3D80bwrIcfGAEIMDF
ur7ww+lw5ojnEmv5sAn7dOsxhxP8xdvsDOSqj30Mse8JLGBL53RMaFitlUqH
74H7H6D3P08h2H3osArVXhg2MFP8AFx9/zESNkhtupZIzqS2RV9q9J08lZro
uItV7A0J0WqYHRZR/zkJnO0Qh1BPyt0MjbWlPk0fvzSoEyFqHQwUZIHzqwG+
j8sTaue3wITfbqvo6ay2Rmcxdjntycu8IIXMtpclsBfVyzsUYi/sag9Vg5tR
bhC8J0abSpyiqXv7lCQBAFrwqPzlZCjwfRd/+4Fwr/1m+WZD9r/klgQ3QIk5
bIXfFhvbJEx8BvysK0eUXUi5/aWrvt030F0Lir9kIIiw3/bse8nLFZUIWCGk
w4gdir3V5UCv4VrfRPOOwK+LWC0JmVXsf2OJVbTb4F106QpjVHqTuejrOJw6
3KHorXvbZPl7zikCejcIQnAJakWs8avCDiTW4bz1XyolfKJ50Au9Z1Wt8Vf3
g8buGHIEfWl5lDNPX6NMEkuQxJ9955I5vjbgWTBODOzZSXzPzuWduCMxjxNr
49Cie4rqzmU25S9C88rBuugJIWtmjzrd9tLe8d9VPyaWnSZt4Lt5g1t3qFPq
e9HLnCrOD3T2ciXFALZzupCw0iz+IFA8PoNpDGo2z8+yuwBArc1Syq2ZUctT
27H4p4ptQ7aW/P6DRNM66oQxXSDEavjzsieqhRVvNXZxs13lVCBKyeABEOi8
57JZxItZ35eZd7pYnk3RzIu82dS7FA2aRFhYBVd+b6wb5WjSpnx3zWdHqqVU
fpzDPcsqhHBpl4xdvfJjUrA3g6sNHM/GyMEddrXWpqXzCSCJOqDcrqKpbYAe
Z5vj1G8qTCGtN5dRzLOvtsmTYTfmx4hz3JU29GAr0eyMACpzvJYp8KcLqnKn
PjUxZIkX4ljHj43Hd6kpam51yXkm5tdBCH7E9s0AhuDgsmC4IPhS41n+cMwv
sbyQRVDch8KSOtIWoEc27kLLRk0bTYVYLdl1kROabw8xO/J1HsgELN1v5162
2kBLeaGmmp+iRSSnsgg0kd7vJIE3+IAF2uyT+1HglbUjxDvIbbSas7rUfapE
mTaLz3smGuJG4DMm4Qklaz7LxknnL0d7KlvY8tkXFiHkMO9BS5Lt2zqDHFm8
C4kcOLk23fRkAR5XPiJtluYyI2JVMhpUIra65OYUQqgZJeUFSAk85I2A7XFM
SDO0koc/fqh4uvyJz73/EyMwuWniwiOzejDVEA574H+wocCZWVK1itIwpbWP
f/FTmMg0/tDHVQXJPMLDcW9f9pfRtJOnbBFEumL7yeWIxCmubfd8h9qcS3nW
iEBP1zA6UshhGHTQqJF+CXpHHuazf5kilrInmFvoVNakMABLFbCnKiYdZZzw
hkNAtWcG1U9+x0hCVhcnisiSD+bqdECkBLlKNCq/lUjabsmwqdfz6N6kHUY1
7MScrdSaucW6/LdJ9L2ucmGQNnrlmp4aILyz8BgALJ6sVIH6n1OLDRX+Oniz
904Pkh0CXpFwtEMPAOg283RPupfgPNSSGCumgJf3jFdDPRLPMY6pOIU8PefY
R50Boh91lrNoDsLbmk3lqQtF7S4tYFzgjdxZSlDeLM5U8gXj56OE83oJyf7w
bzHaApjYSQMUNGu8bty6iFSkzN59wyv1GDYHr/8CZqz1qWG9G5GzBXPG/Vq3
Mi0Xh3w4udAF2kX4YdOYrfefs6SrUZOCH4VSAOeEeImV42uKGYp2e/lPFQaX
E7ti10LeElirr4CcZfxlGF/NSjDYFdQoeR+2K05al+K34BNlIYG1mqAUeVEi
ri4NpHQtCbAOcYNKcx/3a0wiYO/myWoogU+R7bLB9EPWbqkpPx+0+lYgVsFh
B4tNn6eWriEfefPNGoJANR4fqHF6EstOXK9zqed1H9CEO+H21Apu+BGhZhOz
l8lCSlj6OppduDmUOWr3ZniTHNMac4ZBR3+ewXhq80049ZkHbNlKyIh8BBQu
UsIj4sThAzS8faUhyqk8Sf99d8bd5Mdd1cQik2eUapwz2JqvQwJbuJZ5TCbV
MWAm9R7hQAS95FlVk4pEfw3r5uK7r+gW99Rst6ihxFnNfxDNTTVSNrfeYyq3
kZGQilvKjjT08R03aQRay0WmzqFBV9r/lX7jWe9NqD44LXxQImIipJKAxVi2
25YiZfD5PVvcrLOV7i6XpRy1quPDYVw2toKbbbhv26GOdc9qgJCcdx9fFCrW
8OqFGowKjzuIGhQcVfmaIj63UoZrimRzRZHyKmKfUy9TrAeerpamWyll+uU6
i8bgOmxr3lfCIh3vOB9/P3SM2ySDrvR1gB4hl9tEEV1DRtws7jOC6+C+2DTN
o8KWxxG5kXruyogoAst8lU6moMrTlwlivoqlrFIMujFx9Xpk8nUxPbLY6Wvb
Gfo5yoebY0XGAsR3NX4EFCWYJ3ZmK938pYnczGD/534/nGPgj3kGsuZ/5k6u
aog9b/x8cvawfCO5qBrgb23u2ZlbffsdRUeinCauKRR+wZHFJBnFssJa+Tov
1kRoKuUt+lLNJoAM8Z9ybzjDBStvKzZ2ISTqcZwzUVQ8eYyitnhQtPW7zxU5
wr75RAXVrnHxi8xEDsQM0xl7jQ8l8amiuMK9jyS5U0pd0CExBE3LVLFBwZBh
9D6NkOkstftW/zL/MkE3d5JBbspHAB1AtbNeu56k0s7izWrhzYpK52aqCXAj
NaBIRk8TRt2Wu74f4zQQFtze2gYNv5Gn/qsm5EHUb2fAoy37Mvb4KdbfSn/W
31Lg3G1SZhVbYzfsZ+Kv3u4T/Imu3SOk+FUKSb37j7lPFjXHwtRcZ3nTbglO
NJaZR43c3f4cfvrrIno8ENwegxYJxULxasuj0hZ6Jvc4zrZ3PNB/Fzor/U7X
/RpN9t4f1io6ahKQvWPKH3136i1M5ANwX3FW9YZXceIW0NeLHVWX+NnAyRND
oPQ7ObVFKFiG/Z+Q2O0PSotqHkX95wWxyR261/w62/J5z9/j87/QvTrYQT/0
nHYneEveu02ZdiyTFmkO60MyAJ/u4rl1s+JKoY7i4HF7hqjBpGtQkGl5gNTN
QYPX55q8wtGlcZvELz3JWJEnz4OOcjCecJw6x2FX+a6rBJMunvNrCPFFCgNn
fxMHiewqCYBQOn+Fh8T+ZE6fkpkum3IvWPtC0+pzRyenaaA3UaMPykdztUxW
iBbmwXDE0JQ1uR6Nl5oot33ms4aaAWyTJR2sTunfUHiYZl3+XqwPw3pyN2Sa
EL2LnQR1ja4QHEACPQA2Q/ga3lbKzoMbsNYq3QTWTvld9tI1A7uaK/gEMpz9
/JcGVyO8tWqc1Bhv08cqF8agNuLQx68nOZcTVPKq2nolK2IhwxaNKc1o8Nkj
kSvr+LJIHYiG/owTkFn5RIUqoGFKgIkV13RtOJVStVaH9ODCm34LxBpWK4gB
/KknIUkr2Dhap2XJbGBTIeJ6/XcWHOHYg3R6waZPhu+yscHxZTKQlXCXayjr
Muv2I/O/gPXbahrsym0tZREtvUeRNtlJl5jTfHIX/BFv1D78cn54tUhS6+9h
FatU51D1S1g6xyITRVxbiEe1OaJYc9AEp1zkkdlCzn+YzRiWm1pGSmCMadCC
zHcxXCdK2PSsAv7RJXac6jGWQ0stVWQsELjmX1lwUbbYgGrOZ/rF8qyuc0sM
YPu09FjSfcgysMMyrNaImUma9K3Sz6qdnRIk4MklIob2YA8Y/6YJoDL6BeVG
Frrk7fFitfj65jQurZsWx4mefQFePXBPCUFDZ4xj7aKCthUNqQtyHgQTENvv
e4wLx70lCdBZjXeuWjkmgOcLPGUUoP483FYAQOjrAYk/cA7q9XC2YCGLfrOP
GIKq7V16kyFXOueKQgiBXd4T0YJQ0XKIcnP8/s43AYzG2k3UJx4GpMiCdlo+
WDJ2sQf5BP2wZy6WW5kmbNovVC06SXK+jJkdKgfUW5IsarcQgsdu9jZ0jmHm
+mx5RjgckZN3uHNlFByqRDaVoiiAKZwWCREcHyTwHHRAWfAfBXxl6eb/gK4X
ap+2dSH2qK4f8k9iPeMBcUzKnE9wd7wJX6Tt/pTBI+JDbk3XKUQn5SjbyedT
mIONajCe0XO6To/vxClbZ1XXub4FiqXBsCmCPrJYUtzuAkDdOxzzcY78rjel
DkvkxtGZVFQOEORd5IG6SZaU4YAFY5bpuVCGQPQ2x+4CIQNtcKoqZ02oWm8K
hWbI8EsvHAFU1CKTTyGw4SFvuaOld1BtElZ0zgWFNUI5dPC9PghGE5+Sp7FS
+PxIqlalgdNR/rcDbBOLfqRkLR+kLwz+7DSvixPHcAjvKJjSMI5LS9h8SsdS
Y/ITvMYizTh5MxjPWRblBhw9Lw+GR9QfB354ZMm724KXasNFJBjqnrrMHjGh
i3LqQlBQEuSzpZdJi0Tnt3xBcMPrWerQ2dGkIogGNN7dNIT+hLFZ3EALPMFb
CdiVNkdJT/YmifCQHPNNRXzJO0nR3de8/LH0QDv0A7oWlKxhWbE/XsyvGlde
QKu22toAVHVsA9uFx3kkH+lhs0Pzh1QNXwmIODUb3YnyGfPNYwVZ/6tLhmqH
6ceMCD/xKBde35GmolGcevHwHJyglMIjTVlix6EMsXUEB9uPtAY1C/ziGL+r
c+Pp3roeA4SC2gGqaUVU7cUvQhkEWg2UOmXAWE1ytyqsJyAWr9eVaDhKweM1
E5een1X2Nl73VU755ns2C7WzwN87krsKCQ2GTfkP3CYiHfw6C7WbGsgued0D
4NUftVyI3FfvnYv+zlY8mOw0/klXEpC27sJ5MGoEMXQKPjbFYphBV87Yfjva
CmwgwT1fSrmZJDMcFvnrxPikeFcgnVpnje2VYCCLFwsfCcy998ioydrej7bJ
V1JISqxAt84aGAeHpN2UPQfAKTUgaXJcWnX34cRHL9rx7ambodhQErgpcwp4
CBPYb9XH2TDtT8L2JlNpEM3rGSCb7o5YcsN9tEkZOpULI1WSPjg/Nls53kBS
z+dyNEGSYlcHPljCRz7mbIq+Q18jv7hvuFkVziEgwYosdFkL4Sfpsgt4l6G5
1Fn0e5Xo2RYxq7dL787knnpNn6n/228ZHx2jM160vr8x0Wd5LUPI78ifbsUk
myLhWdULfyJTqJeq4h2lxpQ7CeXSwS+OizkNAOAOsFnaaKvEnCmp6EG1c+AX
B82yyG2vlTZU8pbLlqjjT41DGh9DV+XaWFvdjrfV0yTnrr/q/cNk6N/UnaSp
Hn2q8Afu5gea9rjiNEbKxpluknvYBHeZsi5+D6aMsZpfLJyKZOw1DTwSEYpn
hpRYDKA3lZOVsfutZUYzdR9k/AHfy3NfgSTKYJRIBIvz7T8Zb2LJtQ4pwfwa
ZpkUJjHHymdJzWn19GB+Luijm0/PL7n/3k2K1+PKTfOv4p4DZWKGo2Oq/dvo
ZGVxQZUdXfn+9pUXOpLB/2Uf6EbfBZ717rNNfvDFgURMocPJTdV2xoxnF0zV
uvr8xMJff05N0JeK1qZyrA8VbY8dgniN/5fZiIOcr0o7EA3xSGQ6TGF4EEcb
6P2/O0tnTyxcFQ6F/d5QBu6xyX4P9zfS4UaEN5I+2FmkouR2w140y6owLwau
HfTpwoBJfYZ5Jc1rId+nqfMm4EmMlyO6UrZxpVhAGs6IptnDfr9F+pndn6ID
f8SUvRgaqE/2S4KK98a4zXOUblpXHmuMgwZmh7I21uL8fkxeA/ZbJ9pTRW9t
TP8ZTF3X3uhF0YYktd5jdr/bpwZezF+yAJ/YXXsl5AfNAH9lKrHXn5KyXmPd
ja3SrR+XdTr8TD6JXjKxtdf2kmRcji9JOxktnMFmq8if9DPnRsggT3moNCT+
17P10W7nt/Wj/P7iapxVndPUoKQCFDowfkHpFqqkVIydeY3hmDoak0IcTYqZ
LPA7u5TZBsl6gzkGXoCYwJOD3/czIE4dZN9spj7WBn2qfrZtu/SaVxbBflZy
nSTWS5PsFrm9VvO5EhCXrMtrOCPotyo/GWPr+erlekENht4IrSTVGiE/wjGX
/RJvwcNf2PWl+XsCWW3hcZOXqz8HuAqnot/WtzREAznGQTXQDLE0tqj7qlN7
buLwt49uyjq/MvaVOS/xGCwHmJetuQ0NxEGFhTZt8GmOQtiUz55A3jTpJaZe
FnNJZrmc376bRsTBxb2IcGCsZ5iKIGLxL7c4s5taoBSIxvT4Ox40yDUd0ldE
CpgCyyaK+TTmHxkSxBTdJc60GG/wWCT+lJZXogoF3NJDOEoMgkwMWhHBR8UJ
N4FsiG0gya2hzzYZ2lAphNtrLsAmJj3UINRR+mrcS0Z3EQNhiIfriIIUAVzd
hRQSf7BRmBjyalEV7Jfw8t4WJIOlefE9N0zVs+CzqfwVxHMy2B1npaQamak0
bABtHufzdE/RpmrNJahLu7UcM3ySteCMMmTMxaGCKAIHmYTSHVVaJ1aWhmxv
U3NPV19ZMl1uDZxHNY3SKv/eacrN9x3Wsj4qP5TsVCSMeA1694PpshPT2E3U
BdfcvPDxSXj+wejuqJgcsXBMpkRNHuZYTtNG5uGfvA4USJSNQ9DvzCBSGCav
P3oa46AR+zPawIcBqYlUA7uIdiBx1q5TQA0VYsQTNqDJKYAjQCTlq6xV4yw/
Mb2zZ2GuuA5eouC/VoClCrXAaEQuSRd2laTa1+23noh2OPDDD1h6wCcFGIbP
O9gHQnIMQ5rnx0sDGqB2i6RqDpnMwN8ADSkQCQF4hz03Bv5QOEC1JqZ5hwrp
ZAKLAQ2SlCRCpCD51HPmx+8hgJXCifcm6rgxlSNJeFRX8nEkwvvYDPrxmbeD
rLuaLGUBvtMr258GaafS53zuhi51/xP2nqk07WCPnQQ8HFUwXWZYgjvzWQjS
wRhTO/lUYN5M5dHYDP8F50C6YKBUCAZGlUMq4fEOTL135SuEspgoIAnwacpD
x7TmpDCY+2ObZQB4wvGEBi8lckOxC7Bml4Zs8B1xMd8JA42PQ23I7QVFDp+E
TrMP8DEFQarQNtSLXKswiHiXaOqnbHkiWFwcZtz+KgZfaHWOAeuNAVkNvek0
BNkfKEITWXxwk438ZzJD9B0nf3328CXFMP0rC+gMVgaMn0KYPROtkYE8UVB1
0+omMnQ2cSKxV36Rvi/BQf0G6DDwcDwif5Vo2yRsGAvtfpWuNtxdsGTH63nz
W9eAtGvIa9cw+7Jy+7DLVad8eYuV5YShEAA/NFoGekPiREbrtS/UDYjVVlmK
iXIQFWUXj5ljlBm1+vD6IEAIhcyVCCwgS0ab9UAsPP9AQTRpaBpivep87drY
1P/DT+5DXEZGDMM4f1tIHdVMQdmniB5MCt2UWloeelicPzEiGqaAOPY8punY
UBqe82ZmQTe4rSNgV6z0eCeFVvBW2v+6EisQ2F8YUQA8E1QDcyF//DaTmjd+
9NggpVzUu5QsvyXfJElIarPMFBoO8C6hGx8mKYSRQUxxdf/OWYCVWf+VxZ0z
QL4Q2sEqSmgnqH+8uMdDivQHIfAyWxeskw0NEPHqeFth3wt1UGF2b05xoVj7
f1QkmZVSAX6NbHpRRroh4HPkam+lfjAajIoAZaODWuJpcEOsKSh37Mk7YPfO
5tnRpFd12fl89JOboDnZRGuYWOmapLQ93RSvVgnjOiyvuraWVpR0orxoHX3q
YCGV++BpXBkuFWs+uQOdoN9wYbp9mVwOLnrRSza9p1sXTE5Q65pteYhGcypt
vwRPeVQ9rVUir0cViZZ2p/B+3gWvExlU15a/OfW9Pf+6mEbY9Pt2Lm8BLos0
HOhH8pz2AUTkvT4YLKghZO/LHYS15eRKWYmhxfJWBci2bElQmIKRc1fHW/n5
iVvRKEpuIlx/LwIJXaa+MgiR+fWZwsNRRSf95Io49DzW18TZZIp83ADY0hPC
lF24fm01uzrL7JodHHgyMioFwrHAycdAy5/n0whmCZIfhofaA8kPGe1ANzbz
HQaC7rY8NlM2uGY9ethwi3jnRtqx8ma3ewJRa2iXpqQJg8TgpHsuiukRSg7F
ur9eWmQ/Pz90vsxgQ7/mEGNNjamQ+8ec9yyktDsDV+dai7Wq4i7DtBcaGkm9
G8Ab6O8Sbg7njmQ39xsEJO87gFZmc5ZIL4ejQqZw2yu8d2MfhlUlpvFCJBB0
HNCUl1waiwvDoq3eMN+Xzaad0ZvrMBJtotg5ubrRICWZGsVDwSdDCfrmLIil
tS+TbEz8WCH10fHnklkg1BahywlzfSiJDxYVcqHvjzA2bgPk+M5gwxnLOfto
Ijg+qeqOQA8hOlEDZ5KcJKO7Tvh+addMtHRgT4p49uv94tiWp4EVpa+sjxAU
InV+MI/AYa0SeVyZpsfsflqQ8DtHLu5eWIReCwJhdV3dvnibyBlWS/bzaxOB
JwXpKULG5UJL6x2CPf0hrPlnJsDiF93Kfp5P+UM4LjrR4tg71KvXxln/IS1t
I9vZnEgHK7WzxtIF+jzivAGWBKy3qf1oS5TaC0gD1RrQC22UP+XmUJdSdZTA
443ZF8VrxlubOrs9/7zZBPkAtyY7zpeAAplZMgo5NkaOUwNjeksD9e8MGNLM
5S9wOcb0ivTaFcwCF16yG61yYNURB3CJEm3e2CN4dbuLqotts291Zou2mzll
wkAozqEM/44nOTm0fSNqvR+aCkWuniLK272zLK+0YuHYSe60y9luRIpV1e4v
HlmN2rz0/pmcE7r07F5v+2lkwuAZIq4ODXNP74Ercxjn1Uyt4gab+65ydcAM
Ek7TMfO5t1Bm/NWgKxBDCkUzbsPq0z0nffnyDPNx7ES04/LQEP4fxIYCxsp7
ITodf28Bsb+jbvFOcAFRxW9KV1aPG05RA+B5iKmMzXB+fymqcGi1CL3/8Ym3
ZQKdnXwxToaJacMmIPKqf3Pwmjp1jS+KoXKkvBdRuGLb+EpS95VTMkLDkSgO
ixC0G0AB1WwCNbib9RAisFzfSUyvUh/Ky2fNFUr1xlX5i6viBHvkL6xaKiuP
kzMRNVUt2YV/ypp0V0ZIp6LLwm6KXLbFLQMWexe1Ctp+uHeY+tqmYU45tTtS
J108xpDaKR6Dm4M1+TXaSX8xKztEpzQ9NlEX+KHY48TaMPvnmSk7KcLvCkPs
Utg74AqWHCDFXWb0FozIJTJUEOBFa47S3phZfvclryOSiMjg/5egaNlu8drC
snVvJIe6GtzDCEbc6OzF5ePp+sE0N982UBQHcW1C0ltTcreP0mDvIwljaY0i
hzRk8hNzOQBhkyYfvjErP0q9Wt6aC1Cqji4ezFQd1roshgCVL2ChKtmtgitK
brcfQ1+iC+byGa1QRvbcQtiQ0uGAQrEdn/17R3vRbeNThvnWgkStVfSI8Pjr
b3fLlDEJbqdT+OqW/ygBAywEfJl/pQrLVzAJlkq16qjvrEu4JlFAuPtMdBcP
G1Ti81roWEp3V/QUmHKsaTlxLasef6dcJOQ7/fiRZ8uYCKEC3XLJif8hNiR3
IymFoiemcj5CJJbVA37LT3dTUwwE4Uw5houjhNpBvt4G6mHzNme7oViKu8hP
8ERfvai7W2KZL3ljMKy1KspRVi5HfNq8ghxXWr1seKzbYDx+V80HDDbywGeI
DbwcTj2ZCGYxSGwjLMJL+AV1Cuhwg0JKHpanXOtE1K8BwZn86df2TOGQ/P9z
pJKTKOTdZZAm+D8xIp90LXYcl2XwKBvdtwdgs6AFiUVuVUAg84qHMPFg97J2
sKkJkiXK8CO/VUJHr6nGHkb5xfE7MIVmd4915n3jUJWYMegcdwRtiL3SCWzI
h9tm4tsKh8b7DxcOElF9VU11KR7Dv0NgC1xRe6BlbYpM3lKGORDQfp7UhOsH
uQcznPrnQtgtoXjbXFqClvDhBIh0Af4yXwkL9eeX7Tn6qJ8UnWrd4ADIoAne
JCD8tm52N0F92pz2w0J2IDvG8JabTi9XQmVqIFkUaAt1k7i7AAQ/tpznE7Hy
h97KJDc1NjYCsXNPS2UaQ35P/CrSr0eKFHAqo694ihKns4vMowz8Cl9HBPyT
Cmi+1Xjnc+6xICSl4Gql7lV3SsJVOG8k66Lx/sdQ0LZG20+QNrk043ZP1wTJ
XAQWdvHGfVZw49tSScmonCOPvD4zS43L5ZtAORt4lUqqHOFPqb/J0LzMp2hg
/yIipftGJLUCuM/fnvu6UHA6yOhh3y7Ra8qz4BYPqKd8fsuh5eSUbZqFcThc
QzpqzlKykizE/F/JRWhwmP8V/IshLcA1NBfSiz32hFvuWk9Z+Gd+wXrUZiJg
J3nioaDDf1Hkn3jtEGxg/9hNi9ZVmnTGZxOoO6hHPAYbLBgI9ea4nwlfOEGl
uhHChfO5T9H3pII6GgBJ6m7LbXNv5c7gBqnYLPcJzo8vNmWTbuM8BqsYotIz
LR0SMfyrzvI4wZa4CyZoSFx6WAqihFZyfG/dM6Jh3KSMWA7MVqsdy9gBwrye
7/ml0VsgkVV/vdyU29ghhbClorV8H92DpS2g0Np8HS0/3WmMub9b4/ErsNWd
Vv2TzgPbl2x9FyMnOOKbOVRNExSYcLLdsXIcy85IhvXHjXFKvslOMDW0b3zz
BoOGuM19P+LquP4gYE0+pwoBCTDXzYNu7hlZgzVbwf5KjJfEVIYuoQToDYbn
8vKRFLDlqSzoEUAwu843T8VIUe9KqGMPSFK8qKiUv+t+Q9v/kyiDXJUxKkam
vMMe0rIqc3WS+lSpkxWLOFH7NrSzjwhN2MbpdZtDP4r1FwnkM2lEAmD8U2eU
k+PlKa3eNn0bmuODayqCsRXcvoYdZuO2Drmw30m51vc3QhWTH/+d79n5ZPSS
2mo4bG2kSK4dp/J0xDPln3wviQ0AlX8T5qDEHtLngUnEPoU+HNlJdVFAaP/K
aDtVGLNt46dnooGwCECkBoXUvk4awI8BPMwIcC/aQZwatyeusroWpYH/gNZV
oKiOJ84Va3+VsKoA48zuRi5yIS5cXs1Gvo2DJMUoMTxqxWzrcRZNLuZCygyJ
bVtStSwrHrl36Y2NGYgPfFYMuWV7rM1ON1OLYkRO0w+t67onK2gRM+PnYRLh
rLE6YPFUNS4xfHkH2KBB6hAPejUukSSgiuC74zBRUTYDqZkzEWw5flh/048t
ErI6cImBdntTkhX3cpCDLCrkN9toswyIo9DcbXlEzCXaM2IO/0Qm7US0lJlC
y/lCjy25V7uLTkUDPSuIL7mJSR415H+Ni+1sdWp2Gwxvje7kjcJhVOrZcH/c
zv7hmwKwJbgaNBIIBhfNhuBOavDC1U5R++2ObzTO3FF4FDIu8CgOPTc279aQ
Lwt/fmQWV2sRHQOfk6xegjkeIvgAUfvKR+SR0N1ZAm08baOgU5J4DtUHTyfr
kDltpBAAwMpVZVuvmmSV1mTawsyZu2qPWAs9WT/OuVXzUK6FbFvQ6+0zM+jV
BKK1l1XwYBoHKS4+Bo9Kl85gUX2D4BvrI7+oL7aeQaDvkeZK/CiXphbAfTMh
TyJ/wsQSO/5h/vdnWYsVxrBbM6oULfYWb1BIJRudqSURc/2Z9s04DQa8eTAa
Bc+TRptA7DMaG6ie4/FbJ2uW+um4a9sRDmHcYitVlQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzd65y1M/BgFaYXJEdI/xV9Xh/Ka80puQoKGa41kmWMZ4iGn4ft03BJvUiBFn4sAxvcpu5CfVefHrhs0GvGVqRP2b0YCnY7I894/CKqZWQv2XLQtkhsLd+fLj5AqM4JW8kH4x+cP1wYVbw7OBJ24+hKaTeJ9IrA/OWPRVtyTzM+DwxTiSUCAMHVHc+IVcywi7dT5s5pygQALkuSW+4aCjulAj9Rb71KGJPdBiREQ5ELur3Ukj/Lf8vxwGAOvixTJ28CYFpVZiz7Viqxne4Pils4NI1pDSgXkXAk3kXTpUFKa5cEgL77zf4AkITtal7qeJzWDDygPgAqC08JBhyx2BzVpbYCuTa2o5q2NINtTsg7TrDC9AgiBQggO/RSBZTYcbAnhzm1lfLvvZMqWHQCcrBFbfBhiVp4ScBAUBooRour0v1SeqkMizeT2UTzbdrY/9HSiqT4wgz2PYK8ByJQLJFJiKOYBRWyR9f5qPptBM6HD35feFsmWFYFejyW3vdcwSoqLttlcr2KF+QptdPc7mat8BtNWYjnn46cMOEQU6sfFK9QOb41+WZzdmy3luudswlsGY9ibShFmOUnaPHJ1GB/m+cdKEPXaREV+HTAnPklXxeKn6eWjAxNYYwTgPK64npfEViS1f/qFQZjjYcvFGpcHckJgVBnulSMXfbK0HTpdlx/2TzWptD8bi6iVD2qMRc591KHb+nSK/VzgiNdI1AqpRcxO5vkyawSMKayPPJjxG/GdnCKkj+w6jSNku3KrpJ9vp6w9QJx/787swUsdnfeR"
`endif