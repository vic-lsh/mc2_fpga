// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Iy3Y8RLCHE5LyNjetwROnBk+wgKxT+DAz+zAPRq7gnw69Ba9ecj7Zoef14ti
jeqmIx0yd5P2YhlkcNR8wBanlUjmTrkEOla4iZzWi7JnaaIBdAFWmuH2Fkdx
f7x+2lpB9B4oPKP1bB3+fjTNkuF4WUhFHZm4O8uEMKJY8hzyhYSgxxAfNR/w
WmzfLdG5Ivq5kH25OV9psHOm+0OOFp7NG8vYiaotgpudaKD6TaQMRZAgbGSk
dJUElrLekUtv0B8ibEV0MO/QMFE4ey+hvssOVWSivmtqOb5PN4IYXmu4DBCf
+MuUtFFQYbDmTNbpY4RCc5oULzMypjAqS+wEHHOxNQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KITJelEfvqFsGdvXm77vmuMBGSImoOpAQNybqXGXMLyyUCkLr8GUYqquHrwM
MaoM7x/FH6UBoi2cCDv+k++/nVEU/RjbDpmXllTj/NMe1ByBoiDw/cqocqJO
3AFQz+W0buZfvI+HAEIt44hJ7l86HP/BqNcqTcQlS+vWHOmM406dAk+h7TcU
6Rrs7kjWzpE5sTG+8Sx3g4mDWibq1v+pDqvrFzjd535etqBgwmahzWDPeXj3
h3hzXMy5+wZjumun/q0ngjfJ2kLRBHpW/FclhxGbKSH9BknxYoj4+DL92mhx
g/uW6Ib601CS153grEC67ZR0Askaw99f0e2sbClEzQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
am9/B/ygd4phWtz0WD+WOdp5YXHBixjlen/PI4RrTBLTYt1S5v+M6Gx6Y1Fy
au60TXYH1ZztDSu3kHuafw3j9KJpBT8RRNh8x4M0s2iGRTEL8EKvVOfAvuJT
Liz6a3QQaYSW0vFJ9sguSp/BRvaBVsQ5DiXEfcW+GkvbCn4/Fm/kH0HztP+9
KzojGblXtTXDAivsimoBLoNFXXorcIy452214D2QqlimgA6SZ9ympmRbS3Rq
o/sVsVIbjyT/7fiP2I1Kr7q+9jmsNqvNearpOWr7kwntofd4Ia7F1doRo5Cn
Nu8z1ZB995SDxXbkgsdQi6JQnqEasonjMI9nD9Q8YQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WnBC8hSf9nmKDDHi2UaCHj7dKT2zl9WFSYtTKhLiMQm3NsCzbmrWowRizp31
J0XS/eAy7Bxh20bU4gLRG9Yq17B8sWSYFjTUF9NxMDmU5GxfRWbTswzR82LB
lzodICH8656hZFjhJdfs+r8wI22gG9gddpLTo6bcWL9O9aBwJSR2Afb3yrvk
5aR6YEz71WpZ0b+iQoCbEcKS1Hv58On63XXFilPo4fjPB8iukpXs/eDFSG3W
8xiWNk9VRmWDDY30LXXg2C7FNwtaH56uaz5u5rTm2NzeUFLi9/r5DImy0MR2
kXuXIZKihVXElZMdAH/QvhxSf4TA6qp8Ryg4ISD2gA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MGGVBJOeICaWm9vZtxIIWn21/K/B2FD96zn/tlql0/gFUnWlS0BF7Yd354Mz
YDrg3SZ7WsRpWe7m1GBEKHdftxgHxQ0MIqgD/6uECg3VPJnyX6BwLwr0IR2p
7OPAk4RFYmHgaMd04wuXj/eWWwvYSTo1HTcOIIJflbWyl/KhaBw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
lrnrXYCAjxOQUJ+XCN2RlCGIdipUQ5vlMRSiRiZlFqNM9uesxcFWTBleaPn+
nIq5U098zl4J5zYvP7wR11BqFtgTMjidj1Pux67xiixUqDOq+Ix82fKqwpzZ
s4c5OLcNMqnu9Pvna2/ZzC8qnQrNyJ/UNMosB5m/gujFPr2WcNjgajnvR3OC
laCIiknOrgHVsnOhtTMEI1yhadvwzqSCMPk1Ih5Ip4cNqWCc07tPHgmx2av8
13cZl4FqqpfD5vnmv9N5Sg6+6okF4qHQFZOP8C/RyWtQeo5+hhPvTwOWDlLA
5+CzKhXNwYFXGpswPK1bfsIvWadEKhnUqoggIRsdNbcTUEdB2BQpKxSzNpxL
6apKDXAM07Ks8rGMTMACY5EAXlJD7y4es6dVolUX2QFUnjdfWs/ACJM7UWnq
nRfyIT0a9Nmot8NxxgUDrvE2oK+px3mIhvncT2XxDbIzNRrTY3v4PpbA9Sbz
eTmw1bppmkgphzQVBZCBizLjrDcUpvTf


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YoM9Fj8W0JDThLOtcF09oVOVMbZbpjl2uGH0xxJO77FcUKH5tBrQdn3+Y5X0
dcXScW3VduYiwaOQHQggAVsi/P8B00GK925q8ycZiUDRw/ox3bisnE78kL3i
m57ri9ovkBljev07v/fM2LhgoJu4fVhDEL1SUiNNfpumv2e0HW0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Q9hXgYh1/TAJ9aEJ7gzrynzRvJwlGrlPQyw5UbPePpGczDWtHnpKDxNlBmnM
Jk/WEQr4fz8T9EVMgUeqCV+3jOdIOjWH7jWXqa2vEfy/Umrfq4HZL4z5FdIu
7uUaRH8tFj8WVOL1p2b7/gUgg+JA5EWEHBP2XNxPLIeGelTLe9A=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10816)
`pragma protect data_block
3hfrL/5ZF40DEyVmpa69Xgs7b6WBvkf1kx9TxMCKsw8/bx9TONO/sfGwYwtM
8d3OImh+nW4qLE5hm7P+p0fQdfPIWgRbMCfKyzAO0qd2kPSwTCW1awlV+PFS
IZZBhmypAfTxpjTRyOcj7n7aE3fM/ovIryEGI23TExWvy3f5VCpqJ9Tr2qOx
o5B2ll2KWWsfXmUv09jVO7gMluXamZzKS/SrwokKY+qcgm4F4Qj2n1B2fxkm
ml8od8KcpoBa8rscT94PMrZHLg71BHaw3AwfVdzm0V1S6g637nXhwjV77Wxc
m1/fSgq0BB53xUzRUUB51Pm/n825cxvlP6qKDCKnDB9AjVNCmdgBg+8odbJI
E7EwUCj9Q1irbXLA14tTMkvaFP79YBCc2vMwF1H9KPyQmXm5DopK/NyZML0U
tHfLdDvmviEOxct29t6rtU9PQiTbDiWIu6xqvm9Vnut/7sfIszl+ipGdgon5
bR4LCi/X2RAuIhqk1rcYZg2iMJpkVU2giwGx/bm3cftjNGJHvnAb0vQP1Nxs
8Bmyi3HrRXeekp9kTt1mvAHJJssIZ69m6vfS2o2gh0IQ+moUfw9pPOfuar+N
bC6FjQMao1Z6su3Jj8cfnTrVhahzT4eo/pjGb8+HDdxffNvLK0GTU+qEu8em
abJ++Gx4FpDX3DKxxPz400rerHO1KFJ33TvgHSLhoHZhMAjckQLHVeIwsJrO
vHUkUNmUG2EkK5JnIumqkh/aL+A7XH9iqyo6fEralXS8nF3JvU6WOyi3uSHP
1tEP5ro1PS7EcH0CghQ26KsHaIr1NrxmG2wyXkp0mCsdJ38KJ1+Z6EtyewXZ
UeDWCIfkFQ2WAm/+pgKFT50six0arokTzy1Feo6KgLidcPVbc/bYxfrXWYt+
E6z1DLvaVThYwkE9lduYB7airlQi9ZzzaVqaQuFHH6iMWA+wJVZN4SXNMsz0
zzUSV3Q0tbZ4YVlQQcut05NSVW5mjoSIjGXrTAzNrxKr0LEkzfSr/S1xtHTE
b3xIaqae89W3FrcXd4GTbY9Dg7V8ULuoJcPpN4axhJkgFNcaeOJANLi4CUFN
naPQkmgHJbqwZ7h7m1n8YSICW3rA8keIqGVmNu8z/VcS/iCuTRO9LR2EI2CU
TFYo15vQc7rXnKDkrhWohk11p33wccJ1XEgyaYLdR4msEnKnHYVsxD16kllz
ZK0Mhz2jao+s0PR8PguMJQ4LAez6zj0k3YOjQl99P2n6ZzC+M2FNJ+R4KskJ
rJSqJvk4CxIqJcFM1gp48rNMnWooWHxRhCF3HilPpOgPa3+Cbw21oY1yEbcL
Cb1rVlz7bUX/1awj9zmMXYZ+js8J7GWk1M1OkOv0T69vFPApKp4xlnt/gdp0
a9AgY+fDBOuQcA3JrVuF+CmAjvkIIYTZ/I6h9fgRCXLX2dWBbkCWw2/sWCnc
EMPh3uTHsBrIV7gCMQWX38MQTuhnK+NNDlHeXxLvvt1xokpoZrswM03Ck54Y
DvTI43GQ2GHmpqITcsdOQ4OTrR4t/iim1Leeu2GSjNsKdARdKA+Jg+5p2W2N
mN9MugdFtT3l+vFv6Ld0jtch3ARKcqXUhlZe1DpA5hVDaSTPQb4qKxmP/Bjn
Wp68cGntx/6IVNsBVPIXln7G37J4A5RmdvfXn3OpncvUIrqRs8ycn+NYvpl1
Bi4tI2vIuTb0uhMFW/wZ1wCxuMxgSS8xqqVJ0AwCd6446PKICL+iW5E0IsXZ
+QbOHy8D/aRgF+iA0JDTfWviHhT1pA0GX/EUxMApB8+ezN5Dn8PRQ8plqeTV
UvGA5rzSkwGrpJOqK7efrZtxRCplGR3H2iUcQMtS0YJ6mOlWZX61wGu58KO8
RHJY76f3dsmuFg9h+kbELjnCFxNSxULOkyO0MlwmNyl4o4AVdKgPxlDmBISG
Pbxw3vXKu8CfFTFO3j111TkOtavq9B8LzHeyzwDK65gXRawgd3Yy/f0HbBdv
zOiHeUvZURedEi6BIZg04LIJDtbT97bno4TKnlSTla4TqSr3T4HxQZAVSK10
LOSlj5bSJ/hPLPyB1F5+MaGiLoYse7pGFQf5Jhd26VZ8+J/V41g5f4aSrtTM
HNzvrPBhsaQQIDYzJ9a1VwrOrJcFhuv8csh/vpztKY/yw4TKwqyFAVzxkIsL
MOueoo2g3zxCzgfhX4e693BeeppUxFLxDR2GmI9vSPiscG4FI0ohaKxs1mCN
pnYjKf2sYi51qTRKEjNjMH7oNCe70XbkLTFj/Z5b8dt97uV9KgrePiX7Z4Oc
enuxjFrxtM9/lm3HWfcPiVGr1sEGi3yP9FO91bJqHqC8JjotqHIvtrwhtvN6
R+J76+LUmxsDFbyc9RyamJwitvKFHrBr+6PoiCN785Tt/w+o5M+r7R9TSV3J
sHHSA7QCGwq5DRjqqBAE/6x1Z2TLWLyPwbk41SiCftWEcN1zJ0jL1UvScSV4
hPwgPxSb5lLebLLnbqAoDXIK9U9PfIB2yILDaPR5A+vIpC6xzAtNKm/oasdr
Xy7YVkek1i2yNtBNlL9ysA2g9EGkXA5PFsEqBPLQ9G072o1V4V33xVZ1mt8E
UT5aH5heHeIxjBo94yfXtP2HcoxDcq2LYbmzivg5/CPTr8RE1XdERGthaIXq
6sZzYqhk1lv+AZezZl3ZXinTMV4VzRAwJ16Ip899wqrE73gXUvyQckbPB9hp
cu3FwgUyasJHCK+BTPTxjZsdTNkAIBeSfth2UHq6vNSM3FlDcNViF84cWbRI
gyyiReodhzLL6kDsjVadu58+r85TIim2wmZ/06DbsgxgzswTF/YF6kFojRzE
Enr1K1xgR8ipi1dTyExP7bK5QtDK7MgK5kw6lQXOjNFhC36pdeeFWXdTD8mG
PBvKb4+bhTcaAbsWmxCITAuEDMqsZIhkgRJwN8YAUFPmyArnPpw4eXpRnK0m
eiu/ohF/37qhktX3FuQdwYfpT/85YV+AeCGMqD4uJIh8aj+3W6+dcdBuCpEl
P74WAgpbyYQ/hW/nsX8tbKWTqvFr3C8L5dhYbrUjS7c9MOAtEl8hEQDJH84A
Sncq0qPMV/gIIDZ/7gZL51YEdI9K/Csn0ak0GnnDj4n6SojZDFb8JOOhc5Iv
vAxbNv2VxYcKu8P01vQZMyzHLCXBRBMDHMr9GWxzkrEBQ6zTiV/ePwAo1Lqo
+GNXsLmW9OKQ0OBr6Ivm2C6h8jWqbhkp1HNRXVZ7GkpwYfRHa78mWqcTBpit
uVDaTnUjb9gDBGdkrrQzNu03MVrvn/DtrhItzVSWFgpyolEEmG3shC2ybVmo
FHagFbGZZATb8QN590kiEQUXL6sp97mUdd4NcVQyfoh226fNLGYjw2bWEDbX
/Y7zYje4nZ3Mp0EliEITOZGA+N2+gXMcThQLnjCxhpHjFeMFlIwyrkFkRNNN
8LgTwSxpChC3j492VWmHv3H4YuirM0bRq/oI4RimilmwLm0/8cufQUtvG/d5
iQkHoCsBGPIoxGXNipOGE+sTyh11r7/rJE1u+2PgQ5sqEhTXiWJf+L2ouy3h
G8Akz8mLLmQjq+4Y+m0jLYF7dRfMOQ5qf2N4KQTs2k4ESug96R9gGn4RoUQT
hnDrStEtwfUxusbcTh9gzv3w/tkAaB/hBdIoWbg2ihy5D0WWy3NtUPevo7TX
rgQIhVB4HoggT19LkpUR03p5zDa+WRlTyEZ41lJzNYRGPcrZRiBaIxuyMxvh
f8P1sjBmtHIXrETw5/6yKA7eQX/J/WtEkmLslRZ/qXU17diDC3F4591HfWBh
USVHsgNjs8PeE3wXcg/LPYqUYqZGh2dtcffYpOvHUvVxOyxIdH8QYLYK0nNA
s9o8C/sfJimpvZ+tAHyrdUnafDIwDrx7GSqDcQPmtRIOvcvq18YLAX7VBuqV
t1wLsRtfAu4DP8BOmuMX0bKdMm3zNxYZWU1t090qyKcLTwR9qrjcDqp+b7G1
O3B2Qy7Kwhbg+zcc3Cw4jEQ8mVBkL+xQf4suSsKLvZ3uqi9kgiwJxgvqM85z
wcZKbNr1OXAxmDZ/5kyDbVh/p3+Oz24xOb096c6IyR6KYuKRy6HBnBSmbG9A
4b6PqiX/Eg4+C4Sa4nnWAsrC1hCOylZwjFvgW/mfpcKWZqV6mJpYTkLbCTBB
2s2AyFHVYSJtkIzlctYshF1nstypLWZp1WtjzG1jdSCwOMhUJf/T1Jb0BoEf
PXe/hiLU7yOOEsziEstXloYjyDcIpD+5L5lahjaOPE44hfSphdP4+cmnQdVB
AeShREn1dUki8pd+VF6x55XGbwCMpZVAXUme9nQ+PKOIrdAVd277FzOQxDSW
+lMU5CgoQ7fFmMZGMPmDACyDAYCeo9dNkf2mlMxXOlQYYTLhpNKqEqVM9wGu
/dzpq7ZYQHNqQrovlKA9vDRCm/LKtnnQ7qD3EJGcgMRZUIfRr5L/VAYWFIeF
JXHOmq30PFIVGgWNqcapehiG0xoU8023VkDnB3fbuysvhHddfjHjqzK/boJx
Kth7U2JtJ9S0wJvUiufDzwfP8qlaTZwuQAgklnJr7b9FFJ3+nxdONeFp7794
NeKgA1skfdor1BThcep4rkfdA6SYQu6xzT8YJe85tHBA5UaIiVjMx2vq8Suf
Ak+CI3HDFiqY8m9Ufoy/CZGcqb+9vFJ//qTwWBdRJeCZdktHdWV8XX0s6Iiz
NdY7EWGAojmADZCL+bj5axntnzW48Q9UxH2IB0qjoqgoh0RvRLC5/BYwisRl
UQon2xjomyStLvhh4EqaRCzjHo0NczA/izcOiaAPqiTdkrt0guCm4xJVZqO2
dhVtLFgqD+CpGb+fsBFP31hBL5JLx9S1DGDPk4/Ih/gCW7pvi7uuyBZTsVGC
DLhOyZmpk99vUWmLIVceg7iZ2sjO8RiLmeUCm5XNR291Yfwt55aNzIXRar/W
fZwa/cCOc25bsHFcEaTFS9mlJ56pS2EG/BwYtJIEzt2wTs88TRw0PG1q8LGm
ToX6bT2K+u7ubvucOc6CKWGuBt018opNX0JdmO+EKH1K2iyNzJJOhS1KKgZR
bCmI77FXsmveFnLHU0qYLXv8lOwg0JpOET/1SdwhOO8PcArtTBlGyBeRb089
7lRen/eRwp6+Pw6jVehYG/xM1tjNGX7j8O7Sbx/JsxXOJS/x6o0U/tHCK8jp
nRpL69jXOYrA4Qr6Bj0CkJLoxXoQV1pETcupM2K4GerQjsIX6FzUa4xXnbh1
GD5YhyYcf1JXtPYC6cS1iuYjsqjJwShROt9p7DKrMF/s63cxI23okyQQULZY
ghzDWzmqlbU0VgkMMJAoPxcY57jizyV6eSZOL3ooD9BVggwwpRqw+TUxgDv3
gGjWbbykKMnckA0hjf1j33EVRTrDrYLPWzisZHYoDWTm/Hz5UOmeltS2pj8f
Rz33zzii84zYsIPm1GOKHzdzUSENr1bMKWl7CxmA27ThCX5ehWt7shkLP822
KIV3jOtUpYIMNlIQGV7G88uuD9BW7mijwhWtatRgo3Z8BdM5x7SPUOYevHxf
vLKfa9i3LYojayatndTDu3hHsO5KORntPZERS/bt6O1TSuddCq4kGu7Y0Itl
FzU91OxA/ecX58+nfPiCJ4rWNtocZKFNZgdxhf3VCRAMNQbIo+wdUSMqiqAQ
G9ejzMMExY35kRgwTwK9I2YuDD75iMEdBWpd4G38uzVrJrRTIqr4G7Ulmsyg
7Nvvf4a95sGV45KxuB9zpx1GcDw3mfEtAyeefwUm93alaV9nGaghzyxSoju0
1z6ZG1QyjvdC69oODpswTEAlOEWgR/GyWYC1geNIDAwz4cFIL0ehGgIeJwUL
r3QDzZxjkI0LxkNzGXP1cBS7C1JN0G70WUDysRnHL89XhcQiNJouQYGhOZDC
bgyJKpzfmiV9vzfgT0fGIIKLsouRHemLpeXIaXOaESMWNwr8XN9pMBeBtbcF
omvxtO4wzUTr0GSYTbNo4W3l7Mvl9uJbIX6MTXTgEO12BeOnndTMUkKQJnSE
lUA1yiwZbiwUkvji1CCHUNoGuMYr3hjf8iBVNfPiFZmSDF2hq6WUFJ3ncPk0
cZKBmM6dsSwL+OgTSocCSGnDHfOHLbBmrUZolnjzfrzaPM87+8Kj2b6VsAmy
kpe3PMr1fT+EA7oftApMgMZ8CbyBS39RS1iRKkVrFL2F9Fih703XEimVN3Jq
0D4mfWON/HgjitTSwipyZHVBlPevQsVwSQGexbG4pzbBzotbu+neypR/JP5B
9n4e7xZZTLoKc7NUZ0O1/NEJzbAdmH+hEruEd6Nlu/Q0zUSRH1XLHPYaoptP
jXJpyx6HZDZfRLLnvanfivJmQ5V5TMeY7K1s7A9zvUY/742oNg1dAHeUvfHb
HVSNhcJysFY8HObCF0y/Mj9HOweNHBEFw6jJV1bxa1dGG0TeNdNXVzBEk10a
jEdUs69l20U1pLwWRzUN9jFmAEQWpucRtNSBRX4zL5FF9AwN8NLx3fi9uI0t
tTyUtNOkueio1eaKUcQ4rlkxp6SzA+r1KiTzDuoG6pcHakwCJSO/j9dMA7jd
pJlv47ivpvyyjEoLMTYmqG70Lwdpf+Dka78K0zbKqyN4VZBtBHFieD5cq+O5
6yPBULiBREvuA53J+FNlghEHxJEMWP1tJkMj7dY4KZyAzQcF6v1w8KC88bo5
pzS/7NfrUcOnugvUrvR5VcfxmIlpjBpkqxLJotuf+AudfaGelalUSc7VId6Z
A85dtBLb8Fge09lG8g6tpkLeoRuAKGPvLdnY9+v3cy6m0lPPVUSC8Fzbob0i
edCxIeNsbNU5SncSwZ4vaAI+TbS+V+dNKDnQYYoqfetTeX5nj7eU98bPR3cn
mk5+HKxgjJc/DTxlCVGcWEk+yLEkB27n5b9K0yRjwu3m0DnehN+O/QOchedZ
ZthTXZTvL+ZbIM/Tg6P0ElIG+av1l78D1Li76nK7T31YpAJw5p0PnIEG/xD6
ekSdsAIw0+a0ku4S+b1zxNfej1uhAlk7eG4/MJnc9VRzFrnVIxlnQAEflFA5
rP/Y4r5dlHeOnjYNil8ay05F3rwZkuwiEo+KNyISLDhP0tl4mI9Yt+rXYLZq
ONgzIQe79L2WP0N1c2r6zdr8P2ipU8DaHikR9wmOgJb0DCjZftABG/gMxBfg
n566ZXtCbQGf3Nk+5sjBjMEEH+xgMPhocUNH96Ye+g5tif8nPRv4yRB6EPIl
uS0IsSewuhwkNUrnJEjZyGwnEhaDb1LH03PqrW+vQbsHC/RaPJiXH9rQY6XS
IWM+DvA7sCrryAJ7nY5z6qWgtYvKcwJnydamCQoC1oLFyBZRQPXosAV06Uyi
EdoGOB3mbYkW+Je0JoKF6gPL46g2kLmlDpau1TVoztCp88QiseVnS71q+MPQ
ehnuo7p64waI+m/2wXWTl8WNDmmtSTLS3NkuxzcNnRPGCfPvGTvY2X96mZmH
MY4sKuk1395oSUv/DKt11oS0W6o5seVpD0KdOUV+jJwdYvGF5TiNufvaXkTH
xZ56iB3rmub0/mpu0wlSKN3dRHtL1EEXOO7geHumhD5E6x9WXr87DSQ8P2pH
AfbQfLhLXmsv08vHl10c8Yz/cE277beeWqwONNl61nq0PcAuR7ObXx1x+W+X
osf5AzdPjD4tWuYnA3YyXobkeq6JkXgOuf7K5qjq4Lm9TBnHbuNw2AH2atJV
VB2XY3YWO76M7Px/oSXmTA0HleNfxRVtyBObUtwoeR7cnJs5s989Gamb0P2t
Nug7G7byEcrdQtULm1O5l2jT0wcUvsFRR3+O+0cfAGdBohSK1haI6Oy11x+5
ajjEVOHuPQmIoFCeSSOpytN5vs+vkDlUfRf3eSE/od5OiFDZH3fCXZxKs7hx
GRO9CLENJl34Z3ixhTdrRz70GUGvhJ65gIg+iDHI0pIgvTw9EfnEhwYxMcL8
YIG8FSG3C/N/4MI8KRK5VlOnkUT4AVxgdd/Houm3JbsTaJbbrCkihv7I+nAu
fCT+cZH9H0CwSuFvhmz/yQZfXsu+dUmwiBqJif0QPigPExuKb0g3XNdQD4zP
94MuAGyKYObHsNu0PzcsZrEdU+u7Z/1eq3GCGB6O591zth1f84o1sXIw852/
XAb1e+5xzz/BdSigCP+wDgM5XK/zAD1gje7jLOFSrs6HGG5hTDwedBOViE/+
pCZTSIOWdHZsrGUIYkIAj6U3mCg2KOfdBP4gMTZISTf1WSn9lFt//YhNzEPd
Aa/R2XAZMODVIRu4tLwO6MuuMThKoEd7KwO2WC5YbUvWQswccZ+9uAOd/X8H
AWqayIsznzO/J7Z/e1HlnrpkGinvBUbTWPi+E3lhLhIpaIELCPSzo6tKmBSJ
53d0xsBcK3E1Y23aCfdAz9mtodZ62RDAEb3k5mtoZj5q0AlRVrdD2CsE8aGU
blQilx63mzGGJ6VbAE67O/kDkBu1N9KZBJkgKTESuHogKwFb5eO5Kc+ZCqH5
x7UHm3iyGW5XIixONadcjTyH/xdvo06N/rtLlbc8+Tm8y/mZcEo7nUDBP4zH
rqDjINpCfqt72itlBfJ4c/SRKSx9HQ02HhsbV9u23Eu6bskKtOlTos7RKqJn
MfLo+PWHUktCW99+KI8/vRXKln6drGqqQj+2yckeb7qrgclUAmrtlNGXO3P8
7IzncGv28D/mCVcSoK8n/TeeXaDe+VYwdKqzI4km//YbUZ8Fo5Z/B67fBPEq
ATw+NJyBjTJxbucex5DKIMaZazdQSkgECZogtx2QcFIGedKmH/XVpirMLZyO
3KItsv3V4x/mHmJX/0+i5K8C3bxBylw1MjDpKP3iFKSsn2xMoFbzA1uaCMXI
PteoMNb5zuHoD8RlJXiplza4ddxDuNdx2b874qE6NjotsrXnE09Li1N1IDgN
g2NG8SQ8puOxuX6Aiqs4dpzG1W66hu243B5oCtpryW+rvZhnjGH99bOIJ04V
l8dzlxXBQxWy5lhy8zx/T+aNegwZi/kB3BZYTF8kRTfl+Ys413+V/K4Na/tr
dlsYixH2aQucQvKrwNaLiZ/SeqIauKFDnLjWbQU0hA40NQduVRwPl/nTj8oN
xZ/DtxgUyotVeYDfEbUDR1iDW3tF3FTOgYtaEz8nZ4Vr3GNHZ8o1hLYlndxk
qLBl9OjRrl6vX6skoDmjYj+lRoDbQjwmW2IcL/qciiiutqxcoePpnOj8Qb3S
AlwfDcdRSJIGDgaDykY588bY9unzXx+96vYEcD8h1CFxfyjg2ydJ0y+/Poe3
xHLMPNCRnHefaxkJ265YLSBGIScff4NgUFfa+uo/njfvr6isytfMqM0MfNc1
QLoMe8LyQSNNXhcnmO6sO6PLVFj5ApmsXbIziyT3mIFoSKmuDAj6zr7ek3X8
Bb8hmp/6Sh6incn1qn6W/tOsEewrocTA4d2oQn/Ttc+cMhYmXcjxBIZK/qpo
QVzwDJbcYwEHR2PGle7EFKHVBcYwU1/AHiP19pwsx3yzGLexaba60rjCuKDD
PitDy3blyFSuPuO0iL48dpGl3zaHCmNSxdx/y85EPizMRcFW2iCPDL5kfrsO
bsOCTyn+0zRN7rxQK+G7GOxZmzQcWnNW7FeDqX5+HAB6fbcV3Q0+s4LfKPen
wqTDr7Ex2xagm122huC58whZCry6htqMetuZqARuSIKndQtNnHdWIqcE6uOJ
55SdTijekVx/rukN5V37SIElOkHr6j4vIB8uGluJTloPvdfbjdea8UAh0nnZ
WuHDOceHGgxg+C7OkMWtLEyZsh8eUQbOIAWOJrSY/EhHK6uyXzmO4whSj4/0
1fqAVc2kZ7oeLU6OBJKH2rrnAIRf3jd2a+vHbUnpFRjQ7qsXR/6zJD6lWEXO
79nMZ8w1Gu7uu82KCt4qBBeGaW5blX4FKjtbMmBow2zqSAP6bkmgYb2GN1BS
nzLarjBbOmJhF5jAMvi5ffgLhGlO0D+SaZK7dvgdUG+PRFQHeoli93UEeIDK
m3gMWoUwZPxi3mAIkWTb/pTh3SzwKOHWAxPhJB2QhNo7qGVwLyGmZ6XKIofy
dZTRX1nCOhacnDJgYyup+9IeUGCJa7Vh41P524A7DuMy1qK1YBkBGkowEBZk
7wiDFkJFINUl/UC4ShHAc6qQxgLMIWrXzcjASo8IRqMGKGnPFQwLTOz4zn2G
ih8EAKYbjnDW/GthvDO0mW4CuXUGegTPgFHTS7G19VXhhMKajqPUH7b0r/T5
0D1NMDKgsW3kZrO5Vue56fYMH7bj1bOuftW04McO+sGt5TYX1wyb7cYs3I74
/H1wUcx3ObMn20gnE/O6EXJPRyJZa2yRLxzLjOZbL2PV7E9pKlJ2+MOIHbeT
IZmD/M8ehENNPzaOuZ5sQlZaNsjcPiT4xkev2lWLYDx6OcLaD91+iizxceZ4
pW4ZuFN8Bc6Q4brV0fM6488T42p864Zd/vfcKBW3GfSr5mUuV7T/3/crNTw7
gPgmekjRelcgc2f91Gjr06ta3Y7p0bfX58U3mC7VZwa42+9ZzRfw7h3s5pL2
7a24jGRe4dymaPNTOkQlUXLYXQwWvctLm9B4MZy+1+tNWXcSNFIiE4KHdraB
orDQ11Fxxf7hd9diwmx2r2aG66y6q7QJp2ESDPiPWKdedyhFM119X4Rb5FVG
mwIETDJ+zycELbXSnTYCBz/IJHsLpxivljkxxgZboP341GMraGzR7/OvUqJP
L0zjYZ3ohnbUltcXochGS/mU8bt/48LXr6VohWhXFXmz65pOxS5Hci7T3lP4
q8D9UzGdRfO31C528NpPiC6a2QZIxXls5H7TQ/6U3KFq4lb4GpJ8k9y/p7mI
EiRmM48PFvFuGaj7HxUUhWvJ2VSotAhEShnYq6C4TiqnHRddWQj0iGst+Mek
FtM+y4AhldE+ncyxUT7QvR8q/DVpk9HKHy0hFgIT1BFQ1PSB5Emc31OuVzYg
aZLqm9qIKQ592h0Nycp7hJzb5F9cLw3LWTvbinw+pgBcTJ88Ch43XmhzN+QQ
p7w9j45tzEW5QpdJc++nNSiwoCJq6qvjEByEvcHtgoJ4MhIh/T0W2YlvtJcS
mfht7wpGJQFxSFKemj6TFHsNXA/FnJVe6NRbIFPR2wzacoLMe4QtjZ8Mntdb
o//PtPphXWkHEnJc0xaW5/pcOu2/DeyR7U6T9MDG7AVJN9ym5i2fezH8s0ZQ
in1/NCHoa1axZlwusazYd5u/i9HJwP8AOJjq6H5kBgL1d/bfQ4Xz/iNsNylA
m5LkbBblJTqcGRrmIdEW46Ljf69aXWxaOdIz8cY+SBYYE98i2GuRk6Gsmv+a
v4Zdgeoxk+a6LkHBY+vJQNHmpNe/IRSp0cvOtmnVEOdbCBbr1qnUZLy2y7Gs
uPfoDmcpAl5twNF0kZ8cULaWJFU8SxyqAV6T/Ee+X0iIVFbQQ3AdQ3l3QzZ6
fQGNNUZq6w1mZ/23kO6F1EeeoTP3ggMNhWgxtRAxmppRuMiWD6oBmAgF/WYc
WmHwDCPPWecBIX34axwLiqdHj3r2F/JbBisYWRqWCOqDTel8GYN0wTkYTVIi
0JfB/vhL+XjI2503e7AU2jY35184HGTFHDhZZOOaagZ2rhnEY32d4mBrhvPA
cqILqQUeUtG49wETAhjTXZAU+leRdoVc6sdqUjc/IGiymqou0osvuyHSrGqo
ojaiMcXuJ9B9LbJ/XVhV2CYJfMgg4Q8Aq+i6Fbqr7XRnAxUCAfHQvwoAU5X7
1GPIjqjyagGLejgHopRFa/mBsUQszWtDm/w5t+a7OqRH/oaUZPR7zJD04xsb
7gUz7sbYrbMvFCmR9NOlEs22kk47tPkHWI/2kI2doxBlF3SQD3dWsYMk2H8a
y9/VsBMxqEl6KbWCWZxzCvRnrPBFxahhZdpbn+/g44C2AOhW7LFgS63q3bbz
DUHK2+pVReqLMTaiLZinwUzgS90xadtvxAa4LExUlhn38EzVtipM/gmTp7h8
Pjs9bANWGg3WGK8scFNqQD8GQSzaEm1CnHFcDD2w+d96bfrTHTK4Qv/IyI8V
5CPJ6WThibTbnRRLZ3916nUxWNsSHgZBlWLojK0wWi+lZPd1meI12tmc0Frw
N73m6y0EcesDLUFcxFhr+qHUUwkoij5TWKnL4yCQ2SBeYz+DCWPNVr/nei8h
5NZ4XebsavpI9Pzk4wSgBLcPr6KHz2zh9lQBc91kJpk0moLePCIXbKlOeAkx
ZUE3UHOwJfBZn7bpX4iFAjLwndMYzY9jMLEsVs0b7ss4ffS89OTeCF+kG7UM
HejfmVu7iEdvYGgZ+EO998Say4yjWeixMVGYwdeLeP5nsj+bQXM03h7RKzbG
rraXcZokqH9za1x1ERQqmZWRE6PYD+EIJF8SlP95/+fPNsFsaYxNQ6l64Lcb
o+FY/PjlUwIEabTT/GWDOubAVPY8vpU9falxbpq/PF1eIRAgCwehDCuNFDrU
IISxOWDabUpyuy2mVUkv8IJF5PTZAIYMKrlSuyyqr2KHwfbDiZ79pD3UPGcK
2EfwGck85ACuc74lZR8m5kbfpZZm11VCSN+x0EEw9NBN1l1ZgQxbbHKVsJEu
5t52vAofBVQTp6dYEVRq/vOnR6eEQ2t52Yo/FjW+wIoLQgeFw2rBz06pBx16
D4IxE6be/CbIGnEZ5uuDtZhtADRvutoB7sBDx5tkXX7hcAaW2JVdvUJLzTuL
a+m1e5l53Xmx8QEcPTHQw85fCdk9zHbrd2YIKlOlaqIrVUBt2XnDD5M+rk/M
7/bOv8PJt1dWELseFViXLCtMSDhjr/erNMA+Dtz+Y9UIqRtPtllMziDSA+DQ
3l1DCY90LJEEVbwLzBjNyhfuVCMYd+B73mljwFigyj7g7vzAeiM7LdDbv+qB
7XlcidTLJGRQFMhq69Sxr26vpezPcmWfIMzjcodojWMeEml1psyLDBfZWdva
9zaFYAvu7a4aPr8XbU5lym0WqB1BvEFJb1x6YHYv0fIQb/GpJM4UjPYob1hs
B6dB7mmtZxU1Mu03Ln1MfzzrdmNnjPmeiDJItdoxfcNfBKybFcACsdHxuSNm
bg2x58NFqvqHw/IOvPgWZCQIbzSxgJFNpihuvEcL+5O1gHI9itedc75Dti/l
U41avBR+bkyuvxJ6uxJaB9aMy/AEN7q4Oe4fOFzRDU+tsH71LsdI76M9CsjX
c7F8nbZY7zmy87/lXNwX6dsES+vjnCgBIOK7qOSi+RC0SC4WKEJWDvNjnmNv
uQRySwlM+fwP7hDgQc1oX3EadSC0ychgZdfLKq6fY42YPhKS2IRImi7ZJUQt
dQOAd7BJtx2ckJE0fw3K6VqR/1oVZRtLfj5hus4OuRc9kZvgab9uDFREyNs8
j97kLJsMvzRT7BNoNICiKW+n99Gb1HKPTfxErh2EVkLbkZSQuXQlZiGJva1+
xh9lmdaR1TlZkHdvhnL5pTSspnf9wES8zjaKlHkhKAi/YnhxZzoQ9Q5HCb8h
9KAExDL5BK+wiyoTxvsQ06B+/KgH1jRsJs1gVS6XgfPw4m2/mOfao0Gia+bN
MNR3GaEjE2QQ04Lzeuk9UEdYKOkmesVScHh6rjtY2kLpXoGdN18b+RA/UGZ1
1YH/pRYs8OwiqzkioXFWlu1rwEnuF5SYT63oFBeX+p27ALANHjYlUeyFjxbJ
zQSDcAIFkuItHjS9aW/nqZMLvbIwUsVs/uvucTaJv5Oj0GOcKm69SRBBYpXG
5pGx5KhlAmYuLeeQh4GMPFYqvgyQstpO/a34RtMMRQeu76R6/bRiSE7/Vbhu
OgjYoYAWNTgMsSgCmWDrj/nwAiDL8hYaAHZJijKd2k+r+V/LWx+rYZgZj/n4
5S2cwgBYZeCIXJHXIJlHOa9o95mQdUGBDaTWO1AaKzIRsRdqi5xe4YD/Ihgz
N1W+g2waZAwWk0lDMBgtStXWYIneV+haA1fq7W4XEk2V6Zr7Njx3Pj3AsIgs
Jw821AdtKNN8ie22MAPkxGnGhMczFG3UMwduElmOjh6VqC1xvoHNU3ikSnYT
H8bsEvz7l7w9q5iTyTz2vFq30qhAoG0B/AXY4jFjoxE9td+sAE8sdFyIIBoG
gD6/lYXZBr7odaCfLU7Bd6+/KSuHm5iHoJDyenHSeMRm6DxiD5nNcQPM7unY
2ldHpKIHZ/SXsieY/u4AoF84qK6fcuD6hL14lucgnS9tLR1gFakCvA7zXzlt
2dhe6VAp2DpmR0n1K2oQIZC93yPvZtpG2o52BdNjTPeufY+UNm60qQceZp/b
3p8vI0uz+s0yHwYWL2nbCCBAwWx61SugblqOiZOtzNh2LeJICmvV2thtduWE
9+aEeJhLEfdvjzR0YDN+m7Hpwntqpg27OjEGSno53xyJH5z5OU+DmMPjSFUK
ID1kog+aasUWucdhYr4gZlczuQw1qgajYzgNHEJ725q+5ZuMqsxqX3T0tqjC
3TigILIeeZwORxVG3AxUjA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1KMEgbR0QOTQlP+ZjcXuDPZWLJeX9bPjxCcZZcqC/5eiDMWIYkFPhcAxUE2dNtWXmiXKmXOsLXBHa9KpivoVtuS4QiOQdK5O/MORe0sEGBc1FbkS3+P0bLSrbna7fipOBBYkwhq6G2S0GxUClniw5NoP2NHZg+ICM+kfV4efrQEGOoeTxHjrta1DFcgDpF4vqzlSiXE0Anx0ILis6ShZ6tiNhEXDttAoLCZP5VFz7qNV4sApr08OUrZ8858L9hyIdxPBLdUdBzIUj/cCHebpNp5NEJQLdU6vA6GRKulFk9sux7HJ80Ar//BT1n5F/kgyTmOGyLaftQLW6pSnHpagMHk1nwVgJvUUmPAlYE1w05GG8ogtfSu70FiuP1e+Z/jdvs67y1PuVQqAkfiTMLnBM6zftjEAIfPOkFRPo/CV4G7SFFjygcDYY+PigL+uKcfENROsoOqGrzCfLh2+yE78NT3TlPsEXeC35rsOPhMPqNhZ+5jwhHY/lw9LdngRNEIgGgLH8hRi8rrAAHLZjO/RaGkxptCS5LKZzaSuJIcrkudGcL4oyjlnz9bVrwBZWSRWth8G6opxT4rdnQB/I2w+CSOVz39QhqAXYT3fdlONzvtuav8PiC/6dIYan6Msbltc/vuZ5qFb9mxI5GSlXV7HvIc8l/xf4TPDCZAsM5lMhZkgeDRPZN02X4KBUfA/5PO9rnjnUrdZKnLvcWkEpogikLjisCSfMR6/KKlXtuWOcHUBoRKlnj80xP6F0EuwZJMPYUhLI5kRdslxgTgqdMwUUCJ"
`endif