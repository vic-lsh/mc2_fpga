// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NDlchjcmtxcQVwnR6DaxOKdaZI3MhSX2m4djTjDlRepptscCQN+tL65px2GA
Ro92D0V0QQTNwraSJkuiPMH4OvdYPH3bsRE03atOlrGoDbyr45RE/c0Qivl0
LhSj9IdiMJ0CH6e4IspOOrtAB8KKjoraApmz70odGG++FEVsOxQ72uIx7WXO
4jDF7MVX7YarwsV3UV9SJXSB6m5Vbrh9KpAUm+BwJWN3R/XshqgmmyWbHdtD
gdZZ2Yyhb77j9TOajcUs6CgqNj27qPswegNbb+ppXcWQWzQs2L2hIWPk1zyx
IwtINu//vnldKRNbSOzxnC2Cu16c4M6l0GvtsbwWYQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Y2/d+gAVVPjiO5C96KUvYWRJdPwah7HhykcnJAqyZ5Pz5LiQfhxUiHxLJip+
vVJng5Tm4mnqsdengQU9y0pQ6DbEx2SUvz0PYLnU+rhqL6uvNwxSCUoj9JAp
s6q5fMlcam7MILKDBjGqrwPFGK0br6UY0luTzuPMWxBgi8/TF00X1RDZu1Jy
UJSot1CA48lrXtaFP9Foo+9rxglVcvSVZuip2sUn0I++ZskRzBCkeGz3F8Qt
7YB4N4Pa7I6yb1LXNx6C9eFABgXMK8bnE4IFx6XwTfj+D0Rma0jgeCuMEbqu
ETAN5XOcm7wVkCpHsAvxNo0PWMzSc+S4f9mHF5uKbQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
L8gu5lay7jTmK2yTm6RG946i+xAQnpevaQ83k8CdJ3DINVWKu2EgCY0Q3+h3
3oXRLk8PsOCrMLtNFhhpYHQAHT0/vJlsT8cNwoMIe6q/rPkyFLLWPnuV8fXr
Z58TeiMiko5Ww6uZa5AnbokU/j4Qy/rKormmWkZOKJeMgz/X18rBcmuZdPE3
l7qxkilvRctMgbieeML+9zRsogiL6XqKaWit/sa9mfPeac6iWxw0I0MOUV3w
C/4B/OIs1GVqOfS3sxdN429tzSfG1faU9S1ZGYc8fCVE8E9FvaNeQR/GYFvw
/ZU1JIudg7JctMf1u3sQsEcvUKBjRPemEJzXE1iTSw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CV7oro0VjBOyWI8gacEs/0a9lUcYn+SRbDlFTZI6a6StHrzqEJJPlbXZbZf9
zyClnbaCfNUB/kP25wmB18zGebFyMTtDjuZAjc5JomjEoJnI4WDWazX/zQdS
dOk0wdMvZ4dAhomzQxDk+r9zSXtCKuzd8Pzgtx/CNlfqy3iucJQGhj7z7g8j
MxjMV/6RaXekl8yYJHHTtSE0St7ehOCQzmHhvTDdpxKXUncJAbJNPzlRFMcj
T3M5TRKXDYNXiyyRxMJXWiB0RLUiDLLSotTJgJv4GyXRFHQ2/lXV402KOaZU
wBxb+pvBpVUB2vAyDo3ehtWm7i3V2jGGqh8ohQb4Ow==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lGQ7fvOmoS0K641hqVq9NU7oZUJoJJod8b2nCNFVdUv9bm0pNWyRPx0DtvZI
rS/szEW1G3+z7EkVeDGvSR9I2M4CFMoEyXGum48ZFVo0VAl8QY+6ckDG+rT1
l4Hx4HI7B2/aYIbKBZWFku1B0LSwTCpD1dKGYbrEHobBS/LONQg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
xdP0jy6TE4FzNLHmSnzsdJXunhqxE2pDofAY3cb+fhbjWQZ9s0fY0/gKon9k
ElwsnnAmDTV4UgbgA7n1KUDgGnDi+xZLr3hX3xTclG7zopK+MtmVP2oTQHEd
txPSfXLhli02lK6dTF902hbVhFDS4qYaOcHVwqX2p5EnIMq0YbRjy39m+4cI
UbhiQMKFCkv0HEJuZn6Vro7J9T7fiCyMyp2SMRG54+02XJVqLcz6ofaxCLPp
2DeinCpJyNmVBo53i0UOU9WCdt5EBnhEqWHrd1PetW2fxuAIuCYbWWurj4EC
fxoZwzTgAMjtFzXRjxHoo+GnJOAZQBd3LnhYproiYxEzWjhktLOcQ92jnpsx
2fnLhhiJFPqOBUdmrhgfZIqLwuV2qTYBfZZzFGn/S1BtgpO8sqJNi2ab4odF
bjxOiMa0Tonmn0IOwQldkZEAp2/e04rZUoU6JzRAmnZAJXM2JuwJdEPKL8vn
NQu57N2nby8g6KhefTRwFxBr83GuGOHk


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IgSvjCyMsFCQ1HmUqOxtQtGx+5HVfm2DtgQw1AutYIJLMTp1RhyLaSbLxmcg
rApPIA4zjvE311pRvmIZuSJTJSK8nmHqsceNBVjYL5lxAiGJYQtwzEC5tpaO
FXcwW5SQnbAzQ+P1Jxc130tHt9B/hsNrwCp2Ra7qIu5Amqovdc0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OF1VbMP3Zp+mDaycT8Bw+OungDIFvPgFJpN1yYeTcn9Yd5qrvZlXXsCgwMEg
M3S/eKd1NNH34MCUPvkiimQPnDNFSB7+PurMgDy8zNMryluZiz4qXW0tJKcj
ivw9ElVxX/sxdac0DJlCR5p5YHdLQvn9GMtYt/TFBbipt8FmQTw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3120)
`pragma protect data_block
HYyxJL9mrQJgKPqp3vCUqNem2hlvtO3Qd9hohjEwjiyrgr2zMZ24b3nbL3W6
3vILpEGKEIZHW3NzX+T3o8jhWw3mtOTNL3vwQkLE3r9kNOSHb3WNzU4pdxTe
RHM3eZ+V54E94SfAXYY14Qc9GL2DJuUUi0zKHONvmEFhnOCa6hnnwXxvC6pi
SLK4/+6Utj0HswRxcJRqvmqapgB1GwWc1x852BxpmkjrUVxt3Vi8sedDj9Z/
LaRYSizZaJyDLcSNaMYtJx/nJ4Azv3xTrpnxqeJ3CaivLJ85xqqUWOF0ddI8
3szTScXAXjGm4rP64z0xPcAVYqMpnKImmMnG32TYBSJgCrxbr4g+zvWQ2ag1
AHKPdiIafXm25kBn77BTsI8SRaePsKu0Em6VSfLdwZzmP5FpN1hIiVgd29yw
NXb0HmYRCIWV4eJ2wmvHOh43X/5x1X4BaBO8e8DcU7lYgbrLCGhp0AVJ4TTd
4W+hki0wYJArs67fDOvJv8Yk7TcLv4/yfQlG/cz0M6vwGlHvZ+907jkO5RJU
k+Bq9AL3mviOydp4MQdxXjEY+gZpWYSFLhuwun15Jo/VbeoI8R5va1OwbkC/
STa91eF00s1JjIGRoaIoXnaR7aH+6FaKNMU/JBDsLC2pDP6gKeDU9XWkHIiy
TZG+kmX4VqLTVTUjNxYU2DQnRTIM1oAhNXTIO1W6RzKmrEmX7EC/qQbfI8Ol
BACiFCjx7M47k0tHxINrVejcCERL5H1o71UDNLNp5IFyUbmdj2yONeVR+BSY
puCDN7Iy+ADys/zc8G/d+KPPuFzA34XqlUf4WemGgLKDkyEre0Z5CNOudA8r
Hm5DaIt3NnYC8LbrA//LY+SmJ1VjvZM8dCBCA5bMBa8CDtPU04pdLqEc4rNU
nCTaBggqM63ybf4BNkrV2hJF2kz8F+y+iyBVFEioP+fqyN2cZADbaMdafGCP
NFKB9MeMppuyPK2IXF8QVGxf8aih5POctV/7GL6coY+OcjpNr7mPDpiUMtHN
lxmy3aI7A7B59ecUs1xZkSIEdKN6YBp312iLPPpoO6CIDZSlq3yS0pTnzUCJ
xWjQvCLn8Ejqbr6i/3zpC42RC10EQ76cHnpo8AMyBKgr7nRkMv9V2flbXrDw
32R7Fno63tUyfT65OuDIgECieeMQycE+XiJCYlDv8IpaaskmAfumHLchrSU1
0SY8TsErObipH4aoGZXCEoY1SWRic5uIFUsysijtC1qi5DxSyvErUcEADq7D
uJ5JrqDoktUOFI4UwbHs/kPTpjUCbTrhmtPpRvCFEBvNgugrTUsyDJxb4ZNt
Y57xFJYYunE8Wxv1V1QHWRejOkmi/uveH68W8Lu8y/xQnqRKMM6Kv1IXWAV+
y3njXTf8qgYobOsueI3hO9qDySozHPRwJiGaej0AkinDJ+6/FG4LPymGo/bc
bLlWO+hVknh7jyvLN557rYXQY5zEqnUZ48nk1xCaOOeaFhK7HO2ffs2CZGAy
PvdaztRY1KE6WkXPMZke2oFy04lPqcxDTGEhrZs4DgbvPakb0VfW2u0GFa5i
0cGBcu/xyekJFqHDI2IUy5i18sM5BJIbk/70dNKDxdnhPNO9v6huNoRoxucV
3+VaHV01m7ChVxQq/t473K12KtAtGe1P5QXeDg59Hoc++zMvEGkzopgyiwYw
ygWPCS3ph9dmfOfp9WcMLeShTv04zbpMZ37TAOngk4EuzE0fhIOOBOJN/53O
JoNDHU6KEmtXNcOCI159m1lTtLzSBypXmYR9qPzA2KXpZr4TC0+/N5GKCEU7
SKrM82txbzZOQxqG0oJ7OqNICxiTbDiDoiJUIXOMXZDq9lqQdPcX5PTUOH4s
alSsEb7IUBuWvgkRPCw9Bv5weSG97SVsqeTrRnh/rH8os94YilKpSFhnSgBG
j9OjxiGBEPeyes7nBIgM2N7AxlLQ+huRMDWG5r1g3YqZWf3OH2Knxv4vh4LJ
smoTbnhdJhaLfphY0knSrogYl8TkizLiM/QOCXjImbmmaIprXuBY8XhdioSk
lfmn3FOk9ew6Q8SiTzvagp9S+5THgywEIjToBkuIM/J2xVxo1aM3+dogn5Qk
QjohJgqjeaXWX1sK2zZKhbM2O+XDjoisKsShsFCf1o8/n7OBnPJ6kYQabys2
IiOKcuzJETUtip6YJLpmWE4ZqB9CETa2FlBDfAuIt6Bko7GLuOVVwNCZIwEB
0K4FXDbhyKIhDVKjEw2o/2weBIFYcfkZmOTY0QafE+Nq1/+0TwMDfISl2KVP
123XedMhnmnVQVBz8Hy3v+p+e6Brq3/RAFhYXi1PxU3GiG6/IWvuv4e906+1
IV5Rb72rtTiocDGESDAk4Vo8jTwY7eVLFsLsg6+kv+5cUTmJkvhPRZMIQ5Fn
eXZUjSZ0X8UxE/0zrpZ/JFlqIy3chTs1ygLM3MBz87S+7FYgR9vCAbK/pEMR
wGmAZvkXseRGZvxWg0o274q0SrVCyIt2UlXNwuBERgaehWSWcOz1AWZQ+eFm
3Jd6Dl0nRdaOicWKJNkqNG06/cOUQF+93IGO8DwlV+zEa4geKHuMQGG+zc+W
NR2H1lWi8KaU55HzdLnhEbwca7qa/TWiAFIdLdlQK0oNthi+KzHDwO+vVtgi
cNo1uBEYWPze2u0FvNH52Ikpt1k37acrqtGZAGKAW8dqJ2Kf4vhDkjHvjN2s
HbvDKtrMtK7NhOV0oF7L06a0geM4OIZ+1pxGR/8dD1lWwogB5agsSQKr0eqB
u/Uvtz6fb0+xsuZlZBxqm+zaMuU78wLXOb/pnKtNseKQMc6mlmbSyGrJYb68
SIm2Ekoh8LLnD27uFxDl47PoL3/044/Y2//KZ8E7UNRecJuPLTdVEapSWBwB
hfLw0SCUFOIqppG9Xm4Ee9AAhJMyQcmU3D71HSw7VMFOZZmG5SkVm2xH9uc0
IzX2/mKw7doQJbPlqx+gYy4kZ5nHWEbNG364S4X0WCguxQ0lyWagXbZsS25y
qVmgojbqRQaKilIebIHamNBzunV9OVaA6t0NB572miQ7g2Ws61bLSexG4vbV
iLoYtO1ExfIoq3rAshz+/Bpvj9xovTf9H6muiZ2pHX8QZziJJnahm7bPYi+j
ZSw/1bhHXiPdMhory65tpbJ1gtCjTHVJQf5yaQKFPLuY8IFitJ/ADsgR67sK
0tVdsN57dBxkfmBLnXkZXLrkz64FP2f0MqeHFSlA+nOhB/YO6681K9HUA9cZ
EIGl9TZKSe9gdUWQPtlbkvGT4ZVP7Y1FJf7b2wn/DmvNHxC0l4Bc+u39Wm3D
R6k/moXwpwHE/gLqM6eqUU4SPBnOCLog+87iU3x2Ql0XjGC4IXOhqV9D/uG2
ZpuFoMVNHnOnYGzm4J0PwZqFG1tczKmCTfLTbZRkxkOB8M+tqKTj6yPwE04N
UbdooPefFQVRJiHrvrMGgsMwICAU67QAFKJ4hflZepz3lgEGtg+TxiCKYVXo
h0KG7g4fzxtb1lMZddDLFUQlAc7IygsPHd3gL6yIHimEV/VcXGd8UXCidhch
MDijKKPtldCphQ7u+ml62HiDz3RC1lO2M3zQBk2GtrZegKJduJqxx9JA0qo6
EdVft2ShJJAtKTET+O14Qzfy2lYWJpoLtHMkX9z/asQO9CfINgsNPpGWpwlc
nHVx7U07Q6mke3sMuUPXE/v6fnmRqVtkzrd+lBu+Q+vVLV3nIR/KtiEc74Y3
zweBfJ7NQGGMjqL1Tm1iyHjCVW86Ger0FkT+iU0RGD9Fk4K33N72KQf9CQYD
NeIZNaaj0T/t2B2ZvqgQemaw8af0wX3uw84WDpaGe2N6+0ASTTLUVPIJATC1
Ys0K6UW2NmT73iK6eQZtP3WvV0mZLjnepAvmaMmY6aXSn/5MvGTGMsr5Ks/K
9wYrtLl72cb25u31iDodWPE1KvFBOs+NmDv4jJh5xgFyEsy7lhQyQMGvrV1m
LC/JLgVEY1Xk1RP7fHh59F4ws46O+fDpQK7iPFuFPXSzNv9FrWsiA/lABzR1
A0p3Eh8AZPeMJB6/+AMbh/cwhVtCzRPKmVexAWFd35Ea4suDpHCcGITjPKJS
dq18xYB++A/a8JuBS4O4eNmKC/2gEMnhxIxAHX2ZKFrkpHTquGwZHWpPvG6h
x2uaDtUpPTcmJd5Q+aNw

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "zt4TNE+YtmLl37OYNCE/66NMR/xqvkEg1QlSZ3mTK2MFNyfkI62wSpS2QZeThlgCnIYR1zhT7IjvJUYLeyuAIzCodGsF1F4ZxCIp5yypQLh7UEeTMkrUT88kUYosUZjSFKaBxSCMovVfYU2U0shTMrceSLHQpG35ClzOr+1S0gn2Lgkw0w9sDPCoTvCeKBS5A65gi4Rr+xXpbnn3+lWl81L3Roc3JZXoB2wRcPRdRzfnR4hwWADv2/N28aJKDgFSHQG8GZZYB92aMNPft3RjCml25INEYTZjlwwKiaX1cYO/ZnE3uENdS5A+M3QMt89Doi+TDrirCc6IE1tHqM/B6uUeHTect3UfLfeDF+raNYvqq5+auszFvbXElN/jEoWpPLBvtymY0uTbVDStRBwk3Yv303dYM4jCTYjXpFbQ/LvRMCmgD7sBsB4FExvE60nJneOIQ7AqV75fb7wySuzhGR4q78S8a2erOTLiEKOxqgnkE26qhoQDsYfbDBv8BIj3WQuiX0ECHLsVDoxz4v3BWCkl6Uv2Uk527x3eDWzF1Z4x5fUeIpa3FshjmaqGjIaPN0rFYri971ZgN1AeOoSo/fWkOvWB5x/nppfw3bAgoP0/XgnUmjxkZfKQTz/PY8w1c1AXmp7/i/RLtFHGk8GshsGR/Ycd/RuX2++/jjxahTQ5143Qu2g2GEXDLBWTHEbn6m4nBJzQHrpZtmdlm/4Miq29JCrFayHRTp9I/Bo9ufBMdx0H8CoTFUhbzKe7TlyAgT/RuGUvLL0NnxgNmiWPyeTX5iO6Q5HhDiPHCkvgLy0mBbjPG4aNmELsR8R2H1rzFoB9p6fpJONXmk2JSxxga2g2ExQXh0WbRCeMNzoeMfoc3YqCZ76TuqTLoKkc/ILqU1+WXRlDg4NyR5pL7AA0OwDlD9XGiauOvQhKOMnuzmkzd0Zk60NrvHgo3P5bRTdM0sOTBV6P+QFzbf/rvkGje4LdCGbhokWQoFLJ4iSKqzbK1BPmuf6Ag7uxQqm8iM4M"
`endif