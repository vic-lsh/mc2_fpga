// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LB/pbE51DfGdir1z1uhxji3BGglQjVmOBEsl1KxmKdWmcw/dBM4UM/AELZH9
8f8OnqZy3kd1nDRe9qpqyl/Nvb47b3rzuBbhT8P8ladP2u5+DXhj0AgnAIWu
HPu+IahP4Q2Ado1OtKJnK76MnbSHhONFYcWnR0CHtgVSLRzyczR1Mh3PCoaQ
Y4E1RJI5PlQOtG+IE9XcLZ510kI/Ix7wTwq69JhCAYmS0gMiJsPqzC5SMeu1
U9JRTdPydSGmeOsy36ZtO1+sUYwPgnx1K9EXH+z19QvlljuDJL39GrRZ+ro/
4pEv21zazu6WUiuerHA+2b5xT4bB/xFn+1mWr69XUw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AvIyQ2Xosmm4mteWYHYQGdqSwpmNM04f1lrfeHLHU5xYxSNBZeHbjq7387ry
zQBEmItTgnzGY9Uz2ClocrYQAHeAACCuIZqDyT9sQclhJuE+Ma4Jrg5hYFld
zFgj0WAs2njIhNCvI5RDVJSQMLgehmyDjGoV7EvrJEp5uuii0OZ54T7ohQbf
qmfaRmQv9IRtztkfVPD3SjyZGN16MSPXF/m4vALhBHNEa0Mg87QFMiM21e7R
7VqfOGsLbsjofA/HThl778x+Lph+UrphO9NubBBjzzaPNVbCGvKPVpPKVIsu
EybgzqPQWaF9LJGwRB5U87NZDDyQtiU5tPApYs2Hsw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Njbobjq+MHN7ZDFuB5MGNoCro8M63P82lS6PY8nSQOTxZL4FGLOkyUTii6iT
81sx0qyrvH6g6yOtXOVG5g5O/qIiMfvpqSqd3+UGq+gftlaYW/FsQfNWFItZ
Tk8iMgVR+mVQHOngmqB2VjBp0juAkesOZgG2zRI70Z5Ez/IADNtSoarc119m
xFP6H2rcjBCaJtGV+B/20e1xAPhr/7pWpzHVj45vCILsbq1RCUQkEK8X5qJl
J6gf3K4cIi02d2U5byuF7YuR/jWuZ2C+bPZVEevrExi72gG3VF33cjoTYkJp
l9bYzI6FfHvom2JhvMnW5uU/Qv9QvcXdpGxnXEJkKw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
om8hkwimafllP05hWLhkrrkVslagS6niKnwlP6QCXN6u6usqHlvXJjB5Pm5u
Mr+XhinIpg+mvC+7flyw6P701OLQbEHjcDGfyTr1oR6OM+la+AIX7Wu8Znw3
3+cupby9klSWEy9BAiw9l+CxoolIiSUOHx1AxpziQY9WVb6I7JzLIeesrxzb
bYTT3e0RoeJQ32ady4zSGAdjbPX3oVpGok+8IDQptqnVmIMasP+MNp/427HH
MA6zTgDr1oFVK2xLB2QaPfRH+KgUX6IM4ONzSv7ciZDYH30eIh9Mv5CLwp0w
DmQ0fGkQ9ow33SqOe7IqWaLddOA9ygJcy7xDRB1DbQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qRhxY4hM2BWbDJjEg95on1G3Gj4NnYbRUx7xAN1ORl0F77gh8ceK2+c5oBGe
p8TSt3DfSqMUqpjJ0KUXtaU5emek81zCePAb5Pb5kxEtP7vI9xfLTt4b4pKR
dRi8u1PfaFobTO1sJwqlr4FKxE/1iSXz/NbQE5+qYhz4s8eSNlI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ZrKwQXC1O8F/BbkDnBUpWFMzBy7jTlLUFBw2HA2hnY2NGZX5E56dXqFUWP+/
Ousfjobm2Fs1JvKveySeMuBfrLkDo63z0PNT7R8t1swnoV50TTd+/ckW9TEA
1gF5qGpTQ+taWSg1Q00p7W/nSLHqxpl9GTfZqR59V4OkoDVWfapcOp2Z8uKc
9wIJ5bPM80j8VJJXkZX9WBG+R2iMW1klQGWxFf/KsdfFCDTFMzbAW4CEnBi6
BzDwyQdC7G98N8qi+OpbcHdiDPjMMfl0MFjXU3PGJaEsLj3N7lYFRV3X59Ue
+fVOfsC9doRGqVd3oO03bvE1HqFdTJkf4qR4aSn2QHu2PZdvP2//PCkN9vIX
KTvZRDGM63ML3n4LGQIcWN+5gNHAytlAjOTQ0HLlb0j6J13CprAW7ehdbtOp
kmvO4VEs71LZqkrZLqLu7qgw5k4mpLt+mL2l3If1iFvSO/rWGDpuq1CWaJ4C
S+y4wQm3CIEAyZVzRpAUyZ6PIRrFFD3X


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PvweqvbR400Vsdln7VIOMkh9ZnN9Xv86H1nHXbo85UWnL++Ly5x5BwFJztz6
b62wIFV1UK27/2lrSQ+Y5KXtKCFQ/vkoc9fcP4kK/w92uBI7yUKEn7Vrd4qw
YCFkazPu6nWb8yeg5XfSYkrUV56bLM4hwFcs8dzdTOoWZpc1cvI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
F3HCPpDXhGICWNZXgiCN/CTSMcn38KWZ2mAvYRtF+ueW3pWUteyG9yvAlC5O
pbFsJkUajrU5KDrNHifmeeU/8RRU+mZeY4+qi/DVD9nqafvArleo6VWE1ceV
MeZzkEQEqMoLSDv8dLXsoNXWyEWZ6rhRZPyiVzXMlhYFPS5zC0Y=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 420368)
`pragma protect data_block
R98KzPjXoXBCXKrp7jDGYXWYQWtLTUjR6jYOOulGcJrxFNRdCzjq2RKjqaZD
xj46yMIGanDJ84cA2ledAjB9Rr7sMG1FbwNC8N/ln0djHHWzxwEKpnlV9zrY
j0HLLieFnHALIM2zwr5UBYPsAmSlWGMIfzlNa3pU6rNWkL4xG21mFblCgFpV
2ANsPq0IvUFs6UOpkItKuPJvzURvXmkWC8MtgTbkkD2xXinmkBV7PkTOZcrK
YNO7Vj18I50kHVkiTbe92rYqPlsjzKx+3LpaWtuE1FuzSmByRlz/1XTEx5Zl
ETp38vLkdffs23ps1MHiTCjMLk+oYa1Wu0BDd095xl2EuMmZm1p6yDqzzjtx
NLFq5qmEIt4WEYq4FCzmKD71sb6iKKK3Us6eBc6aHn47dPxLpr7VEGHlXq2K
AlQPodsgJHW857G3U7eAquINlElRdf2cjJbLtX70rdpkM6Ukjxf1wA79v5Mr
/t7j1GnUhqx/HEUNB1nrem802rvm4cBOJtr2X3qF0Xyp5ijNCkaTiowQY/D3
bI8WHG5sb2AxorURMB/on6CZrVKBsjrJbYdKx4FD4u8tb2kZOx+7CyZF+qnZ
wUcRHHpQdlJ0OgQOFzAVuxj06ri5yF09DrGusvre4PgBQDBAo6gKEGyJPiHE
tkS+fe+ORxpKqG/3Jp2cf5Hs1Gy/dmsXTFEH5PpQfsQL66OyiiSM8dbFgqnp
FpmOJfwPe0hxUzIP4U7YoL2Y+ShcDHDGEkFG07BukWhqYX+mPLNwTd3UOFW0
c/rt9SEvOe/0F/AcPJW0TpKdO6UoNtbjqHLtZFwR5npa+ITBcI3hbmVa5TpM
QF9IgSuj6Reza5oAYncednIw40ALqgwqFoYx4US8h3o1GA7GRxf7U/duvuZH
yjK+FDsjYGPLIRD3yoFFVo6ZOnWb1RdJELfa5nOqLJjzkXU/IwR2ehiQLHm1
HznVqvwxQsMslLmCyDPV0c3QYkL+fBX65jIZGmdpu0n7O43TKvQlU91XbMlw
nDnpdWJRuUpzUiPKEFuo33nVWDSb1PRrTg01nZpaPHCe4Q07YQXFXrr+Zy2Z
nzR5wuUckN1K80wrA7k7w+c3Y1Is029up7fgkrGo9em8Y88eLSxDAOrk25Ij
GWVzujPTSccZ7PLndKT0x2EVubPFIuXLLOw3meUI6NeDlhNMXh49Vn5DdXw4
l5jXqVYk7tFqiJIayIzWd3JQ37h3kC1B5WW6OvBj/TRLgTuM9LY4mhHQ7LbC
47A2IrTYHtVDWqSGiMDVbbbAGeMKzyYDRL51AhZFmAt9P5mSFL+As3rgarKY
SsANtmdqt+vSBJfZLEOxOhl8YLeMwm5BSeC4yUh/PcmApt1Ms9sGzXFcvZlu
sjZIJqhtNKI+DnSEYrVwqu4gsR0VOemYCnQxRw06+arBknn4DtVAoa/Jy1lQ
E6oJFv8YM6jWWmBcsxgq1jZKReAkWsyqdf0kXPNaVz0LquzdLQR9YJ8rlndf
82MqVUBYKQqSFz8jlUgJc6BVoMoNoHdId5iqxAB3FkZG9o4dzt5TAcK/NeXB
uQH/WZJ8EAdHzM0PfdEj+8FxiC8XB/MPSXJWFsJbZqTMg8RTj3ZzUI6u7jfz
KpG13YXcKGAV1MUYoCfuZ4+pmNXwVxvmGebwPGUj62AunpwZGU2LoYXQnYO7
6htXm/xF7mD1gnzkWmKsICA/svImoAEhHi696D0UgzVmxj6rkaeq+v3siCYf
PertFpsPpWfJ9B4cM0+b4G3kTuUDxgi0BGAN41ByJLCR6rIRN9vw8uQztAVo
hYIc6TS49dPgCXqbYjL/bV2bwJyP0PPCJjZrBwy+Gd4NRD1JhyScMX2N9+qo
+u6aMM6LipZrtzZuWoW2JqiAPRs0b6RC0tXLdlA6OOA9GR0JgIakZ2Z/qBqj
Z1XjN2ud/bJgo0Tmy5Olor20ZkqWxsHWopnH20DZR6JWauRb2uGx8vRmfaNm
lo8RmEWHH3qUe3cwOWcFEal0ZbE7cWfa0JgbBYnAPA/vDUaBp5tJino3X+C1
VY84496DMIZNVIK+Pq6pG5R4ejailMAJc5VP38Gc1rEXWAJpusZVtwXk/Qm0
FK5WH6+jjYbrozhLsmV09l/YYfQVREM/yWqd7i4zioAdiyBi0p2uvcjLk64X
3Z31CiV2d6VEcdqEacbH86bwMEbxMFECSCeyy91ynRNo05b6NJ6Kw6iqQ/rk
Zs0abnN6tzO7Wigm+8B2v/Ax7YDLk6U/C5K56UuLhO7MvtuqBLr1uH2GuQva
TSW2s1zmAgRmUwdWb5ykemufsL/SksIKN0hfcKmYF+V+DCpQSxra7Np1nf9R
F5TBSB/RvLBkYjML+Fliv4lYajn8s7pYl1C+ZYyIMqqMRgwyXPKSZKAQ8kPJ
iH3boOTjKzazxztPXCAWumlJpgPqYbO04elnHn522DPj+68siBZ+4dRko/q6
uKZiU1Q+c4BZUUNcvj86dwaDyA86q3OIvxiE2yLs5k58PJdimzsJ938FMme1
RDpAV6a2wQ/9+GA7YTFcZkNrrhzqzK0YdhP8oI+heaId6oRWgGrFif+VbjYu
pVoIK8/DbdUPB+4DT13tdisRvT9MKfzCpUE6Wj44NkX/gZJIK7DFXAw/tHL4
PzKx3D6AeVBezkGRiEthHdvpEBUzr95p2LC6yQlHa+y4dR3G67xYrEUSTYL4
tWiVAMRXvf+MmFAlSaLa8p9fMqKHO4UtI3lgRs3VSwDU+fGRAth/I3z1ateL
Pgs9P3psDrClmfx7+bqG3B9YwyRJkDd8z8w+7zPz8+n8GnQMMjVMxSK61my3
NwW4MFQwHdjL+YYpJEwPB0wTmw0t/rYm4thjiGjKM0kwh3A9in2laa5ngaLB
yzuoneAs7R4t/wZsVHcc/mnyW6vJ8fzybMMEgXEMNoSYDVQ5GPgMPqKKHyLY
eMdI7pk1Ta1+ZIcHX3gKwW46gt/Y4BkO1bShCUTqyJTH65ogCakuD+LxfJX8
yq9VJRp07k8EI2zDcFN2zc1O2ipetY9K5RShXGuSDbhP2fOXKxou7NaACLRu
exolzl70u6qs3EZz1e4QBfdssYua6pKJBHcYfBaH3meFqlEINkiPhPeLQOyQ
lL0R4XqmZCq3C2X68R1YZRG+z/c2WqLAE9wqwEFSoa8MVEgQebeGWMAzrjJO
TZZz3a52woHZ+twvWJY5YDTd3RMNNOVM7fLF54sY7rEQ4MNOD3k7LziATTtN
DWHhrohJBbwD6q/+bZaHTiQJSyvEq7WcUYyEymVqxRMZ/7le8UO+KZpC/vfm
l0ZFrg+0rNU8u1fcFvlszMGtGXrYTOqp4DcmIvn9Z/tEhWkWlvnnl7XGXJJX
vU7dlzaCo+3SvcEjSZZMbGxplWbkQFvQzkAgqCRSvq9NN2knxILOt26diXr4
u4kYxC656upzkxEZdqEo+OHjUndHVOaxHrMC1A0FuREdmGqI/2AcdVXmER7F
EuoZpdpzJM3UmdRW3vRxCnEXtTGHFpiMdr8weCyjVtIprocAqvHE56fdWX/A
9G+7O3ga5a7xHIK4eNb5/ffBmwk1efz1Ik9LxJm5cnWOkCK1wizMjq1ZzGH8
hXi4aEQ+93qjMWpS3VYAI7UefgPJrCM22pDy6p4dx5amFaBQiD40xGTNT/CQ
gCNdT3xGCRUGT+roly2gle20lkTCxgkkHupkpl0CA+V6rUHhxG5lBnK0Kcpt
COH2kbd0fJGw4AhGyAJ+Gn7/zMIwyip0IaqPIRdBQ/1kGhbDMrC5WtZ79M6l
jrssbbC/N1jWkT2+rOPo6ntFX/e8vQ1WsKLeQXAgmo+nzGZXRolIsn4ML3bN
7JT7C2PZ+iO5yEyw+lKG4XEt3LK+P6NaRI8Wwnsq6p0KbzBMWz638kjFwVtl
AD+rMcfkVYp99J8JtbOIDzUVyn80IrSAm1LNgUpMSWtIozDRAzfcFZ2Nuip6
YDgmohWkBrMVVmGcOtHJSN7PCyO4KIsNAwCcSg8Jc5aaKcxmCll7sZxGWOhw
b5xmD6Wl3WxKQOjsNl+h22IHAY7jtV89wm1X3bJigEy+dqNAl8FE6cBpqbti
BsLEFCYNzTGwZulgSW7mUsPEw6qnsamEvYWZm0HWGq8qpRu2jTOcsa3xIgf1
GV7L/KOx29LwtyNbNlpvKLY12mLsaKRnx88c3WBA0ySnMT1+7TjceVWOev6l
FiTwbxpvcTl+phb4gNQCTm3CL9wokR/IjZVv2kfYDYiog0Rc5rupObIccOY4
o70H+Fql9SpWvP8DW+2s+MzeTKSaHaLb01a07UNlwDL7qTVf4+24wCsR8X1X
iFaASPk3jS8XOWlK82f31ZNOyoL4Vwkd/rx3rAarHayCo4FxIGHCV2jSmcbs
ixkhF1U9XIpNsnY1yQcEFLBzvj/RW93+x/JDkEdTu9PIDLSfYvzbP/N9I9zo
rn9kXwA//5NMUqSirmQ8Oc+Cu1v+wyITwfY3zlB9xu/rGYVRpx+i5S2a2o1k
Iy3nhOOfMHmw6uu8ovfZQRobUJC+o6Z5I/ybmOiYxn2rGaeihqr9VQS65IFE
Paoab7ajE0X+6A8e7J5kw3dMEuehB3AtNfnf+m3yiqoJ+Uj5ThsBtKJ9vCYz
59RM6Fpx7KuK/6W3qESemIdbNnFNXcYKOlEYppX4LVBxtqF6BrvAuq0wtLeL
7ogsYP7tEmQQc8DewfnPh7cqnWnBGfdQ134MPb34n2oNdHfWz9lvFPVTFabe
fCDO07O6FZseiAz4PCJXkCQ5rUdfaabp0GVZ1r/OJ+qBxAXL6t8KC/OigDIp
WkOCRCsrvzZp6uxax5YanEVYcHe0AsHjiDA32vTRmPtMFmP8C9/ysYTHhoHn
v+kSWXWrLNhBK4XglJW2GwKOE4s5aBVopR0qowwBG7TXAnxRsQx3XKXrBz0L
EwqrvyQMmZfYQheZp6nsjoRAIicpjuDvisfRyj3KPQD7C8M70FXNUJAgl55b
FO/5K8mkNi1uaGIn1r1FHVbvSCjoqkxwmILgZp3KDS4h4tjev05bUnJ5ZXIx
Fe5bj5/aV0xhkq+GKcHALT/NAIjSmejOEqji1F3CTM2KuI0uDU/eofG4FTfw
CAhRUgS/lPk99ltLStEQNYKtCM96u1AZg508d96bHWTPDd7v2wr9fu5mC52C
Eh32NJDjaWDLWJkM6LNk2swiUUefz/E9ySfryv8OYLWU6UabJ5FwaVcTB9d/
7CMI42LUpMt0VQ2XtcOP5k2I2KmevtJ++y93DBTpkWXyJcegCcytfs1eXjL1
l/077VHgpWUNLofVVi2uxCFnr7iJi94DfwxSYe4DNMU/eqzijSSWzFLO29ir
mbwMEN2drVtkxHm34xetqcznKj1fGjxWJhT6DC19xEX6UZcedffOjw1ovMdV
D5QuaYdybeU9uD89YT6Q04HWw1jqaCeoPS/3nw6otpFwWFGv/5Bfwr8NSTeD
d5i+d6sNwoguFNeTZvN+wXdiO7zULya+oWHaXAsWbtYfMqyPC0Yut83gUl8O
Ag6eWVdVoUqlSbxpOJEB/iKbaTDkeM24NCnWV01D12St2FKWlLClsx10QLzp
VSD6hQ+vUQoyv/8cEcLyEw1uNNWerOBt+bTC+HA9aHlSpD16qaQGkvVWDMtb
r0u62DrGRIucK1q5GbXIE8zAGlqhPCFS5jeU50AtLS8LWRjQ1GyCFEHT667U
nRVfQn+7Ovef+dBrnLpLHviQtS+sDGl+zwfrwl40yCoY0xX5vmaxnD1ExRBq
jPbp79X1pqP1bKsxn9FMy8s8WcdkfTtEZBDtSrj6aApqfoao4md+YBx8flO0
2R58hwytZ87DpecMK8UUwa2WinbWYNMMnrkdEmPXc0y0zGN/fau2PJinqQy9
p5guzpV3s7JsyJ+20w/WKQoltEyUptn4MRFibH2JqPxVG5mi0XvTIV0e88iz
DVWeKTkVx1h++3cOjUeWjtumJ2dR/5hNTS5xmBnWtJUEAFbUTN67M/mSW6jv
azHxe0v0gluAe4Ta1mz72MDnN9UtbBXDdXdceM3OokoxrDMHEwr5JvyNEq+p
jc1WPE0lNzt64cP/ETmsRjFqjYw5f9BBemWYg7HKIJGA4SIli0ydbA4JxFo3
WZ7scghoRcbrLrARddfH8uA9jlHCgTBPDMzh6SGLkKEHN7gJvpya6Jic7wmW
cuLniCQrWNZrv7zn08VyOuPS4dV6p/6SUMv2MLlZaIY2SOnKV/Cq1LiclBuV
VP7o6sAdVMgEMhxuuadKze2jmvgTo+JT0/tB/pRUn6R7aW4nZLJzAxdmrCNc
bclc56vOoh+9U3sJN0+5LH5P6Xv0/EKf6xulfMEfbBLY4IvjDmmNyBGeqBK3
lC+AXw6PLnU001P7oY+ZPqYK925b7yTQZpHu14KRUrJvA6w9Lm8XzHSwQyei
szP2pmjVLlBo5pKVhKhSmwUI68KzwXVVKOJvlZzF/FV1voIgSH08ca76lMP+
6bDs8dENNcuk5qFGPIXIGqteF30kz/RZlzDq7FVoatOHW2Ww2UZY6BGLwuQT
Sgskxa0DiZPGkb2LoQUvn3FFAAmkkLiH27pXlQAw7nv3/CDpvrehhbiwoFO0
hvHeN/A8uqip/OxFEnpKvMg36BDB5BGRKoWEeRlgb5LlsZGPVehKN2Ro9KoK
PqnnEa4EE3uuSRsA216Fed5oJZe+FsvJP+x3iZT5gIoHgSs9npjUEXGdyn8C
5qUPUn4oeCF183CnXo8w6YSI+CJd78eWnw0njekabNJkOeaxvHk0jgymaB9F
ABkbB/FOiz91t1lUU/ZdyXXlFLWwfJvXLdkYh4v7DQ6Bzhs7vH6fwHrOn9lE
Czw3iNSjDsVBMnl5UAY38qk68zY64MnH724nf5M+2AdL0hF6cShO0NqCBQjK
ALFIm+AZaNJ/hyCFzyz3n+IYb21nRvJNBDFmpK7L9Ds+uDy9cxjSRdLNN6lW
YYXhJDb9osnvqfJb9awHAIJ8HmmgIdkfOVQGVgDogP0kjE4kZtusHDSeq3XM
kisDYf72ivxRBCxhtdDDX5mPKm8hXvTebwCgoVnHBR8Ow4I/ibhXn9fqk4Vb
MzS3qel6u3UanIk9kQpO573Rs8JfrU1KwP2+ZTngTFsqik1PYuOrlDEIg9Nd
DxivYEYiu+ZdwmYhxu9AOhiqbNaOcUh3qnfw4l+4/66X3lZVWSHJXCh7H334
GsOYggTlbZPnZg0ukq0N1cY/6MU62DhLPgZVPPFaewN4D4X4EoaH5r74/E0F
3HIclS04FL8iEi7XNXHbE9Uyv6T0JAugjk2299C2kdLJUDluIph7FoluJb1S
BN4gUqTJLDGZDIlMZ7OzyiGea45Sdy7GkCwKj2O+nvrjy1bHqKbb8f7lNcr3
uhfnHlxuzmaOW9ahr6y/zbHwvt8ZKktYrck+kTPabZey8kPNe6npKeShTBU3
fncMZ/2pdvRBsNM0izkcrkgj286gym9ys5fnk+XL5BiCUq3OlORKSMaO0Kt1
7y1jYPFt/OcvbO5MrSBX+I7+Rm8PFwUfCOiKZEJdrbs6T74Vj0+E/W4fnBfG
7k/qqWziAYa//nAehpuumkYkPHwx72kVeb2VeWf6viJrJHx6ANgMQUA3RM1X
nNAH0NNO6Fuwy+zC7aSZib+c+LzCAkGgZ3trCkRxukgb34y1m8Hdw6Xu5RnA
A2AyHRg0swFJ/f/u4lSEHux/kGkQyW/9/tDVyDpK9QJQE7XthJMTtPgpt2LJ
Y/VUCyaZA9TuTnwv5NOtXLG7GTj7KCLNXWo7au16bDXVpKNEF96/WQhkzK1r
E+AxtTvJ2dtoGqpCO/ueZw2Z8g9oL/jotR2kamRupetLjRktbJNowNO0iUQO
yq5gKfiqm/h570UBDM88ZBuKU4YW8NxCLormBgJ4gIYptTwX6slT4zyIVL0l
nEG/R51sunncL+mKimGimXhOWqQinJjqCQM+FXpUEsq+hkU6iWDUCxZt6HMm
Z2wSa0qxL8MhwEBf+t4uAgCHD6U14ko/xGBRPByVTvxaM3Bxfo+POHtTRGer
v2Q/8i/PYeI44gQ9ARqi7u4uyrIpF6/ds+xsbn7q1AV7Kz4EqjHMw3A3On/K
ZuUpNH9QYzRk2vE5VpRuG6PUhRb0iImo0FkhS6Kp9SRM4LZoOsHmATKnOJo8
SkjuxO6BK2IfQsDvYjVUnwQKJEqrp9WhAQwFRZZvqZto7xDe5fv7a2DLqNFh
wSiwgwggBeDIJuLHZff+gbAkTaDOCGfYwB5fIuUeXWyd0vRw70H6tYv4TEEn
IGJcEcx+yqYVponJCVekyD6RbxwRNjE162GrrA7ZY4gHTIP+0lzgXylgmyRy
dEZSoB2VVEjkmtVXednSgCvZYAcL7G6rRa+0vpMhzrhSv9Jgp7ytWdhWARyR
+xBgcJBHivNtCZUP7ebRYj+5rY+GfxlQrlDSfk2skYGkksioCpr2d1yhweUF
bC6j7+K+p/m6s4l1bJUP+iSZ+QT5ylXWGtktkhZowx/tv09h9It4Orf4k78q
N34hN6FKJbRda9vKJwg1qHOQItD5xPdkrNNo9jw3GtdiA8H88xoXz4y2O13U
kj/a0uAGesVl2v+/tnl4DIaBuQzK+aPrZeqtrIVltnQd/gJV8FUz1Nslhamx
P5FVzXuiA+KqXpFNbw8D/hZXbm3kMQioirp97gu3qSGfLtPIjOG3ys9yMDdr
SBswud2PeflMJuDgwxMFo/3K9bnCbQ85eaQxQL/nt0W/6b6U6BgFQUVL0R0n
8gHqmBbGnoLnNp/0AqBlECer+wFrhqowpFsMIF/hPBFQLDXG+CwYfYsIQ+Gk
tmzXwXgkDyrKSC6QbSfZ8U/el69VEF+kDaayklyAmrNK04YdP89ajEoH8LZP
PxpGUNK1yEHDKAamWApyiePYZFhWcpwi4fDF8ph++Secp1jsUuO2a9CARufv
jjQjTBaiZXCFJM0jrCijb6TX8ulSOhQ6DL7P1Pr+rXH7XgiKZWD0MS1P6fFx
TBSSxlplzq4lnX+PeNf+iKv62mA5ed+fI5RHk4VYRIQgRyZE09yPueVe29zi
aks2q5VwuAXOCT2m5pYD2LoqPwOXs20vcad8QocWmbXAABYYFQIfI8o+yIyr
XVbmyk8r656yTtpm2gIQf7AuiT2OPxkfcSfEpdxbPHt5lIGzrsrBW016rjj+
bJ1Ki0zDC7IVXjVCbJsdRXMfHdbIbrLACcxV4uCsFK3KCUqMqdBI4rhUp31u
igLxGr/4dVot1JG+AGJY7Zm+QVkMU1KkzbMJMIK7AuhiNRSwzVII4Maut1Pm
Z+zVgdSasbMtCrK6P6G8Ob5Y3ThhX1R1X+eETAo2f0eBOMKcjONPq86ACDxl
iykeOTqMHyD9XaXx+Z69kXoVQucBzCU1OU2Orki2rIsI+RJhPPJUCstM6Sas
F5LcZgnZnA/k9xBEx7bYBoQ0k8qm3oHBAFn8W5oJQ8hn1Wpg8rKcd97RDWUY
EsfwGIR54n+U2d7+az7URxnNSiTlqNYBTRIQhF21SBpZqcxr6+eZx9NGa7Lw
PXyXNiGrLwbEB2fCQXU0blNXXKQOm9sIUwWXN7r8CTgObisx3nPpNTN6g34C
HOZxH7nETBlOJTvqurCHxZOEehYgM9c9XDm9ycp6gGVpDDD0dSYtXr/X1sgw
/tjJuBxUxl2ql/HM91D1CYkI4fjEGMKlIgzOWy34Dzr2ETRupkRO2aQsI2bf
OKo9nPshsTqNjPcm+FC7obI+AY6z0tpjqoauj5llxWE4YeHkDkFjBrVbceDk
6Bc8EhPjBF3UjEnvYTNszGuOeMulbB+vUuH4EnXZpPtFbanMMOu1sbFLJ4TQ
h9nU40Wi9hP/yfq5dT38c+/nAqlGvrZ6Mx+Rl8OGpMNnNuuYEO/Od6mwxIKT
J0/E2egHnbH5g1G/gY5LluyEMTiFNMOB0vRGvQnI+zNbkw4RXZKdJfYkpmh6
VGeHrTKcjGs917TbKon4jDwmv1kjIvXyOj0e5Wd3ZbUz6MaQ5N0iOl8TlIbH
VvddrsKfEHg3tx+glFlslAwBy+FY50JDc+sIw3Tq2BhFEB+1keVLZuQqEaHC
e4NreWdq+n8qnompMcOgovY8y0+856XBPVFaS6h1kLbKeg9HoFzordRpbglX
UjZnkphH2Cj74o7UqcWXue04XqmWKoP3X7TYmEQ4jUncpRuSARJJF6Yt03ey
eeP4t5FDaAhYaqyHwONbbwvw77ZcE0Mr5WWLU2TBJ8X5PNQaWto9wmBxkipY
Ye7UmgJ+yIZPaWU1E7WYopqZaYHr9GVQfPxg+Y2FsVzjg7oiCI0QBI6ZqXmI
T14Z6i+Ql573DyvgQRPG+vFRFb8OkQHwu84RK2loNT9hP2t1so3M+S1CHeCJ
O1F3fO7kDA80tBzFf9NaqPQm7nBuHDto8HC6hU20BcyBIgzLfiSrq7DYciL+
XSHPnySFqncgcbkcAN3nA6Mhu6HCC7P7DJB+JHkjeyJhc24dPQj1/uEq7Q+D
3lPej04z1M1mTPFL2mP97//zFYGAvSM33vPACc6El/werqTmeumC4cJpG4Q8
a4f3gfTwWQzeua8hsrfXuvHaKVbE8vcQAjjVNGei0sr5Tah/LNvqmKEwNobA
XBRoP5oBnhKxbXyDSZ6m+HVO0KBnJvfPCv1xzHb9R47+GQm1l5bk5Oa0+DF4
6Pj7cuN9pYIcag59FZJ1c+Eo03zU4dyjYuY50PGuEd4dN68vQXzPIUosqEyT
1CfvfcOrOzKA9MQPn+7MiwcwQ8HgFeH7j7EAoNe62ZgCVeP1Qg+rjk1/p28j
YXUyqUbz/RdnmTEh14xZfOkTNP28DDJ/kA0y01KcZM7MZ212UEacox+HzlLO
Xl8ZAIavuaS0esFqKzgMUMx2ZIheFjcm3uN+ldN+2bE/WHo/wZeQJ+fGBa/R
jCF8tStZwbXi9A6lrwVC8gKgk6BSgBZSeI8U9qaCPeai54HKqRdYSSXs2D/l
ujelvdueoHMh8tbG9mDHqWl0hMT/aSwvkeRu/GxV4jhQGu2UVCzdRsp0Twu+
OZjh+3xCED+PLtPozIBvoGdbljXjd9AIHapGkWV9/TXxRBd6Xp5ZiYhJyfT1
o7eV0Du2aZQVt+vxv+0Y7+VbCxpKqdaE8akG0B5BLpLR9G6kPi7KMGXd0gPv
2HTZJ4GznWw+IjvFnDhkugjhvMeFTxfVTMu4oxYZeHGfcpL0ehwDgCqLLdEs
YQeF9Bq6vcPBQ/lLz5OgnOinbuIIoq4UoI+m3IcMYYJ1Ija6VazPaVBuGW15
TWzM3o3ON934lm6nr/v7tj2NC+721nbdp72a8i16WyYGG0U8gI8VLotk1IyC
uYN2XeSdcRxN78wUgC4jYdtZGzKWukmyuLUiIA9KSQs8OZj3aAC/V0LS+7zl
uR97aL6F/pzRNEexma3ngBbECEECPAPxBjRQVH5XhsYkFZiHaaBNB1pzms5d
XCKkvkf5i4X8mq2R+o8PSZtivyERTiQJpBoyZEIB8R6QEE09Y+Ao3GPdQyt0
/W2CaYxeylrT8SV18Ub7PZBUKdEWNNPol1RJJiXV/NZcCZ5Kfn/qddu4OZK6
GXF925YJegpmBvURcvCJR6nATYEHPNlr6knH3drsZaCzDfXlSUUAHQ1A2kgh
B+Yweyowp/BM8lGiNlNUAXk75Eqqrz4B5waZM+0JsREFmTTzxImIlirB+zXc
NPBFXCpwq+Ip6ryBa1kwbUSACMlr0QEo9/ZuO6YeTdw4EllcaGf98kt5iYmI
tcdjigYZz3+Osd5t5Mk9KHlGEjtQRulZATukf5LNF9Fp/4cLcdiYsGwpvNJN
nQOqOwpte7/tyV3GrhBPg1n4mmMf8AB/nmGnpDAMDzUd+DE1ztkItZW7Gbr5
UJMW8wRLB/L2p16m9G7/7NwR1wvZtbI+eYvA2rwvpd+SNYOAWcw31rAd20Rd
0+PKHtCrulL4TsapHO7QilVxpz4elbKTZuISHnKmgVntMcJyt23zwtO46dBV
WEGuquJ+LP3krk9myp7rugaf3+m6HoK9DxpVV8ogz0Isd6scmcZf4ZSL2SsR
lY/Eh1+pkkWsSDAxDl7NMTH0zIqT3uOwhJd4jGFxzMMMfIrCEV6k/EXOfW4d
S2mFMtNk3swSkd2yrQYXpOdKDqBa1WF733iumdFMLH32W++iElCKqdNijH7K
G0OSpmUw5ng1fibQ1nA1+cPwF2YI0Owg5wja9LWAAlR2oJswGyNByQ6GPpiz
KMH9tcMt2BUOmqiFaTrnydLUwbURhgzhcT225pO4HcYt/a4UupQWxCZRPVrE
l9OdizCTQE+SNUIn4hqFiufKp7pV7usRyhWNc0h4tvJ9Bx7fzRO2pt0sYq5R
XG5xPm35fy2kJipF6ycQqvMmo3b2LfZ2lpGaOfOawvZ87RUSOANRqYFPDcR6
yCxsntXXFX7e9XJpbf40kOnY9/U3NQ8i+MNO5yeh2t2qVtJQ4RBEDvNoUJkR
TCm9PWI3Oyqvv/nM5Hf2oubQqaURVHoWv8Sz1mTaj+ijuu+MCSZydkUkrCji
SRHfDXRpTtNsH2pb1nR0rJhFIAs2wNOmIxAAMcl4x14uNhPW8V4nDvqc/UDI
ccvnZdBMeHxdPuia3jHqyaW5d8lWwhr76NMivTvuzynXPKq2JeEvCWJipwDY
+AX3jQi6bgW3QO7mfpaIRKjd/2NWnldGvp2tU20lDNZ5dAGb0mTqkYnc03FA
akhoPR5cjE2aDIG0sCju/ZtPi0DkQ3Hajd19hMz1xMJbmtnLaUgmQbr5O3Oy
gEbmaFoUpZ/NMIDt+rRq4aTk7qWQZCRJXf5BbOP+cojU+padbTKx0fW2ly4v
JNEpMH0qz4WmxtYVjmK/bZjNTCzRLoLPgY3mpCJ4B++KcyHEqTJ/SEj1da4b
2qIJniYI9voXVEkEpADQZZWwXwF1AXJg9Z7Rx3uGbQ1HPfFULoT6slQ9T8yk
LfytWk8TrpizT3deyDt9oeR4eQQEvKHDZxeAGZvvTrVK/lfrnbhec8HWpgWG
A3veiVu46VgZW9IayxYfcbC1fO+3fe5UshnVvuTVk9AY8zYLivg+xKNH2YxZ
UI8VcH4iQxtqYNfKTpxyzHkV9RQOJ9MPkdUo65v6TwlhwYfGWyk4VBED+qR9
rrOgVo8E4ZILyq64xyxCFcypE86qJ1EIud70YDWdkIEwRXq6tlKECGsFP3Sr
eGGjIZsI98kMZ55AWY3p8R7/Em3q/AEQTA+54XBzEnyXihuMZCb1qbCMv8pP
uxcM+vw1oQYziXI14faXRgxXi95wJZHs9Esv/FUWgAisKQiiepFlXe3y2czD
QsxQvuwnD5AbPuM9a5WMl6DjTY+5V9jWf7Fl39rc9ktSbuVtAOtxquJuRKht
gbMFi/eZixIZoJIHa6XXPn4fba9c7gKzTPPqYuKbY7RCtXmwNGkl5fA8pIVW
v289Fpy70NKf8odGd9kXEvJVbqVvS+yET0Fg8ENYhcFtU6hb7BT5ti4EAryn
KNZNyuEejTYz1jhYUlVpjrnh+t/QtCrSTifL/bWnpRWyKscq7sj5Dt2uDyvR
e6lBOejTGrbQ7BFf8ntFlyqj14RF1KJtJ2vLSB1Qu1Z/UKdyjvWQPiaHbGuJ
PAdMlkjCPNlkmXeNOspwYqFTpjB+hM4PCypKf7dnOMetYU+mXs0UJZIl70r8
bqp1k+dPU+XAzJ+FsQTze2dF7pAmIEaHjaimkj1AX3jzzSICJxpsiN8xuKKt
AZ7gbVnsTaOElcEDfrmWhKSNoanK9lQNZG+bAi08Dx7r9icDATfgtUFW+2hm
ETx9MArm2HOHLvK/3ZnrLbSmAC9njZfMnoOU7mafJteVDEK1dPbHIEOFuM3B
8We3jJGJrhQHMjsgf6YAvp566h+V/xE/69xf3PhAGvCJ/ccCS29ZqGLY79XM
uEfC7KYbUh8H5yLxQlNKpV3ITuhssl3ZGQaf5cLFQtgCo3VBzXJVR+Tf2jkx
03ginISohHVeoscY7675TvjJW7WfUZv9XtMVdEP5KSk2p3ek8CIuUZh8iUfy
OgW6oM4z49zgShFQRWz8xDHAYK8hoYRdYJJX1lY2VNELum2AFPpN6GpD+Wd2
C0OgDmEPASXHRyQE88eAvEyxY8FCBECjsTxANrm9/cG/6inks1pGh32Ojvz2
wyzPc0e4EWwtVzFfsCbxtHlGz2MoVoXFMm3YMoK1PjB2lPCj5FPLSTIfHnjd
UcGp19oDFq9rYv4v5d2RIEqIGINYip2cNomXHn3/WF3D8IY0nXAAe0egACFU
OL67rAb1YGujkjTb6md0K5Ekd8bxkVaVM7TfpIz1+xYxa5OhkZAF/a+XfXH5
6SrbROdIxX4iXj7LOYW3cloK3XhKcp6Wi3d7wUdLPSI8shmKpnIdWO/eoO+m
46jG6yZCdahcvwCaEYs7xCCFIbQHl444bDqmfdW0caXHEl6aFZP1gHTrdLJ+
hHULrUgh3p/ZwVrTVim/32XVADvvrRMSOW8FSgjXZk1YTUStrLPnL+G4SqKb
eDW5znoy12CP5ydRyxJP/qdWrRAiYwhwFirXkwToDJnk++fO/Evw4aJd7chi
iGNPw4NG+LfjtLfhY/9Fz99Snrt7RNTW33eDubpl6SONP/ugRibvwAaVI6yq
G9XNLKZB8HuKmgbHrYjNs07sXwRqp7ZAWCHgSSOcafH8vKf8eR5spBZMTGOC
XkCOoK0V5ssYsxUlcsUj0harRLu24SiSFRpAFSGmvbsCNREXmyZvMYHS7EFT
3oo71ZlU6OiDGJERdy1xYEyKBy6EpicHEhhFwbi5pefYz63AyXYQUNj5pfOE
0RoSL3bOo7x5FTYcM2M+TZFHDC66Nm1DtHxv3KUg2g7DfFZ+j1xMPUF3j9uY
ofpAGJeUku/crgB/Xb6NGBl8JjOi3knaPcdpi6WydXKz4PF4Qen+JGwkJwn+
fzq04cbJ+eHwpx4Bk4fcfx0w4WW1DVWglZdvFyievvdN68G3Sa25b3s3FU9T
S4EMYj8IDULw7J3U3nbEMI8kKIMSG7c49u6QhKmBuwG8im3KoGPA5YjUm/M6
jOYk77CfDU1OFZtl1h954cWfJf5dsQx7oi8/m3hZZTFmpgUlACHtscX7lBan
l/zfcBlbk+QI1yoL/lb0pMV0YDhiWUUKLqAkLkwAfznGHxc/D1d1EMgaacXz
yniG3mi8qBzL/l2yIArWrvWYPAsNzrOaYQJ8m584erDPa1G34WBKJsOTXfm5
dV/pkWgkyEqbVvCaeVDLKg+KkoJvm72Ym6qgFeWDpOFGH7mio+HKz5Q662XJ
XJNwk+5vJR41XFHrd4cuZeb2jjzJDz/bErPaMDA5XgQXzHr7uMV3meCBpEdB
7Qxq2T+McpYOVoafQnq5Ju6aLSrRPc4+YYl5Rn9cAYFuCbn8Rzyvz4y+LdAZ
WelvN/tmnbz+HXBCI7sr6Xx8OKziEqDe93tnq/1vAgUiIrzMAJq0Rzf82Z7z
jpH+L6JlXt8h5hjlD3aoKAfMzKtJfJoWwbQcZ309Xq2Ole9IFg4ygoz6knjA
q5m3ZisG6aGOqgQiHCsXSjQb7cK4xdhZTgPw7vW0WQqgxhWti2sEtA1TlzVp
LFKZekukok/tzcWlj41WveuklZPEdv/U6Hngl872TQfyL8OTG8BMAz4poweR
TSx364xeDysRj2C3Xghexcirws6LG05+t3RiGnH6xxB5nDpTFkEpHIUoehsk
9FrQJm5WwpETjgbsfh/ZZzsC2Kor3kR/bEcW+HE8y1X0fY+0F/5gLcE5EABH
BhRyHcCsd1CD7J59dApA9oe1A/p4EbCmBbjPhTDwwWOAIQuJu/05Rq6/pcgJ
au8s3POllrjGEAPHh/XTqV3w//9kf3uAE4r4dPUQIfeNM49mICiL1+YCuOuv
defwBj17hJkDnA1g0n9ePoGD+gIYYV2TzxzmPDw4Thh29T4OsgsLGh0NhKpD
M9HRWYpx4GZY3dVVHmATyA4g5W+o07W12lTD9yhnYMaNThieb69DKRpsUCdH
1zFsNJAAFuqixminudOrX/ZmlXaHq3F7Uxs+wwSknKy35maVnm5pugODVxm6
j2wwNODnNvmURvB0OWq7sbSsEEK4/5x3TF/R4dKT+rpZVlEEZIIyw5cq6DnD
IzF/zuDlmq54yY0TzjLDhXdMnMdeaLDVkbeDAUDdR9DRdeIAFnlHbImy/U5L
NnbnCwWXF7tvvm4cS3KzBa/7NeODF39I37ymdjhNQQI2YDr92YH1fxLXAIC0
4lVQBq9RTHnn/sKCT2lP/ukR/A0JP8zRyzu95EWDh4d6K5PLri/qz5YiflOG
wHPQmQykO4ZO5zvnvv3MKpxv3dYywU5l+lqfmWL4jLbzcpMtCRIbWvGB0JPC
WC3dnLL93t0ycEKjUzIr5jOfV0UVk2W3+D51EGM7CBrwbj1tcszXVwqK0zKa
GKqdl/QIhC+TaOeBTZXMtvSdmO5SekpXiMZC5jci2e4Cik59dbsay6aUYb7m
KDrCB8FNIWp8Qfd2Cxf2CTZJNib7frSKClRsGCeg6Gca4a/9YxjrsXQNsQtv
1JklPe2gOZiOWoPlaTB6U9kQnluGGTjplq/r8jqVdGLsi6gNYtyKTAf4MAGO
HK9I/K9jYbu+CAveyOP5qhnhjtHNj0xj7gkvF8fCXHFF020Eptd4v0YBW/L2
norZCCdpojHBg+Sv6aEdbbOw9FT6aFhocdcpwALPLbJAWNMvsOmv8wTW25eA
ljR2JFxURd5A5WbK1LCQpEeWJtLgIx/tTptx8xnHcZxXRUHRvHN9FWK5SKEE
TyhQM68tEJWiwt9Oi6hFPhhQOU7Mg7862OpEuIFTGJ+Ksbg01rtSz2lqhVmf
tDcAYqSDjFnKQYXSqS7jgHar6FOipHZDzUnxcyOmLKEhbGxLWmQBKOEErQEI
tdKLmdne3iqmBJmU3jREiGkMkS0vYhljNOVvCSgRJcJAB82pypUEzfMDfQTk
o0EgRl+k6zcvEtKMUKm102Uckutndfid4GKbjJ0bINIVKMLtHjAEYoECz+Ay
9aRAZ/UO5eT5LIbroLAQQSk9R3D+mp7AW6E7Jn1+IrZ6d/ukrx0OwO78ZGTz
RYPei9hdDnHSK3x6JposTZxpMljsvYJ1pJ+cZgqASsoVePDZShDdxhP8TGke
Kqvrm3RFBBWdiSaeF7GOldqD+rlx1BtDGsMaDUJ1HY0Js7cIm0x/XzyT3EgP
dwE4aWEmOJBuwl/zZ4s9vm3BBOj8l9zSNkgf+gxbXPM1wP5+3eBP68eDAnTv
OUx0DiR9uhjPvLPd95k+kRyJgTQIt06d1b3y2EKGzLBluGAyG2TGN426rsBi
UDqP5WyGViPcia0zuyeOA14Wor608qd6P1ymgwkSndtouX5L3Sl2ajVTop+q
sx3Jdp4iG/3yxJvfwnA7Guz3tQ3JocRHcBHxMPoPFkX9mP34c4RBRgzrQB9E
PQiQMyxqXVUH0JiIKcdni1YFoNuKD3d+Q217Tp7XlDubIdqJs0GZUGY+3V7H
rJddgflWvhXpSE2og+wcy8w7aP/BMosnOmuZOc7lTv+7ymmpYH5R0UnMzHgf
82Uzou0TijnpJT7aXczViV1Cr/CAPeB4pf81AzpSMdmGFBluf5Cplfw9RuuV
zQvtmUIFb4ma0oJbPc1Qk7YIEoDEX4v5BKEAmVhVM+A7avwHcCoaDdCUiHIX
BmqLYcyyu5Dqsc0SpjoclyiP9l0P2+Il6IUzJGg6eGCoR392Rs2KX7a+Gh/T
RdP9XOr1SqEJnxQEbkqaddAzIEVmq+ypGlj3HnaFHGoK2YMyoyMEAtVHcTSE
RSpd3tJ9IlKqo85+Ymc05k+peG4To1OT4oKhtaC2npAvWMoNYuQRZvKiy5m7
eXNdc7Q/S5G2YYOXY/1FoLyuTCtmelX2LHXxHeqknWm8QXC+u3a0emwIP+x6
7xE8b9Z/i3bohApgtlINZVAZ8npjT0ucw9kAiNtGjPkOX7yBByWa+LWEhmXP
ovF9EqNPaN7RVCPydqVuWufGB4oJ1apSmkY2ioEClYKXEfgpX18BFpU6GUSQ
YCkNdAlWO8GJPVf0//2QrcPrf3BPcdowNbUbgrWAzFriz+1LfVfbgpvHEqPK
GxldyADwQ/3cyXncxz04PB2JRbpPelKdLYpU7HvUBoY/X6X2MXC1X2Y7JE5G
gLmhBYc25plv3yE8vAdr/vUuBmHkmeCDpVJv506fiAehPMcFOFbDlhg7PL4N
yWWdYjhtaevkG1UIz91ZBZ9XBoBSsQKW/EHfOu4nyuMFoTFC8cOZ/A9Pjdqu
zl574SLK+AK8zM+xJPb2gABffBIuEFtSzybZ2iHNglZ+HWvX2l0MHnacTH8F
bq8zVC1dPaGJ7AA9g1gHLfQhkEudCXizCvC2VY+z1PqAyFUa9v0fWC1gkFju
hpedmBoVR39oB7/KH07S/TjeU6ik6Z2m6Qk5LAbm08psHYCHGng0OnG5NPjR
M5JeTHUdblCYHYvBK/AOPzcLCOYATab9IhHDxTA+biXXFadwD0JX6OHc2Msj
tT+c0rEFMn7RoyXrmm6MF3rMSMXe72DeqSi7Nt697BW6z/YHt+3PbYTSaczG
CbJwyGb4TTRBTE3aI/yn7PuRAf8ZYvZWfvnmXeUIonlmVkxb97rnAeMQLyCw
pSNUeSsDY1WBaV6hYvnkLWp5ibOG30KJXs7DR4G053jnBkLDv3GvNVENFWmr
UWXl2z4yowspySdw8FIrLlFP/S1jSCR4BbEBi5Mtd48B0X6wB/p3qnuj2Trx
xoxXjcVlthmcbKob5X3fyzlCA26RWR51c3B+LxyOms23/PMT1mCsmf0WaSWX
6qFV/I4PPxmMo3oCQOSnaYuPdU+P9X+DxR+PD77r+q0YgiGsqyzb1SRrJ2Au
hjK6hQFeMd26iLnxRQwp5dyy8ItgRuNpaJHTQhGOFcQ053JKzYCgWt4uVpEF
1F56sBPKIstyCD0Ax7ibsI4W37DUx3ZnLYd9TXbbiCk9JkuOw3AFF7/ps+8E
gDQhFgMhYQf2WsZisdmwdN34o7eXgKUHs3Xg89fuq9MTZ760ungi8Ytp0frE
3eCwkBCjN98VT4CGUhhfeVBDKUAze0gF4ey58GbJuD6DawRT0csV6rqqES8S
0rSkV7LajAM2HBSJnrIsecPZueVHPyqc+p1YSC6LlHfUrpl4i3x9DtfuBNL3
ARtd0ka7VApKZnPRvKun7b5LRKz0xLXlufK3Qqv4AT39Rlvf6V+rpNp8zBfO
YuFpB0Z6v/5c9TccsMdR8k2ZGG2dZPNkj9KTMOEFgsSI4f5PxH7xjO1AXP51
9LGYEKvqSOFcIQJmxHHkEkqFecjJtzJi2CGDmP5WwOM4P9cXy4wxKEZ3QPIK
KRMicYRuGJj+lRYSDMxpEy+fJ4GNhudDR9Raqo5dVzZwfmov9Wg9g+zJTMzU
gD29Zy6buX9YbSJ6fFse28IdyUQKI5lcH+4ih7PCMEOOD/li46vsJebHRU1p
w7dNleKDR+8WCB4IMQneYpjRN4uuApqSOF08LQTMqvwrsCl5SWqZDQr9CBeT
FwhBsyb2mjZ/fwqVEVcVNkc7HBe0OcFOgzpMf4OZEbpeS01veEIql8Sl4jjB
L277+6AAKl7foS5XSMVVreWMFD0jBMr6R0mgpfi7G/3z900yBqLb0D6ALuvt
DsbSBixcRUwWbfdq6RqIJn+Hn5PAp9y41mn53rPtkMiuQPBAIrkfTB/OWlag
hkEif3iFR/P/lYSy5Gz8EkfxIiWawfoxL/f2UJot+k9QIhom86i7+k6+Qts6
F2hwe8NyQX+IVIugVxXlbVOSfA4c5kQAsUXQTmoY5Isthi+O9uXA8g15nQlx
OyzCGG1tb2ceu2d4A6o9UkQibzzCoDReXCQ5V7p0G+fOKq69F+Xd0ep01WvZ
4fmcy59pkkwODc/2roeuZM9clU0MroQB7HldGmeSOegZNwQXbghwAJcqRKy5
+MhW86A6l/Vjv5I1/hJ2O5QTQW+Udsl0hOeVrm7/WU1EY1GP3xbTyXlNpmQw
Hh1SmSuDwp+SCoRNASZWiO1ODleboVrqL5eS6lqfu8KzwZrBLotnBFSzSpvT
gBM7ViZ/j06D4dVxLaaWb6GBU/x5WUbiUa8f/hcmhPLk31GgbTqlUR4bkoRk
evyPBorr1VcZlPXN/pZ5dSQBnNkrpyR101D6jRmh4UFKgYx2n+QOqcT/JA4j
d6i2FdPu0JvjRaXcy9fwAmBIAMoKs10jOfrQK9d6ouTcl2IEmNGBB8GP+f1n
Egc4Lzua6kOtEH1FnJ7niEm+3JV2RqPB/M9uBafUDcvkGfpSyYTqDF+xAT0/
gZkaotGyAKrdTGDWjSHxqVJPotz9e++BMdaB2eiYj8JFZXVJuv9FyAXrkayO
vwc+SChId2bT+wViVXxw7voBkwT+5JAp53VK2mbAVxV2WhN+p8580zmlWc5h
DFgymvzljdV12gGR9RZkd4TtxIrByYT8l2VyAN7uFdQSSSZUitTj1Q3nz9hH
WUWsMUZLLrRHvnTewxpJdH0/eovcGvVXGk6+AOS/hg7fBzn5hX6VDETXM5z2
OoikqcRyu6pqhp8oMB3mAllXVpOdLItCbLu5FNK36YHwXOTJ266ini72G0t1
8C9kZbGf3GAjjuLA1PdxG6mGNMDanHiFn6mBJhmf/RqU8jHHZTzt3DhwoGA/
Dbf/gakk8NKqFf9g8kVS6kiP6KTROQoj2eJ3oLVlS/pLjWlmF9gsIe1AxtTX
/s0hszuGVvA+nKnkx42Jw2sj2MUoTbe5QNgGmRuStvUBqd35Nv2GSKNEH4a0
XwPsVNSARZOXBDhTUl35R0iOwi4uVPGo1FhOL+zScD6eV/gHPy2UHXnvXAMm
R01uJvtbHD2AlHdoTBWqnIWhx2EoKtm4gfG0PFXqp4KiDKutB4FUSLU3SpiR
/N2vjVs9ML3h+9Ih0ogOzWBxjfIcCogZ+HStAP03dPSL3dcRqknrxMwY960o
llfG52Wlbdv8yvB39GXz6FwNYxiNJWE78BovhdWlAPxBs7rzo5Q3OwGg58Ok
J/eVEvu9D2dDcoUoh1+2rOVHsYvL2mRlWcx//1veVbdmkueErwsQbaioHj6r
SRwnaeQu25QmSw4KIcrgWVrUC4sccewi0OG1R4qOJitmnbK1vvBdATkQlpkO
OECCOLc5o6ZzcEKPL1HcW9qPZ8BRvUz3+zSzyXc6+Wzsrbbc2jjOGvJMRmQw
b+XK361JVPIqWDoQU8LPiBYT3cDOh3+DMAt+L63DlTgcIRIytqTETL4Ggapi
TnI9wqTbW91e+wgCv06Lio4GRFHPGtaSysIikPAwDbBJ5/nD/Il4QX8mbqNd
B38Dh3I29NhU6tg3bZ0zlkh2PAQ3JVzpIbbEOgQQKFX1DdaamvnTDPcgZ+El
PGFngKN2e8bAuUBZUqP7D1pDMC+drg/WN58k9yZ48or5uIcvuRf2JnMq7kgn
ytp22fuBVCoqyT7iT8zdJIOEwQTrABVJUW1XxhBSgj5dQDfIK4+/lWmoxBfE
g3r0/CkZiOcY2fSj0iuh+xhHQ6xmTOo5G3luePnKBn7NlhsNVdkfAMYj2ZEI
IbSeLtHas08phS/sPEK82RFjpSD2rPZsV9iyQQxZRisj7v3cPU5+roSsESqs
COy7oIjjcvFS0U4wRcyjdjPT16g6rxV+M1x1e2F1TXXc0S9EdhZPLApWhfnY
+GODY5HYNWJEK0YU90krda2tPxDpQ/r7S2wRlsEvlvy0xQOlWqbvU7xxeNvg
hvZESolkjO93Jiw2fwTAFk5i9v9qupyLsjSSGLm7lD/0FZckngFKCuNqLLJJ
AkqI/QmnrrtI0+TcRIoeaUDDVeaw3z2PZdmR3n/581bMd7nzXLPlPRLSikis
GbmOlo93jvDohU1LW5UFP2BogGEZawmVP9KcwN87hqNJbPHHKulX8Axk7i2W
agbvOUiAOgQlOVEUgOskinhsqLDOSAee32yp/Wg28DVox73v9Y88P5c4eNtE
+u/R/h3TeWARe94QK8/MUbZLvoDKJert2p+VSNglkuVp/sJEaQBZiRGlEsDO
ziA4msv6osZZAScKhFs6eWYPyWOQQ3vI27hxXCeGsG+3OVGdkSMM8hhRRr6p
uCTFHGYgJv5WHlkyjK35jijsUQqbbriI8BNSoV2zhLkbPu3CZeGuT4bB910u
61bkkUlxtNpVWKGCYOP0HNk2MeYqAf5il/LLzV9uZZXk3Pa+wLCtid6jh0zw
3BhYQ0nxBJjQww10SK2WmNaUGluQXopGgbvDCSn9Pr9EwgVMBP09XtY3DxdK
LUqrYlKNQ1KP2EaMyAiPbnSz/M9oVbncq2bMeynNAm1z8JppV7uYOmJEGDFg
aYFwZHlR9C+rKqTgOCdyvUAb+vGcBhA7/DSkpSxd03LNlhWO1NCyK0utLh5e
qlSrFRvz6bPLcgWS0IhnHZP51zGPRqiBQumr4ZU53JAzUCMEcLR6p6lbcA49
f8d2ShsIl8l9Kv/dgJHzBN8+/DlT/ff2IVh1nQmGaYE5uIghsckDJ2GlZj8+
UFrYfZ549a6nVOThtT25nb+t2pAoPJIKMM00se9axqNhUwS6SuHUzpvVQuut
0kI7yUXEY5q1OSuTJ/WOjaxPV7jZ6OltjZf8MSXlRAE8mpX1BAwB6AjXk0ZU
QB5lAxrthqlxv94isROFGngvth5VuloDF8LGFcrkxSJHwm9tfkftSVxJ4Rv6
KqBNZvjYVo8THg6l9pgHNdAW2fZtmAJi+Bi0djDl7uxwZUGfy3yENvL6W/Os
1rtQM71xD9yJTH9IvqYo9JVNU4BTNZ359/LL+cNHnjPwgRc5v2Zg4S3eY/hy
WCAJom8astc5PKrv53bGxkB414JSONj0tkkBBHm+8KPW9vO5GHzDkb3f0k4t
vtyIzw0OQGfDCKfMTXkW+TkPcLmcTiNrhD18pesBqjgEsvpBOc+90ght4R2W
yCGRHbrgy8vfF0GMEUZip2mwlVo9zARvk9Ycj4m0sBOF5fWqMT5hkplHYcwx
qQ0++7qVzuT9oPtM906sguNI9pR45qVfxgZ1Kz+S9UYp+wGFVTlCFEB/ag9W
vGqTktYALtF2aQGW2c5kqxRHRn9Cwzb8MkgrWaWQC60fkqUxh0htElYqbCHd
Nd/O3hWrSbHm1mWEWn812SY1HS11ETcsy+3U25SqBqZKJUhEp6Pw0cgFAN8h
UEeZYip8xXhuuehcHA1sYraIOhCmXL/Catoe7rtU36DnBZ9V9Qx5OVIudHzk
FMNe3Fbf/8iUCJZENvvlPFWXgLT7JkKeumIwlTaHHupdR279mtwmayLelZtQ
+2238UlemTf3GLTnwpodv1yU2pLVrU424bZrIkEUORTJ7od16b8OrpI67ZBX
bi7WT599QMuDd0wmNID4SkvjhFShuarl1qgbRnEtC2AFC6CyOpVq1fndSNBw
QPtiUjKotfqerVliUmEPSVDHBVOlLzQPR4xRCK3z+FotYyAsqNitviCjtkZr
ZvZg6nydbLBwmmsyqOERxeBTmH1xNFASAF++I2jF+BWjdBQwfvWCri0M4LPf
F2jlvBVNG2Wm3eYm3Fcyv0Sr5zg3NOQBIRbl0kRsIWBZcGhRXVtcGSug9EOx
GkvbKMwKQ4sfI5/Wi7r7H4wRvCS4DfKtCIXiseCYJNR1JMoZNmCjku/UxYgX
UsM5aInBNCcX9RxFr40jAiEHDcrzce9Au3lYwNPVZdQui/YQ4l6lE8yLGFIW
Yi4Fj2e/OdPjtxbLvvG45Zy8hDpHyJS/b5oD9BSksI4e3kN9aHpBLWzlWEHS
sZ0MU53pOZSGq7Nr5UAY4dy+e6Tp4vBJv2kG9XXLoCFjKIdS3QBdMSiIXEzG
1qkbqE+C+d4sOiGFSpqzAsqwVpGElpdg40kWYUdOzr9Ll1z9L7wiqliISbIm
9KyFQqfsGiFyFRx7aNJI0G9uuQycZDyufqfoZW0S2416CguK99QzZymjDFE3
n1YwjT+7FXhi9unLHIf0EPIXlXQ9Uc5pjVFKIjVxY1LXXSnHJupXUkzVjHYn
Cge2+QNppL6VyQsMMReNtvb/Pu3o+QhzaOg+gCsVBWFhPp/+/esHP1zBYXRz
cwn8MZB4DE/0pCoyx5eiYX6k2XnCWO1+Y0vKVYJ1g1NlcG9eWAlrwh4miepH
In0MfT0ZKbb0hR5xk5plFEM66bKOjIU8ZkEelec84xvF7jFNUIsg+npgmIF+
sBHsxgIdl8Oyc9DVfM04wVQ7bQQIk9V/L8tRKz/I/BuyNOPipDynP/dJ3s1s
rqT8fzWmGV41SFZKjVvhn9vnzcBzYmbf2ObuxrfLHa8VmcgltGWjBXtnxri0
qR8Fd0jq6njp9Tc5rgOAnGT2Wzc1DuXcMasw3ueqQaEAH50/6wUOsSpZfRA2
nYFrpHw2LdYNG+iJu0XVS4AUHLxYRc1MFm80tWb3XCVCOuwm3vLF6g0JcmQg
yBnYqCw4yxwCQzPUylHMxLjZjVBMWRx8BWcMsifa7ym1+hKtw8+M5jywKWqM
l839lN4aZ95ITl9gXD1vjAxnxFlHlnqmO6UGLw7+fOKJcKXrDqtyFBGwo7KV
djzbU5aJVdnv2xCw6FLgN+GdOmeJI9JFevp/ehV9DMfzdj82rZUqbbTJeu8K
5Bma31uN6/NI9tFfZeglRVenqxtVP2Ke1oAOciarxqg0ozMgenc2sc9JlvnY
KlvutwOAThrMIQEzL6M+PaKzq85HrhWTo3G3GZhlS8GzuAU5Sj1onkhtdLAW
9DK70myI6RbEfb+Zr3hdG0QMHJRyDwM+E1UkS/rjdFcjc8LOkOkrH6OILZan
HId7ZExUZXlUEq9U2PBJmlJxtBrxu0PHptxy4lVePpVWvNk/F3Rr22Z1HS/H
XrYaBXhmYPFkgMyKkOWV9obdD3SNmsYp0Q94njuWDSGhYb1bUXSkIl9oferD
XHs6dtXrjQgAm+PcgDURIBGYZ1iJpnjNw1oA3WYzA4/wBtnACiHrmUdbjYxx
6+NrYwucQ+hw3YHMCWZZJ+VmVxtqKtJTLELkIsEMWuGAF8LuT71j+QGAVWGd
LlgXAfwX6wH7Ys89WW4nBD7D7rygwbtV/FkUyC0Uff7TW5Cze131xJRHtH/e
CQdj2mf4pY25hogZTRRC5zOGYQ5wbm7081lO2RQ6Gz6woMadwMr7G9kAqw2c
vdA05ti1WKeIk9+MloynGRhgg35Q/rsZmLSU4PkgqU/Gs6CV1WNnS1VmbQLG
SUuXPGJmWUOTxABGm2le+PLOX0NgjskhA0EcK5gXBMfFybYjljicCUD2p3FG
+WFSeihwxoX7YAUb5suW589E3ar3kSSuKnBJrF9ZiuXHm400pxu97ABTH9yl
pTlSbj+R7Mx14vnAYvybLD5XMH7MaJiGPV1AKxqCOiPI2JH7UlklyuzqrPnR
qOrpxpruhltdp3JccHCvzw2FQa4GYdZ4dfkurqf/TWT3AD52dlMZk/ya3XrH
aBmk68kIUYGAYfji7SRDwU2YAsWuhDw42vlhrbaIU6dGWYUtW8G7tn9xsyqi
9MZoODOV/MhptYr9exlZHLPfU/rpTfihWmAtHKpO/9d9ciSZfMTPKrACm7mo
nHGYZZQfEn/d5xo3JseF4LQ7wac6sYdOsYQrsd4gvrnnrMRmlVaJk6LqQl3g
xvdz2JDybYD6S0fjAjjq5YNMYUMx3IGxHznNsd0hBLrYx03c/o+OJVfk+26J
5FV0cl9vIrfP9QjHdSFxvktID2aXBahahHPsRpGLqixp/pj5tY+pt+Nx3ge3
oJMYJihHzku64SgqJ1xtuABGR6Llv0GYDwLmh4rolat9NAUxrB6iYEOMsnfb
b9IIPrzMLITTHSqGyU4a6TINyogabXap//yE2/QR5/86HFVDZ/vWFvl6UpWw
7/hO9snAYoww79VbtNg9CyLFx8L5Y8UO9SSXdnvk+UEmb8g85Rt510XwubMt
bNVPCb5G/NA3UbPN78n9EbdLeuSUcR6i3RLEVdret7jdvC1pqgMgPKYHipW5
A+EfKgYrdqQUxN/rkH3PEiRqd8vyVGFPN91QznqZh+Yq8vyO6RDHgM4i97E9
iq8tG10MkPtCGuw3auss6LlP+3FX4URd6TCtTidUn3e45fnXK3Z/X9e7vn6c
5hFjwVSx3KP7eE7ZDA8jjfJjNb244ClSaaOBBoKvNwgLh2pubN0eUi61pqwV
i1YHILygDg8MQMhnw6lCDVnWhwlffkokZknZ8CYfNoHsobZUyFP+8MNV8eAH
PCoESzWVr34rpNa/sEHbihdyE8VP6MzOpzW7zQ/x9vhSvEKOL7gtkSezePfX
Z9JN4mfOdj2XFed1n893Hqez+CAKcIlhyklCzb2UrzQnw5U/JZtFmAVc86yB
DfegQA/ORrui5lu3t6pMrE/L81n0IsXExjVuIV5RsVlx6hVgKTedpXiuIZQ9
12VDn4RJYqENTf9UIsdUhe9sGH9V8lU+eMMR7sBAxkgoDgtwySYPZa/08AGD
itLobZGKTQUf6FDZrisWtQgH6Th/WOWOMdO3ASgJMtyua9FrjLLAfRj+Mu/O
pGAwO86EkL1eNNrODeVcW//v9aH+rrefObp41NQ86CsxLYrwFsdTctONkQFd
Wk3p9Jg/y38CwQJfbMSO50j7+E325EhTjKsr5cb4dl58v5mqo2W8WmyOP5Us
EIlwnuxnW0LWkbVs6VSnW+Fo3NtQXIGNXiYNK3JRGDd9vx4ZnPWEVbykwRyB
McVb2MQ7sadUdtWSKWrpYBKEeXoq6/opWz7OSa1EbYUVeZiJl0PkaEZWSYvt
9FpP2IB2LSp0l95XjNnz1fBkwn5sloFCVfMYweVjMouolRRmmpuOvaQhrKqX
gPSrKiLK5d/zcRffM/ptz33OuFDPSjWdISIRYabppUkZjYNE+Ypiw2HSymti
cEKNlq7Vi7LDbDz4ZLU1H5xAXQuwW/eBpFqiNoKoAuwQsFGyHX91Z3gBpcyT
6XzVBR7oUb97UEg8d2we4mdaNHlIBa5agOWDxTmY4CVvXe+DMgHsaiW33bJo
Vzb7wqQZ+Z8ohV1xgoRYibmr91Uh6rFKygSYZalnwQZtkle5L+g631YFT6u6
YzUxbwGNP71q8y+1zchrMFvVQToXvirkUMCjI5npfGWlyBJdVbs2u+OHkI//
ZOOFi2pOjI2Ix1bMRXUItrwfS70m1+DiW67l6Xd8ra0SZWG+DNjnFcOc3LY7
af0R3zIh9ttsVPc/BCwRu6Q+0Gh4obse2nciH3VgPbH3PQAdbyLl6Jgb/pp5
hGXsyLBtZ1nDMGpby4sDw/z3ARKLgAejMTCkL5uwSAk5DTGfzonUR2PCkcnP
TLdpSx1VWAdHdtYIlXxbbeepwkp6qpeqnaPUZ3ycJZdFY51L3rX6ZGLrrv6B
mYbjLgVXQAneeDSJV49gErDFOAFEgmaqYntL/VdFpgOqu3COtXEOBdkyZ6U3
bZ9UGeQSZV5vuUQgtYcF1GW6keEe2lHoYU2JFVHlyqAI/YjcP8YCspzhLd1t
GehXE3ObgyxKEINJMERkU2G1RG+R4FUDuIqJ9qZmWYlCT8xpU4Bk1e7mzwZX
Sm5f8tD3QcLYaqAxVWMiyWoD/MgBUVsbPZklIuQddEG3b16dhRZHobB43g5L
uR/iVk/xmvhmyhtStHYjIx0sp6lB8YctxGdLGfgMcjCkA7uXrc/DjyT1FIYY
zZW45imY/hamoZjlFfPnbp7udVsPjHc5NJdi2EVTCA22jxk0QEK/LWbGwK95
FFMWGUSc/VmOxt4afdqwiG/uqbiaoQl5S4LVEAGi2MkMKqLu436XsGwtTqxn
vBDqqOsH778HKwMkYpSYdIv2nCpIoEK/aXXWz7HNBkuZ7/tDwsWC2uhvGQSC
kGO5QOME6/x1CYIrQQQxxUkgushN9ZzaG9A7zOMkxy4ZMkM6SQq3qzGn8K0W
L3xe4v4Lf6AKTuBfpiQ9mYZB1w0zQ/24INL8ryrONhqFf5/DX8/wMh/EVK+M
SaMXdsEosxyLedXbb2APqpYZXUYruz1yBt4MVYeCv8H5I91FtcFt+etKMkPI
Y5MGZbgRviXb0AMmQ4G9CZidj6O7qoAZWLUsl7AvyjiXGRk77mJMwt/tW7B0
9WroG/wF4gok+2bqquy5bZMOacN05JfBHPCNmpV7K/6V/NhvF6ZZGARbiYwl
XaqD4uHmAln7cOYLiI5K7SYdzR7kWzYrzoN49ny8H0Tc16yNi3RsPic4e4rh
b3mpUSlFad4ziQ+1ZOsMvGBc19P2uH84JdeEvrLzRNVR+MEXN1/zkgviuH78
TWzazTIYvzstN7q4zbJU9Rcq5Tkz6bFe75LhDUO1ejDyTwwWSAAxzrGspacG
hiLxpKmi04gcrlIeT2DrqR7FVXHTV64qTAB/7h1cb+Z46otJ+iIcXV2LJelN
ecroozbjaeMGKHyxDnlR0Yt3vrGNv98pvt0FQfEgKJFaneIrGcSIQv8HRXvL
pO2vlcljaTpge44fScad0AU/DEpRN52EfcLLEeupqU8QPuLPOKcCQJkHpZtS
uP/TVSo4urXfKX/whwZMSo1LsE41n65pgvG2ZbQpSGttlbh4T96XYeRwMGlA
PQtgUWDaTk7m1vl7eWp6XhXBeOVycW6SAuz8fMAtrw2RrlK7oiOjqE/W1bDD
X7B0awylFgbRbOdEjnKk0fKvahD45Z6iUlNJQO96z3Zda8c5lyqMMh1Es60R
nMHmuiZn69Ji6o6ll4eg8wj4INrr9613eMEvT0e6CotEGP+h+ufp/W22mjaR
uYN/a9shtMJht7Mk0Uzpvjf95Kdt0uRyM0rf5JTMNgBAutx+uiVOzfUc2myn
eEAwDmDAdgF/KHXMOFYYl5gNHtntNolmV1m2ZZ2b3jo9WwG1qR3pQbJpe99k
pm8CzW9tKRpAITD/dQiYYV5i3NRZ0QfBXw2LsdNjHB7O4++9unfCNAPIvy5a
dXk+agjnsF7IXOeZ+LmQ/RsBWRqZYrkZ+FD//t0DS3nJcb+zy2D9fADp/85N
37a3ZJJBZSjADj/fmOYHuymdAq9BD1Y7JJHFB5w4qPrqAgVW8nkRlDNKVJNH
F5Yd/Up4Mh4d35VGqxhYtu5ddgXiZ4p3fhc5elMIbnt3jtD6XfO2jd5DzFYF
wzQJWsDa57B9UPMT5XQ4Wa2DJX2jLYvpSEz/FhgiurKXn6PsawetK2tGGika
y5SWvswG6KhJA5Q9UPC6CfWVFQGZ6laMgcygdrw0svnOeKuxJv8tN7nF8siq
nlxTKWm2xWJvAuU0tmOgaPlwelB2VPWu1Ds2ceOBUt4zratHvB6YOuW4gVSW
/fnb9wj64CeL2xcegFs2VrkU7uUKEejfSvaX+pM4hAsGnMKDI/oFSnqZtpw3
d4xH+whXoCNNTpQo0ZsNO5nqUInHaVNSQ3iPPfGuXVv+6XatL08jTymrtLex
coTdAG5PVTovE0N6h8WjHyLXiRhPA9B/3ytZCVozLOLUM9IJM72+R9ORAjQc
kahW/BbJ/h6CuNQDRk8SS5ZPOc9YeM4CnT3CEhZeSlNoOPEJhMQSjfcjcR9a
PUn8gXyB3HaUp8HILWFmlxnM+o/oQ/do+wx05RwDbbdnfZspETvtbd35NqHb
kPcjNNL6JCfNiJy3slSiWGelN68xV3EzXYZPrgRlPwDhMuTiz0BsC1A9Bqvs
xJa4cANYRs+KVU3Dl22auat1e9XbrNpYQC81f2+vzjZNTnaFQxaJv7vztwHn
gmX45ZncxODd5RTQoI9D4bN5nZ6AuSqVTmhc4uDa93GUlDgNgkh0vB26A+wW
4ArvEqUaiCV8IWiIvGw+N2yCJHm0MHAY4///gA1M4pmX2MUbO/PKZVqS7PRY
SUBGMxadIIQ21KG1nnAut8Yw/vNmX/0fTgqchuerngjbNHgpuL0KicMmgKwU
IJq8/zvJi/KY3KIsESQehNQvdimVKbg34n4J78ogVdNIGzlxeAXY6pTexH74
LWVBGAH3r/NI378Ck4YGxfyANvVmVcMS2cYMFyMvdj7SD2KimcH5R1jjmwSv
7keg96TbHknP0ZrCWVWiDD8n8LHYyDIM/95pq4NSnJZ/8Ov4FOUYhAZ3NzYE
O7/RcEfFKU1gR02MA1Nzu9NPnRmoeqc8u+7AgUiVw+uzpfnh8GqtWDZs5gTO
fYipi3R0Brjg1Rf6MkGKFHou2riz53BpSiWMkHhQOaIFJGwIFuFj8TMxgzOM
CllnvkLarwmZGglpYoNPmTHjIeZakcRSkNEKLx1NZPbiIwD7mZfLjngKeHzL
ZIC1qydDbu+6X7NDXc+XwUxMQhAR/rDzzThia6tpQoif71VyAvcf5zLIAFK7
7BxzVNQsex9dUT+HB4gv8qNSlGDP1TY0NChyNpCAnKO0hftZ6Rd6G1Alp87A
yiNPv3WatmV1SKo2nF1bKGQYb/WJw3r1i9MatW55Cjasi1dMtr/aQ+ZL62Hu
MWKWXx9p17ESEeX/PbcbJ3UaWuqCQ+lvov6R/rPv6MP/G5wEIJ8rlVw+nCtP
ub9VEWpJxvNaAdidtuegR828sJgThBhTzz7ebOgbh03g7o7oR+0gEecDkxHz
suTT4nx2X7YheW0S2+84BXBnFFyPpGoILD9m2Ao8gBnb8R2Fyf3w8U3Od9xX
/9hAja7ztiuyHMJr9nIRPY57D+btROB2GNhFpp016UqMO4dUUaGle+zbh2FB
4IaNPQe3UlubhC4RH+qXR9YJMFUUNm9cXWFqJWhDmZEYtJsxCQhAcp0pfQ24
2egHEyRwTdgTGucGmb3fieItRgSgHgI5Ww6xLyFzJoHUxiGQmEkHqzbHNZl1
lnGDQuXImLvilCt5fio+gzWsU8j1qiR0UTtNWU2CkdJ0KurLO9FpHI2RDMYG
6zUMXi5QtmTehgQd7vQOn1U32Bq/y8l8cZ3CZSFEDE2MdLFqz+5fhWpoBOSF
lNszfp0ARx/lImJXbjoV+W1ZoeJhmfY7V3JLxwFCkKvQDl5uLOa/yeUzN7bB
h/E0N5J5bBJcrUN+ABZXUvULs6lsLA5IZYwNG1dnh8JjRm3ISY/Zc4v+6arG
QoFkUroTrpWQZQ3uhGTZubfu0PnIM6jxR4BwH3BWWl5cPiIgeTkJyk69CL9K
kURkHBHER/L75arDLhB7Gag8z5XUDSxrf4+0B/OlgdbBNTRFreLltPD+mCKc
WPv1jgiqAjhOhdtx5COMaYp3bUOGUyJWDBNhozqFnu9ntSajtnCpNB6OCR0Z
1RVk0KEhSDhKQHm4SCAKBDNIRSu5XjYb0AS61BXIJ8lLBXUv69AjNicpUKuC
c0FXEg6qnzLZyh+FbiXrI7kzesn8kGfKRTEhus1uJJWo2sXfBLMmPD4C/xPr
WV4O7m5hBZepAk6dIrtQNB9saHZTJisSYV9HDHhX3izvjlF72fnRqU6HrTE0
VkpDICvt91pdjv8yyP42ZhR/+GZDTgZN3RLUJS43OXgNalKrSm+193FzJxRD
rRXLmWkH7qLugXDo7XUJOZ9KgQx1wtQKEw8q7tE+A1LnMhum4Dx07Eto+kca
lnUJAbZvkO5e9eJHqRyogmBPkkOAUf/7MsMCAu4Sz9xvXn8iU/4iBkzgQyxU
jFIFr3OVhkPnqGs/G5sDnBGehx72bz4ydsFtD8uDmgpuSe5Ec8muG38FcxMJ
AEhLvW/hhFt+JpfrEqpvI4HQQszSf5GtXrGJMM0vQScR3vhpJspdoseRhWJz
ozZ9SSuRQZ3YMPNxgVxAVG6+uTfQlvguMs2E1wDGgEY9hLI+tVbAJUr7HBs6
wftDLggveACfwe2TOf8Vrv/2+aWDAdHcIBd5RTOGOdNgRjXg2Sn5dULzDgA3
dTA485HDLnnXIBybjfz7g2NdrzqI6+qjufsfGu6v/LJaKbxOPaC3h284fR1R
oyHqE5LAu1f/lKLtcJxwQLqN8U6YmZSfkXLhQ1Iq9+XmzzTFjseQCpzydN4k
XW4SiONUfMAgi5UWZxnIsMpzg7MgckdMUKO2rCTUnNMJPwV5wEznhJyAvGhf
1rkXkEKCfjfjMY+3zfqrDpSeTTi2jhl7k3vusAwhS1NH4o1fa4NYXqZrlWNI
JhN2b2638xCq1N6Db/YMK0XvGjtxtV6aXu1MZyQ1lNwqXloVt8KGd6gUw8Wz
NorIeLQ4jsiRT93Tixu7nAC5IStFYJiTCoUGMcFfxpsUuB9vTkg6OnI43OUK
r1vAZG1RJnhzYk9rKpyFWFCRBPbcoOfL3l1mvjirsIktXTsA3hmJy+KxUN54
A6jPxAV8H6z65MDMxjJ3fgaUFEzuTeiCp+OPoANVSzevciNi9EE2/yBIxlGV
SuVDguOyI5XDmmvpeTNRn86INWL8KsboGrjpOlLXV3fJhUkmp6WeP5Z4Joy2
kOd7cmIZXm2A6S5vpyakEFzTqYxlr8IHw/cRdQsld4IrWVEPt1mgyGgOfvhi
4ETed7rKkXKxSPjmCEX0pw/kfmBEcZJFzZZOymxuj+3AJMiXOGzkaKTjr4ED
P+gmJz8av+lNVBryWyEyKQjbghfjXI0toSEhC3ngXWx6QYwN76F7kPlsIYsW
08de4YM4CuiBfWv+Hza8dQlG8faBOhDHqZftp3tsBy4Ik4IvfCTNZKV9FET/
0q9QY3/xClliQvuTmIN+t+KbjuDW8Rfkl9DFVnJZOypp9DTia5gDaAPATNVZ
aXtEGg7kcbjnB0/aPllAEutxla1MqMvCdJ1CO2DapKNM2WBLLurJ6nMOBLPW
4EeGoRIUuQduf0sRCM7LgKpUFuUC7v1fPXkohQ4qVSe8IHMRjxgKemfDIFxP
CESS4ovoSfPIjCCMVIQ22bpLLplnllNJhdWbmdXrG0WyLlNZn8HnnxjBiqbP
mXq6SpyBop4v8caaL1egmBlvEpZU6DO6s5pQxhCxaSWfcpVt9OaoVgphey2U
Lq4IUKcGd4cK20vHuw/rW6PyEz5DILdGy37NrWhBQcwO3nWUCRsCE+ht892x
gcXsfX0vEXwLFlQwPNFLEzGdqK7D2lRe1OLHF7uGUamz8Evwys3DzbT3v8xD
LgXL8dvpO1ju8AsbHFCWS1Z5b87bK4CxWAQgbKKKLhYPIcaLZGy27RnlS+i9
Iqq/SDlN7Znb2YlhJwOSGwUAcRJazOheNkB7qXSqlK9eqVxXJD56pPK//l2o
kC8U+2JJt8eF8N+8egIDEfHHNy7bkcTvGhDPTo8ysoqp9fsTsUscXSXCiiO5
KY7kLvzyPb12kgl0ejFHHBLFNs5n2Xyf1HpciUyAJktKzCBnKVFCa0hwZhbY
jzbduF3wbG93XjmuNinYI5gfQ4MOrpv+igiGvx8b7S2IIgl+MHtKana8qJkr
O8xeCPhxfmbnCMWrMiGIYp/9rz+FfKDRaLUALQt6aXVeJbPcCGWFDxUxczya
mpfa7y4J8tP5qyo1leFYli7pGmGOQzNzChJyi2Z+Hf2I3Jo0XmAVHUHOTGib
5P/pFG88GuJN+dK4qxmfbSbehU5nUsummXOkEAwCaX+sYcWG58j20m3Ti0AD
DJIZW3pfCSR3vuIlenrq9h+WlPnVuxNL5IiU0W/CrpbNXghbVcJ0p+Mg7r0U
tNhGiPkqbhmmv7o4fpePAvXGfxKsY+KM0L5sJHyWv/UVOp1TmscbmNYCasSr
AKQWHG9JRiPF3w0xd5Qjm7CD8OoGtudtVD3Q00fzLZQVXszsi+55wmDP8CDE
NR6sl+hBcQS2EJnrLNs9TozfxLjvPgYrcrrYMBnsYLVAkEGMTEmYlC7lK3j4
s2Wk1jdPfQ/Yzm+yQF6rgPbU64jPTtGnEPR8xpvLIzNZYOmZApvBvdi84b0r
iqszzDdPj/6j+s+2lWodkGjXFU7cjdgDCKgTXaF284tpXtpBPFcSFfCxJfoa
AJGEdAXEvL4ZFFAEp+Wiqc0QQ+MooG40c1GcTQSElOIWADrsqsHIZr/byCb5
BWJK8Yrt1dIcE6OXMQYdlcA4QaAZEhnTdibblZ2r5QqFI0hJkXRUyyJJV8vc
7GvvMjZeSFsyonCqiFsZzBS7hlH6aY0RrbVf3OlLpmxwibQilH6nsUk4Tqxd
JQFAIc2cNiHSUCRCrhAt1rbUVXd/N55LFK/0Z2g94XDS4BewA1zJ1ZgFQUG3
BJxuprVFIMg6E6lwrWi232ofhLWoTxoCzTShgjGJvANRYBZngINJgjxGNd62
NwXR7FIc3pJdSUrToRsZbIVGzqHvMrpZFgFYU9GSC+6ZzzsqxW2B6axG1Wk2
sLZgMIQ0Yv9beFsX49Tp19G0NSV9j9dvlN1Ykuro+zxr5rAxoL/NhyiciS7f
KFPwcLE5jgng8+agkbwCL8Qx2BgnwyKz+Etf1w26Ob0PRQsdyBiBclVwAxtB
vUwZyfGW17bQEI/xde8GKgT9NLJPUYBQAbD02ewPAo61LFsVcenTQ+iuQrLJ
9KLnHlKGejmh9VrhIpxyBcwUr3LG7MnRhCx40VE4HHiq1jaYtfxkDpba/9jd
Ex45tqUX5voTgqnWDrxHiKSXY1WV+hRXZ3UcGNa92gqOYRLZ+dEIfUx7rNpa
jmNT5DdXxeGmduggWNxwG8pxFzKLzNBU3XXkoY05VXMlg32pZXxaTvU2dLaE
Tub5nJJepfbbm4Teck8TIUidd31TLSh750nwAmhW2/PBsSwPOI5X5B4u1VKO
E961ek4Me15FG45dRiUB4GQUDIPDeQ0nQua2ivp4xAHvbyk5sS/JN4QFDihb
ogVHJgbZB/1+mhBEfIQPSn1xa9jPMAXhN/7P0I1QwL27FtD/K2vRUB3DgtzU
jjGxuLM/sPQPKmnp6UF/A1ieQJLkTtVaki8+SK+nLJmp3xzz9CvJvHsRN0jo
8rhHRg/Q//j1D5Vrs1sP0OXmAAY3jPoPf+idR7QUopLT5+cSeT+b2gioNuys
xbzNeNq3MBBmqwRBsQJSQyauE+CrEDeLVPpvDguMn0HZ3bsyGret+8AQOKdd
5g4wvMCS7TKs+4JAexL9EdE75eIA0yH5Vn3HkOphiU0qtW0iqFLXTgyMq4+p
Omatf3FqmS/3XFY6/eqbP983Ye7INGQzfU15kMupexpfwn/pnB4ESGAIIima
/z1sWB63OHRF+Ogi0dJRnaB2CgvfS6wzO0yvW6uPKn2hGsxYeMijcZ1vhpmj
i/Ox/FutujZG57OQkL8gM5dASc6XCLZqR2Tz29Mf46UsT5ZPMSeiyI1l/Etd
VsG7V4p4s8cwvjQd7mJDpxRxpBqbCLpb6fYkD66mKI/FZBeNd7l1R2aZF3+q
XmOI6aYT/lF0a/JsWvVrdZQ1/d1qrLh8ih98t7SPh6BTz29YNMqaV3S7gIKQ
wi+Z6XpFCZ7/eqOn0sLCDp+xaRyAOcvXgBdMXTz3GNR0cCgd6Dc9qL+JsY1e
ChLSDDHA/EUHK9+Uvl5moM0QkY0bcPOQZRwQ4V7t/GV/SqEVD3MYliivSdQt
6T5bbKAFfE/IYMZ4jDdif+ImsES3VfBh6ojMcp1Z4umzV8V6uhsix7HMWMIa
CVag6tJYTPap3gcBUR47vgMushPlIbQYf0JJqgbSki5Y+bgsraDxpZiKquvn
JeMWotAErJOQfvNouUVeImctPMgIx03BYb6roiePe4yJK4TAtotMyQt7HlI1
0vmdXIE7dR6PY6HWx97ALqUegMAuwnVEQOTZXxTyLBjYKkLinoy64z1v0ywz
ucDhDZY5VAcnC8cTUbGEPcLUXOAx4cHNK6BP1eua4P7K1qaEEud9t9cVST6x
Vi/jh/1TmNDIqFP+N1uRj8IDLCGkQrRC/k6rlg0tR6RzlTLec074Hq02tCQ6
nsRBTJj9XsEvkabgnf1RKgMao11E6eA8MwhFQdNKb1YCyrIkdEvkw+DSRaMN
zVhmEBPJTVnSvCOufAOAbmUQH01u0PvpCq6Y6lj9GGFahCsx67jOM6XQblKw
uuIBeQ1leeCxp2RM46hRnIFVPh3yLl27bDCTkIuRJzDSmCK6IoZH7VIILtWs
SFPuh3cNpY5Ncb5yoAnzGqtBdvY15PJw10olXqUN/6QNqbl28C5O4M49ViX/
H1KMi9vLqK8YPpf77KyMNcP14xSth8y55P4C5lGgN/ait3KPnyT85T4YuLFX
JsxjSpLjDXfSPtmSBMmif4N6O4iwpk425xW0o8kzMQAXhGCQddD9NBZyJ58A
W2KNbH7Q36Lo07UsZViMkf1xGmiq4XVRoKpVFKLh7/HPL7w0+Q3gTVX0H4XB
rU8qMzQL534h1D/grLGDrzxAe5l6nS9q0Nigfxs736OS7L//wRLXBYUYjxMN
BenLJt0opq4xDkd04hBB2cD8Ex9VJxeGu07JYd25U4H/EbW8rifqMQ2xnnbE
VAkdn9sOwjoqY+dbLkYzQPy7Oo8C8mj1epKFG6jLYNgM8hHGF+duJ7ZNIzMT
slKrhyv4pr74pUHcF79mbCTyDbNxTRtm4EBApDg35urW7/HPNimuMo5KT4hv
Yiy/8Z3sYtSD6Pm2hihN7QqSeyTX54S2Z93z7HPB7Wzyh1S1FlJcg4l4ZsX0
ls4p6UwN65kHAz8lH7Qpd11NzidOXcgG+CUrScG5EZPQDcB5/GNcwF98/9va
D43c90SRu6jkUHTq1hYQIiDC9dZqVS2yUz4lTQvfIQXIunhORALi4tprUTp+
eWzh7a1ucMvjnRSoEWNWYaAyxUSvwdlJECmh5D7LH8itI1ymgp2VolHFJuc1
90CySQU73e9lTtFcTO8XSU2I+8/murKWrPR9D91WX+vRxvB3S+SZ07Sclho2
1hjqcUfb0RRitwIBlUwT/78FQetYY8L5urL2T93+LrPkNcjvbrqLHoh5Pmtq
65KqTU9FxLIK37thI9uXslZ5KwX07guJ0d5YuA56Ykn1XTY/lUgSUG7c8aF4
60x4aiKoRKl2TZ0ZZvl/99NxBu/CR84TUot+yXqmw5VJ66tzCLwW7U1+Pi52
pgeWL08cAQaeWp17yqrY8Nv7I3G7t/moS7TiD2nO+9hn33iX9X6E/sRDbg8z
4XeY6jqrNvNwmLK6smnPgVMJ4OZdYCYAbECuAxThUI/1mXyENq0M/1yea2cf
jPb6I0UxRNaWLAtC5KowbWqbO8ZhJ2AlcN8cMX2reVxVeLpntkvgdrtgteq0
R815mfb1FOTCvRxk8vXXx8dc/3FdvVZqTvH3iB81651YI39SPqiuha07447z
pxvp/GUq+3uHfK3kRlJyZ+Icu3HqA4+L5jlGwH30sYlhPDlQbLEt6ACTXHf4
hdasIT1jTwLTOUDgMzTZWunRkyyPoljr6mN/6TsIxE7QuvfjZPthTf6rgff4
d+trPljxaGEx/k1R4X6nbDUGswbvbJ7fR1HkSjQWzMm42VLmNetqLe8sEOW3
9ibu3KpCdCdtyeN1wQLxM+j7zGqZoPx48zk6jR+qKJL1EcI05IiL3DGRxJPj
ySuisxvElrBvH6/5MtGg6QggZtrKeqQxSrTgIyDsAVHhEQvwRejSpamLyrys
f554/5zxbiMA7mrPs6MNu+W5U8Cyy9721OxKJCtz3kQlNnj8HF66QmZTRDzF
Ltzjg2Liptg9KIiIYRwYYp26R9D/ntl5VVzjm3YYnxIU9B9notgT0gd5sgA1
hzd3ON3X+elsXRDLAQZhGN+dtFEYw6hkvry1G+sOoMhqM05JsiIng2HP0hnX
zeLqJhHCtYa4T74Nw9PsvD8qwCJrV5djOH4g7L3FNeSkARDEfKec0n5qQxQS
kXrDF3iBPOpfqpGDTkvSu7wYe4PZiLP7V2j4jj9wIWksIKYCZl9vH0V4J62D
QyQ/4SjdL0H+52HYQGV6I1lBpjtNv1/bOIlFHkF2+/T8Zk93uaNQZomjuIQS
4mH6UnxGSYIxxoo4orFqn+52x5Kkr3whaKL2tj7nFMdwcua7ymFB+14Flb72
yMgxqXaU+ygAXTcyGv8NPxPFMM1GEcp3w3anagFpSN8vbgFqDSocjeFWFHdS
p+8l2nB2XiTjCvDUwzTZA3FGISKRcGYf/ALW7yggfbOEKtpiN7P1SCRLvrUI
+3JEbCNzx7Zlq74Bq7wko43nVFm/BGHD3BixMu6IhYUPbHUXYbDEYBE1wrer
HhUVwMG9wFpmT/TmnpyvESTCFeV91V/b2Oj4NSbEcubOibnD+bg8IG9QHJ++
Evo9ltskb79ShSnCKepUB/ZIqkcu3gBsJA3Hpp5D/W2xfkC5RbmXcoZ/2YQH
zinHuItMhEcvdlIFiQ2JTAZFRiBhhNTTCrI8O/kmSsdeM2z8OYtrOulbyF13
ecpXjkqvGz9LwZ3mK5uKPxNY8dgXLoEPvLbqJi05eQ9sig4/7US7Q2m4BXBq
UW5hGCL2I91R70LnPTdHMmBgp2iI+ax91srrVhxcXBmmoN8unhQkrHVSw6gk
E3gQb+jaSTR5qBml0SjmdXxCdTZZvsJzulKKC41Nj/4q8T3D/bR010Px9utZ
RQJ0AwzlgH1S7R8EWnowZcuhU619903eW6Y4aGSYeFVHn2o7s2R0//j2kh56
V5nLPS5LqlQZtu0RN/K3MELQxc4i683YliDmRbkVROQC0yZ6i0g32Uc5pzpc
yr5V69JEQLFksUBc+VTl0ZKkQQdXaNUHFBMBVE9R3mnF44ag3nkZvU2I7HDY
Zpa41a2W229Agvo7QTdkwb7uFN0DZkFwTZ2m11exx2x/atjTf2ahEe1QzLEH
g+g4He6TCt8GivyBRaqvFj0g1KuVJ4jnGHzsLpCwwbSHaUWRbGWOcXVHOms7
dvJDYjr8YMB8HFEnAw2iBeMzKDMxxo+f7B0iq9USHdSVJAjj9t/7smvfrbjs
0F3i6dgddMxPghU+teilxza3hkWWEbWD8OtMDcuPGfZujxN3BHeB92CwriNO
OPX6D4RBf6Fn3XwF3C7M7kIQEkT9JFbprdYpMt90dgejej05GSzsqvALITQy
oy3DUjNHJMnkCRUmolz8lWkP+QtiXfgRm2KFhjUnG+bNlWZKEtGiXy9rixLA
QD5H3/8DzfZ3BIRy6zHxhyQdufFLHUBmtLqzRK7PAxzmLQ0GPFOmVdq6QBBE
oK1SFBEaECK0nF0Dj8STZBLpCAeKGmBz7qrE8Uur5FnKij6Bx3mCaJmONhXL
F5qaoxIUJAO9MnQTEip3HmvoPC9TKQM3+y/ySDhwh4WI/tw/OPcTa9Buo/v9
Rg5C+FYvauRVFRSXj23VX1o6KImORvtiv6OsmLk8YXqfBXrWlskqtwWp08ko
caUQW3x4b6+HAKPTd63LQ7wPqDDKgLGvJf9tbTvWAkpVp5RQqxOfPTk5rrGm
fygSoD2xdrsRTFVOfmT36vm5iObW+ImNkihB+t55bRPdpJTtQPe/yhzemxSL
fB3CFcZmwWI31+EQw2CIfNFxy/AmhFejq+Yp6OrqOTW5aOI03LQXoPwgyTfX
oP63tWUKvAyMJBaOwlSQ9mScyrcD7nmK7xGsy/e3E66HfUbSdoPAmpLw5cAh
9TPqdrfJhjJMpbomgE7gKcO81fV4u91I4B3fhoknzhIDDf7fBAcY1PiCyeEO
rS6WvDJPPhQQSHS11K0ZBrTkUSV0TMvtNKzTUZkco0W1OaHRsYCHVmkjaD3C
eaHp9opKZCMAh7yqkteUc8/MN/EgkgBSfItbPgfi9DWKdUlsbipFuXsTSAb5
TWbvqdTA5DDQGIwlFHaFfmCr2PT9xxOJXHtLJL7IwrQ96L1isEJmvFQrRapx
zbdDGOI+1qXbmefqM4YEUmRec6PGseIjymbxAYohuEm7UBGfJicq9f0oooAd
H9++FhrX4Q8FSZWz/z/vtf9TL2yXDVz03foXbOpqHMwyKOFg2GydT06XLKt4
nAb0rso/5mjrdSVElNotHVxnMEl0zIEd6m6JHQAocZSv2PUm0YIoy6oPgkf6
I8LsdWdxIAQJMH12T3DXw/Pn/w5/Oi5mP3AICd8TiRC62TC+Oe+jcL/82s3G
YlL41Mf2vt1IUB4T7y9I237+hCy6QOOMYxHChEBoVmP+68aPLAE3LVl/CnKF
egxiIvOvEJeulGHKjz+DYjW5tt018wgXWK6+I4X9iRjYSTxlrXo2bNTVXQBs
HyQVkDfXayDDRAKOiqEwvve55PzU7Z8QSouIIP9NIp4pOqXZeoyNuKiXM8P2
CAvBv6cg9U1uUM19Eoh3suIzvmvta/twJKhjtq+qDPTUnqna4sv4G3CaRjd8
4jfeMZ4OQreGsjbSpIkVBn1potgKTyE1TR5vlsFtVTlqbT0ZFi3CBnv6pRGg
aVlWBNVAA9YmCUNDAUQlcPsWWouJYHPsKz94169YXyOIiNSsgr+626ox+Pw3
5oNnkxlDR+lNx1zoMcdB9gX+TwRBLYT5exwpTuAHbocdRh+JGIAgWLB66Pef
DBL5XfU94SOFwqXoUqpwlrLFJ0tRyq440l5KSjdaZoFpndKaCV61rSpABcuv
kKnWOq20MyE1PXq8A1dfzBOfoFTtbrtbYr2V3UuD7Nk0s795iUkHEs2/jKWc
pEYxbg/vMbZ7Fn3c9Xb3utMU3iTKqj4HMXFkOLZvHe4otNpu5lrGSXniOni5
EuD2YlKjrd2trv1rezyGozbn657NAsHTENvh2Jc88Yf/afMFGXlZB8Ha3m7r
aoDa740FCSODJBP7ATCX3Q9QnjNhPZNrWH3Wb9I0P6goYn14IV3+GBguwEYA
DiRV3KIeQ9lpUAUHS9zgtz5Kic98zAMLIEA7wg/f+skaOZjU4yPAcATULTpY
LqiLBxWfbZXmGmE3ueZtP39ClO+dr2dSrS5t1UAAY2+m12J+SEiL6E9kc/Kp
X0O1COXTAZ7N86Ks1jCeII30Uvfv+V6sxlBZXnxuajBZXTO699J0FQJUvoZg
raYE0MLi3vWutiGSVVXTXXLsUlckPauYvwecl28ArPqCspSQlHgfX+3T5+FN
j4y/fK+euYyDqlb3chJp9QVOzw9L7ymJiPm8W5n3vNgrAQPRmkbzw1/WXkCo
7YwQAT4Vz1Al068KSRBTCRxZywPhYJSLTadaVMRKSMY1jEByFhWCWp1Q8wRu
pnIHGbePoCT9d9AX68+ps/OKzVfn0tZA6jD5o5k+/jH/DxY328j1WNErmCC0
dCj9fDecoKLvTUWGTWzQqkieFk1g8EU6BaSC3ZYtiUQHYwA3QwljFNkPi+7+
tBbefkBDQ6ZSo8t9LWgua+MaRK+VMcdtDRMi3Pix5efWVp2vIHHwmp5l5fmT
x2bronBN8zt18OlEgejwkGukFEFrYCJL0mNX1P8JL/5P5D4K2E6Fz8kyE3Of
DiADxJ+ZIs2zMk8oLSbvhdNj4eCfSuHpvl6+eTawdxYQes63IN0W/VlhsfiF
c+q2Qn9f3qoLPwxaEo2vvj9A4Teh/inULD8INLGCoxl28HNt/ZITpKh4iEx4
fCIb7CqrIwrt8RZZvyRxYc0QTSuhPp8Dfst9NnxR6Y2XIH68+wmDax/3XwGz
fGhcW1gr+Uv6xQmWj9n58pwb2ngOwmscG1t6I96QG0qZF4Ot+CE1b198RQ8G
0mJa/s7deBJUMGa8RxlW092deusTCqq4EWpQFFl90t6BdPkcHxAM7daknX9p
jMbsdEAk6ADrFjbdDXXLD4CRAlEfUWCYHeLaEcDc3V/N2CprJcW8TVpYGYcg
uNK7pQUZwA2xhIpufJMQVbo3FSQZTLVyEwlerEvrwycp/9C9EQZee4Jc1GkJ
qNuc4wIcurEsBtPY/KjLyi9Sew9G5RMitg/Rz2kczBuyTXl8W0xTm0f9mVpN
H5cOgHXRdB4mX0bjUQ8stpbSw4EvfuapIFwiaSDn7mxBuW3Tgs7y7r5rdD4d
wQrvbOYwzwG6xC3AxXCBTI2McAKuHSMv57JDe6yIaKrAszGx7spEH01NA0TA
v2I963sZEIFhjjF68xAMOLu06BozLL9NS/qnHmkzzZvMq7NhTi7XktMbBnJI
1VbsJtbmhRfw7cto53DyLCBU+nGvOijtCJQJcAf89gHq3Vh/ySQuIGrMm6yj
SJi9QmTpNwuRxnwFFNcEfKGK7rw4ImxAlOUr6k6ALeHSieAaa8z3FkWDcC4O
eklQXHXUp24l9Kjpzc4XiUUeCi4i6JJda+KANRB+JrVNOoOPM8CaCx/THj48
eoBomDpgyam3zePVhFV/ZOu59JkqdUY4ujxBzkzfRkyXrocy2pA0cvBFQrTc
CuArBimeYkZuIpBVC6RtKP+NR/L0Iuw6auDGZHRdvf7CQYHf1QniQNmHoNe7
/YaB6i1mQ/vdrvL51taocTqA0lpIwysiCipPJQYuNxQX0Ij6Ogb6dNoB6pDk
SnP4UuTgCtmJjgUltrPOvNxT3FuMmfygGiN/hNbYsw6C8qlWm/Y9LLB1xbnf
OILfRUAAYIxs6iQbm4lVegFRQtFbaLzi355DRyFMGqFZ4cniHw0FpYopOuXV
A5n6Nkk+9+fqC/aSHnrwAe+e/fvUWrnIdzRI8GV9C/hXdPNeYVoCQ3fkgcwa
W3N7hVMqqzdVS8tVWrkQGl9cOtFB1xphnZNy8dk54eWYXsfizosrbLBL4XET
vaMDNJcW0tMuD8sPWhqmzOPoEJE54hbPOwQ6ybEVq3c3sVSjikZLHsLbbmp3
eLV+iETCG3PcI/UPOIEcsm6ThCeLWyoXbbMtPRKfw47XNrwakXfBoJc1jSSb
x+S2eypBY4dFZZ7zHQnV6ici8PdlTpmOLHlaYwpCIDVB/FO58mNQ3unFWAqD
jd2a6AMewoXcOt72e7VimSyc5Z6EETSzEMCWslntwf19fyeEoNHZkef5k7id
7nZqcXLbEBKI93V8pGZSrCmClehHieUAgANLpoeC3CotAxhZ/ICMgqn8Wlfa
H97Gnl9/tojJz82AUFRc1w6M6E9PRDaB4ukF7loHfwf4fJGzrc7IO4o8iyfG
jq4+IH2Ov+58UhuSrAgROesIxBDq6SMexQGzRVV7JV9jGnEluQynuzinCB70
oUAJROzvGSCmpbrhYxcjsYHvxxzhgikKyDSeg0ROI18ZbHGiqTOt+fuX6d4k
iJCLS4V+il7Id18+NsfIDJhLBssaHrQR0TnwQtyreANeNsowCZXnf9rntt7X
02c5pCl74uTLDu1Xif7nuMt1UKQrwPI9iEJlDB6acJ4W7CJo/jfkRAWRVs98
PpN2JpN1HfydKFKBmOrVhvDLp7NcPEnQFz8zVPixdg6YKwAYGaPCNOXeyy2a
wxWV+DalNSxQDKbYSidtKKI6XUJAYn1hUDbFJDJdiyOTEP7C5nyWsW83arX7
SctI9dozhYhj71O7sMJjaTVUyTzGnoycItwgxQ5e5FuvajO1nF9x+4WzZgjl
4BQS8R5wwfQC/pO6txTzGwXIMxqNQA+vYMbHAnKHvUn2TDybyufg9otR3jrY
/row1p7pwym6dlnlKiSqaqiK7AdSzBj3rw5Eo1hvHcIGYzN+fer0l+OTqfJy
fsG8wUQ7mxOmOEfN6vAvU1wo9l8VQqk1ruHfQC+2QH4r8NnERaliyouV31PP
IWW1OAMXLE+pTByV0Ad+qxNqiO4qXj2a7c9e1733ClQt404ISY2JyesG217Z
NH7SAmdi4l0+aQSEneIWYerH7eGTxCRvpFt/wHqw8m/9K7CUgT32c8vJozpo
IuVMMAZmZd8gJXjMBKatwazdNhA2OBhNqEBfoVyBqIMasCN1zN6Es/BMS8JP
qscbQ73dUGfbHMo+5PvHl2HcqjN8JG8c2ynSuHbcWU1b1vjd25aLd1sn0ggI
JdRvk4QGD/ZCU8YSL96Td5AQSZZlNhS0VSgWAfiEgDFCX9gA/uwJXHpxq9WV
uq4grwj+jJPzKa3lVVqTw9DwmqIgdpHL1aI2LO013nCPFXDnfeeZTcoVnwQj
9QQStfuk3CuaWT+7c5nzzo1lk/fOiODLs6E2+yuEzwMzX7vO2SD4ct2xSz9d
Rv2/DUIEgSXVgb5MP94aTp74GgTNNtELkG8lqXU5YJqg53UjTfWUd+HiJQXt
dVmnFWxdDc8MeWutLwuvg05g603WWM7BQzKR1/7bI1vJUSA+eQy1dZTgRogd
3JFz8oqkaSO2jqxHTdnUKats7VTCiadiMg4kqWRd/9Fj3u5wf0Tk++k9J59O
C+cfkYF2ZfDN67g/4ae5gxwkkqFmIb9581/48oJ87tbuonVV3cZxHGUMTNDK
zaZqlONxbsEi2xIZWLmYRp+3iEpCteeyBjlGavEQ1PTipcUDY97Z6PtQTFOc
qH1dy7WVj1VFkHnN51hjnGg1wM9lHTwpOqiLCJopesQg/+DQlcV2FSMWSXbQ
QtmCEhbCyyB7SITnpVFikoPdPy7dc2ahmnNKGD/03cTp+gJ7BQRnZq0/dmM+
jht6rfrfF30R3sjVkr9ofusUX775qv5D0iNSPg7hRqLLaJHI9dKtxvY9sAO+
iXzyUnR/MJYEdBThSWmp+nH57Ic3+GhDT9RQcWyr4IFlkACWeKhAXXat/f8n
hdgyHOMGd8+2tjhfUXu1hItLgGOWk07YUCx97Y4IWy0VXa4JBY0wqBUL1ZXb
OoXdQegUBhsPgUfU6viOjJFF+dh1A3KAyMXhaagel2viOi6fhQBlrYpMLTQF
tMnrBQdqr1gBovJB1WOdbLNSlxx45r+AaCMEv9/XLbQivPjle81WPECBmBas
LP+pTdzNemKQokw5glT4XIEq72eqmK7Nw8NDz30jOOON/gtvOYcxNJtKQ9TO
i7Ks8nTMGIeNgyZW+w3TyNwV8860EzsrwmCGsE4gTozBGJFw0LYe801HfU4E
pfcsmm6HRFD/mCHVUKdLY+lAlr39hPGPevJEKF7o/rKJ743mCYOswNwmRIib
LSQQPEIfwr1Zy54IOlF3J0rQU1uF9ns0V85C6dZZBhYQMqzpDnY78ubFYFw+
RL4go/TeJIUITP6Oi7bwaQASegpobYp1jyn3toBhCmto+GNH+S3snI12yOmP
0kQbDgvKazNhAX5pz9AW6HwNIq/85WKYQ0LuIdfZYFrWE2o0yhr0db5aRy7r
G6Ge/A2c4QhGxRhU78FzqHpX5DLymwNjvkq1KrDkQ2S4LxAggFjDMKy7wZVJ
UsAvwBFdFJBdfF1RPkDl7iIHevp05UT+rY2En34sXy+MKmsNFRx+dO51QIMZ
P6j2/o50zbfToG2VBVmNRdySh3IbLOxuQGCMe21snA6Z2E96eESGrWZXNlTl
HBlOoUQ8QO+WKzV2r87Tzsjw6iSCJZaUTbopNlsb/Rj0VM4psTVkFb1slX7Z
n6Fs+WDpUVT0vdCCceGRQEP4Pkb5jtEv1QayYtgVjacBJ09eLkOTpnFFaMX8
IwvjB9Y0LR8iWiRATltQitqc/1gBUS6W702smdQ3GTttTYSReGXuNz5HAGG/
w6greyzc8MkBTZ9LTGxSLrmaeX4Dbh6U9YIFB6hiHMyqfjbM+nrgPIzXmH36
3IRXSF9iEWvJ+928ia24VuQEXW74kxsA9+sq1mdp51qgFqYzLaYtWi1nJuiO
YPaMsLeHHCPAOsoV20mAIxoCfclqKyCaQZB0qu9nhkFxiKte8yKJ+Q2ZUCZW
uNLl8HvfXRDqSErv1/CNTTXmHu75PaVysaEWidpE3Z3sdDDUSNxqgFgfeHRu
om3askVOP8F7QnUpYhkouRC6+5T2I3JXPI58zSjbXYANER+Hu2f12HuGdRrg
q36gIEbjnlJrkCUVMDMw6V16ws0isMwObHWqfR34gOpSKTferBBqGaVO6joO
n50hgoIBMK2fOMPW1G+58zTj7JKN5WcSjim33i+aTAsUnur8huWGAN2ldODO
GhXcrAMrmk7iRR8YXvZGfayYtUtyQa3Pl4HbhOfEpjm4+pV73xfabmwLYH+3
sO/sCSdWlPJPV0UJIK8sFBtq0DgWMb7bcPohbQ/f+/7uS3uARkFHzRI+Th72
9bHal72Nb0V4sLXPovmXFtgdKt+y0xhFAj+vOHqLFdIhi1ekQzE0reRswUCi
kU0mW8S2IP5uWK1eh/sNgJLNmq37YD1gdhAPST60xYQolXG6M/yPZd8d0Cpa
vjOkTt/Ix58+OPg8gMChfMUTR+T/cTckuVwdC0/3OiE3sE6MGqvRfMFv0Vp6
h5Ov52rEfIQExFKoEWSvAZIhlcEiiEdfqQ7lTc/m4REm3qIXlTLKVqUu1pvM
9fzWUkV4POB0xkC/5gQN0UCCv/YvM3MCSghunBiS56SRNh5Bxf9jNeKqeC4u
xGlfiJKcOr5AzHRL5aB86mgWkzD09ei7M6oufw08+sX0f0QQCGTNoYFyHRiH
yd03MJBVuTKWnfVC6mVIAE1pYVeHZa8C1yZ/NhbayLYazxgzunvWGFYqvz7o
qkWE8u+8kZnHfiswlpNhcUwvZkbNwqNLkt0wVlnJwd6rsy31TmSS3EqZEmji
ljfpD513t1KhJhwkVX2DNqun2mSprYR0ZdCznD5HEgoZxOhNFzWTdCkGjcrj
/TW0YnMBn1qASr8Ln13EkbScHvngZX5Xj071qHZj5AAfGi8PwFANZ3uan/aW
BYxE6jpmEuV3nVciiQfLo+xQXF/32XL0QRFvMODrsygbp0tSOo232t9cGw3o
v2RYp62JKun4Q4ZR1zoGl0LxaLExbz8/oGYcPlGs+zAjD14bS0A9AyJSVJn1
pf0tZntAPcl3qzvpkhy2a9/FRLZl4B1ygQY9VilKIk7DmLaeYaW3vXQ2Ze39
nN14CDgLrz6ZyV8EaKZSFHk++Ncb7dFsHRkeX6kIynloXX5tc0LF4P83yEDI
ZFVA1w3DatRlwwA8E9IP3qye7g2RK4NXYy/ZAZQpg1kLB5d9GkEZhMupnCZQ
de4Drz9SJbRN021XFCqiChdWGfbNjJ3fFIwZCZ7CvQdH0OWXfHM8jrREscAv
pYd8pcs5PBn53P989t7xFAzuYNNLsyjddcEK9b5JLQawGzBOFQ0dmSjwjC4c
e2C3c3DxFuOC4cuvZvz8r6YPKmz0FkOwnQQ6T4xGKu9CzSBhunwkcZEYRds/
+MwJgp/m5A53phE+15kRhFOJDEF6OSvz7+CjK63lLnfy1UgeIFm0rkRxkYWb
qfIpJDe0GNgMffkovnTwqcYyDFnU6vbApo3omzIyOT7k0G1qYMgOefn9fL2p
yOxUps/bbQMuOEmn3dToN6GSSW3IwvVvjxx11gpLKJ3SmOhTwIpmy8q4LeDn
qTJISnxXtQngUu0eYZo3015oOnJR7+jiG44uZzVTKJX9OOnRV8OM7mepiZKt
LlriwcEgCYzvQMAm/JIT5pnEzGfBJtgg7DXMYP/IsLgWOfIJ9nLmt+ejuxny
iESpJLVGYoi+w9P3QbHoWvoPu0v2dwng+wSjZgThZLhyA4Q2aCQfl5ZMRC0V
agJ20FTJQkbiHMfnxp9H3nG0Abxu21KvDmSc+GJLkLPLvHv21oKAznei1Sz+
53VvN8/Ncr/0Nxg185OaGYaroZQt4UHy0+vNUvHucm7QJVO6lV7+WGmNgshN
LsaYqw3sugNmLMroV/W0aoWMGUl0SgW6vJ4+s/7Qn1k8DTpz7du+Y3KVTkjf
0Zyu2pfB5RpeOn/GUZEitg2DKxMvhaAw54EZLqNPA42eb30fTA8tn+vFpi1S
fg8vHduf1l5S3WorrYNq6aF4bP4hFm4MWIJ52czDXHYhxiJIji4rZ1H9fy5c
+99HfJfmURt09C6p4EdKMer3Kin7EHDI2KeWiI7PStpW2bcDRfWTPcoVeJAy
lnXwHm0SrhFlMmpaTb7u8uouQ5jNmkLCNoyoIQ131FlAG9UAF+vWFQB0HMCL
2ETQcfX8TE7NMdJ1fdGEcf9LNA/DXic1q1+wZR5uNvxosDdGHIbNufxlCNc4
grcma1EOUI4uNcXExlWeGPfBXjlCDRnAm/W14ZZvEjahr23oQIc1te7oYwiW
39Vyb21GIPZTJUpsArbphVHlKlDEnlzR/6XDdFiMzgiRnXtCLUngQGF1mS3x
+aRgBNcZ/R4v7g3EjSfBaMFEDkTmFvo4a6zEj4zF5EGEFBvcvWtHpAIBDvfM
yCaK0PbY+pfe0Bk6DNxhFMucMeZaqKT3oDLCiHvtTkgxvDRdFQ4RBylPps9m
299a6kPEE29g2UxnKwHBajf2Yc5DjjWPhrZ3QBOrQmI7++5pYJ3xuaasBEoN
GHze1Wu2AhpDcYSo2IR4G3WjIDvPIo4HjSL+TqxiyV1lT3EKGyrRAv/uWiud
m/YnUQxfpx9jnZfi6QLZJ0gBR9z7mb6XCKFUuvFvV1sRyYfl0IzXMVUDvuzi
q0222LzHlt6BZcxOtvHrhH0xllD4xy07eW4aKnrkIHsvGXID5GxCqoXHRTDJ
ge1rbm82BrQju1iWZeUysVuTvdU5s72Zq7qauIWd5UVkiep/HRQgDaniVt65
E9AZeA+1CnFQ8Nur4zIH/0kM9Th3Mi+FEqqIK6vUr37Gzk5O6qhCvgKsJNh/
JSfVjWHjhbohSbBsc7sbt91ZHF7m06WIPIl7b7qJaXAstMwyYnBlRHLss90j
YiEJs77BfXuApHBGlElQjxUpvNPCzWnG56n3JRddwwb9pn+IzbXvSb9gxMu0
wpArQnDwkktPQWtz+IJQSq9t61AcoQq7zOE1gqEbWqA4cReyZtyxhzoRy9++
Rl1blCEKj8S++VZjImsW/OB5Ffg7eR4K0/VAxEDaUdkVr8TUYof7A1bBp+R2
7jngDTklaO44tjAdnNh8Y28jdB3SOoCxa5zSUuHv8YIT7ot0tuMUU8a2Qzw4
u4nFdVjOwhagu3Li+7Y0lxxJMqzPExgwsi1EnH+DdWdfgqspVQa4M+WsT1t8
QssOWre6ooikoZz1NLQWh9+KvWL1yKQICgohuMAMzKf2ctXUmCYOVjxOlSd/
Isj0zgzt/i/Nh18POHXpWahiTTFoveW8DTEVXiARvaEugu5UVFuDiJ4ruGP2
9qKii5QiSpeHSomUhXKZz0tbRrW3S4AfTZCZGczAPgkHNRVFPcTrW4l3zR0J
yViEqqdB1wynSA8BD0AaZWmg2T0bQ4NqOshkOpzmlEsr5mqOpEeM6ph24LPq
OO6Rl3zVcdPJDDqarX5up0qB9Epx46bdOg6zzvrzUHSyqroRuSLq1glHf2cz
BsGPh55qjOZN/H70JzqKAlYQc6JozZPw5JUEufmGLV8Ju6lpMgd3pNjAdb83
Fd6tbKa4amMTjATzpvoQmMF6l4MSNNpRiM6L2NXOzMZmq+cN3jC/I55wgRNf
Ydn09C41Cxj9NUtRnLv78RuJ1/VgF0sfmPF439pmSRAy31GdK/GeXRmCq0ZM
eEQzQt+xKogwtkTTLorcelsO7mkkEx6nYyd+5mDu6jkZ44ibrlZPpbaPDZkW
G8GSnoMCncp/KRUTjMHeHP+FIanygXZ07H1iTBN+c2EgIaxVN0z1otOak4eJ
cnFy04F9kn607b7EWtqDb98ef13Pdblp+Nat+EwY27KG7zix0pyIE0Lt6Rax
ZuYAdMG1eFyEpl1ihjnfNTVKjbrRMaJq9Gevi4PUiAnNIUGzog0XrXu8Mwut
W/mWZXDdyhYZT2dQVuevnlAI/xl6iC3yOK1iNxhcKFwKxC29+f8lAtwyivjg
0e+9ISoIpg6THdH22CJvqdq7C2x6H7Z9AM8J6+h9T6nHItBK4fBUcldyE6zJ
i+VGAN3bOenHkgez1HQlSeSk6oJJGY+u87uScCkcnIU+WmgOcbDu4RUiNHVn
xgcmcFF29Eld3I5OLyVk9hcugxZ/w6ZpYyOmIHs/Dg/WyDxyBDBikTWejvgm
GaFV5fv1B1VxRs4L4uyd4iiwedOLS+f+XzwlR/DeVmHewbQpBbKhGytx2wNx
jjJCToOU+vktNt/PPc+qY5A1eVZjk1DCKVD87X5cI79BT72IbZtGGeGNdPUw
qiwdD5r8SzfLEZ9L3r6Zss0V2Wv/ZQx/kdVNyTLQ0qTLD067P64ClCEu7xlE
dbI8odSsrm2Ony6roqnmP1We7T+o/FwvB7dFpKLlhUttkuCAdWGJ0dqJ88S/
7qiX4FCxbvmjM8xEaCn6ZrpI8hCl3gRMq2OKO7cxojTt9UeT9q4CQc8O0bsL
lkYAEkyp0hBDtbtpZnAb0TVtTizivBM2DClriDwGKsbNZb6iAzRY1fMptKu2
6gvcCvs4OCN0caQUMRiNmDYWkG83trRsH2jmAogR3nFZnFGVTbyHFwpeOEPt
869Wt7b/ZsJ/Fo+r/AgIYBtwECOR42G8/HCEbHZ8tbIzgNbVl1Zf0+SiFOsd
SREVXNphqC8S3SdyD9kSpdVYXBcgUkCot1PMeXyoLQty1sezchjssmtoz9ej
GVA8tqGrqmDiMVHjkEHZr5VgqseMcP0XcfFdHvlVJ4pfT7Wnh6El+4Am+P9m
RpKPJQnNW7Xu0MPdwh4P8fB7gXgW31R33yJByMQ8SnfgC9q1ZWPvf8VotHhG
b96GUYxz22+7JVOT2ROPnJQaeodKsWC/LEzkkiOTcFckAs0TzgEL33vrUXrM
k01aRKo78MoqWwAlHWMwwl+GwOonM/puKzLwBVZYSiNP/gPmjWq15fPgmAIk
Eqiaq96uqMM+yBsC8n/FgglZryeLuaH+SZuWo6kCbsT2cPEmd8IUrRTi/G1X
UkLHEIxZjp9/S6oXYcmasa0YN5L9+g0+nF+xoLQmlfkITzzmpkiK+uboxz3E
28ZlmJa1dBaX4/9Bz5+0ngfqpAI4yAKuMC/cs0q3RisNQ84+HqkXRIVpi49a
lUAPbVUOSDrLL6uvxSjINWcl8tP0YQJbN8G/utZwhYEoLlQ+cnS8dl8d8DVL
AV1+XvHJeXFluy+kvNgMJ3vVjLFnuB13ycU2xASNA97H79TZV4no+/moRRX1
MzeScWT9W4zzE5xHgHKYYDZpPWNTUDs+nodgBPj5eyWoTePot6xaMZk9jn8G
+1/xpK+lgEKzFnf1uZdAW83ahC78spHRrua6vqrHrCwJdXm0aOrSJO/a/Ieh
Psfh5+pEg10UG3B8ZStOP0rTyOJ8FkpyLELIj1xUPMGqHka+KI7E7hfNDhmq
TRBalj2ukwmU7JrHtf/r4XXnsY3IIEnI3OlOilU0S6iv/pXI5amP5AD2Nz8E
3/e4d3Kf+yf7t3ClNk6xuNJuRpb2HaVtkfwNNoLT2R15edZy/MgrV58NdYvg
iQtV7unJujDxJfEGMn7sGMu1Z4goimNshLmkgfZh1iZhetlAthfptQPshVs2
FdCZmv+Mo+5SW9GmcOcQEbgGuOFkZlPBbwq1KJLI775H6WWMr2fjilXO/Ipl
xlr7K1xM9H9n+36+RWFmD5LG4xnZ+K5DjYlYy6pQ/OnImiMEPDOU3VZXIwNv
jPILa4n+XWLjSe/buClWxYGHeGXj6BwVWlA+dXLcIuvFqk5g2WF32S7N1BZV
jYjfCd62KcuLwwYYUVemR6C9hV9tSKhgUh0Lh1Ty6MFbTrqYxGWnMz64/EGB
p9FSDvi4Ky3aIhx3BaTU3lFn9XbzlFL6fnh+cG4EGuaQ16VMuyzYVSXyE1G0
kTull9JA/IVbDLvzS6ZaLkOxu333gdV55/SC38W8FZDo0FklfBqWLInI3GCa
63Z/JL17Pmw2r/k0vlP9RkkRljlOzhfKtDFbjvjZuUfSGQpi+mvgQQD5nPM9
cTzk2L+oXBt9t2ZLWQUE/ZugrNMHoKQvBMihxnpXOyCDMOAokmLgiScE1+Xr
Aqqgcq1nH4ued3Jkq9oSUQkcZbflvrLY5rmahh8tcQHEhOEuYOYsTPi0nhcl
HE4Dl9C2nHJff2I3oNun5J0KDr+NBqEpoMSwmB2Vqy37qL5h6M6TqmL4FAw4
b9xlve0Ba2LUmPGBZsxdvAPCGSLD28zixmapmtUgonn0J/V5bTw1DoPd+EnJ
25Qt44XJP0ExgZ+gWSGC9WHmy3G/XqKDkUbvQ71Ir9bKSM1tZAz7ntPFV5lh
UiFE2iQDKgHh4wfV6gpHK8BcibZHKNzzedvPE7wZ5/PPbNoic6WA7iUhXpVE
rA9OQVpNt1LZ/t4GZnuTRaLAGzvKYai3Ukdz632T6w7/b1W++rs10oM7TfSm
SpiFSnt/sFZKUxt2e0skC3eJOyUsYW8MDd6ZQXUW2gwfcw32ePYLzoQI/VhV
rFwcGOEvZhS9PE+7xlen7TL8jXwYoA3DB6OxB+2cZMS7AiO0b50WO/fYorER
0++KmYsSgoR3w959OFCT8SZow+e3GL55399Fq8cpxYLRLML34MR7VnQRBBGF
zAgmMHWAVT6SCE5lbErnBbms3tuKhHlKE9d35HfjOQz81avr1GSIDVJ2ndmu
RQ65/kTVoJz3nIUlpO6u4o98Zo1e4+B2kWPIfeZdaTi1KCdNcIRDSgTelyUw
JX6rtP9uhR/mRgStyJEOtfGzVt33XZ4KCCjLRb480g02sAC4WyrN5PQ/ghnm
MkW3crQrjQTFomCmJRLk8fN67R97R8iIwlihn9gJcWTGxXWTZStmmilef1BS
iM73Sj0veweCKDBnytWJ0xrU0iKTAtqxQqsc/KK6W0EH0al3Jll1jCoT86AD
+qtzRHtIEdZI0V0Ga4qG+A623inpiffkO5xXAtu6xKh94w77TK0pupWVUOiI
GuYHcOa30ga9a0b0uljU/H3v6SkRm6hDDO5aEaWy7XrcByOHohrIDQ+Knl84
7/Ixta0OM9WHMwmeIQRCnqBic7b4Px3RSNoOIqE5G4RuykiWb0P794XgOOOv
zkt5drHOQzSRfl8zLUjRt5JiiX6tA6ain50ScjTRiZvK1R6FleM1siA0Np07
RmhyloUQHHt8ouIJnrkDaPwLYiloSu48GeTA0uEk7WKHSTLMQlI/fJDaHbJA
HLW3C951e7/wd2t6YmH1mGvGsVrY7/beHcB80pYiS44uI7C7DTgri1WBZq2X
kG3Mg6Z98F3IniT/4rDrNsXlZSjrV9m+2SsWm7ppGoAGUhUvscCgP/tcD9xM
p96J06FVfQZgn5cmdThbzzgA/RQ1XIoj3XKIDy5aoDI9sm53aKVaRy93c1v+
Ck+51ciKVKF5Jq6MfuWJoaO2FwxPwvogOHNwJes2Jq/Bwfgo+gIGzuCmksd2
mgb5BdRC7kpXk5mBbsHfLhCYQnE+pzmGAUrFyA64GD21mw5r4cACa2B4L+sZ
Ieq7zJjg/t2B1F6YzucjZpISzMPkrDnUgTBlG5HBWHGBrKo1jk0rJWj/XevH
BREvVfAt7xxOJuO9rTsbWH54guqK2EWpdz/w4xPF59IrzgG7omD6YwfIzFSn
yeLH3BGYNu4TxsKhAVE5L4wAuekDQlL2yHxBQKIXip2Qb+vYBiMXY8IJMRat
h8EAAQfIZczldBn9VABCzz65UVqXNckRB0Jau/RPNYZI41VwROH4kMG5j7Ip
WybRNwYnvFEJwIGV3gS2fzCCamHC4Lb+AhfwVRFCdt93vmU6+RDKJlyCLTRi
UU0cI+Hfny5P6ZV/J32UemR2Ghi677qw2Tad1QYW5VEzi/oN/IA8qjzxjDQ5
wdb72P125PeggNgqc8o0QaRk1FOyoncGlJmgUJHSO6QDabqdECIoGHk42TbW
CFUo9bhz4SPoYscsxxoQD4bOT9J2Yad2VHKrCbvhDcB2Yy7GaMcmLcfAXlbR
iPB3ZHuBF+jvQMg1HCwBfgyOT6h2vXiC0/ctua3TS3VtX4+uAlHHjFhGlM/c
SxLrgp/BKC/C077DuTp5jDtQEgiIaoCnklPC9DrdkLmSBxtmSbItMUfXDpfb
HeuOHhIOsxd0mCZHx3rHaZDQOlMj1jsKpiqlmfBWHsKUx9hyFpEiIOgt+WHB
PT4O8ZW2TD9g1ranQQSVULJcyN5OOCnL9hlvHHh6BKlalxhgw6iKnVkZpLhf
kR6deXlNVJECwdTI5L2lXOI6a1qP4OaDPZcDL8xutmZFd/+oIoOyNYEFoMox
oTcXg3I2khveJm9NvAV+ZixA7gPcAzkH+DIMVnL+xd97Fhao2h6P3h0IHe35
pgRA1d9Zhb1ndzaWUWpgjPimMY8IMFatNbo49tCNC5Vov0ku22FaF/NZti0y
GyscYsOniYJbyVz/YBI9pZUciuYdsS/Rnnzor3ry4f3WpJWhvdFxevHhyC9O
bJj2QmeCDYEEbfTyGSYF1Y4BEfWAp9qD0ZVUYwHLiOMw9whCrP+a3KF15hWx
UEuppt8vx3jYndZ30F6D1h4iwSCU0YUNSZCCGmTMglZL+yJb4nC/GoPRNDQR
jFMDGxuF22mio6vS6x5Wo5NQ+SgoBUMdBiml8e3T7N1tt8hRZSLTyANa9p5Z
qBRcM1UifOzKz7FPqhkfydzYlmgh0pLJOmsUjEvIVz9629MNYr/yNwj8tdaj
6Cm29lvkzOxS+AXe2xGhuKbwSizIvpvu9p4yV5npRcEIg77xbEr5H/ALI9IL
jJSeqF6ow86vTQRb55PIWlEilB/kz/uQym6xanj7KamWdvZHpWYmdgigE41d
t1/7h0xVPKnATCchxWQ5MJ4VM2Lmyx5Gwnh9GdWobcamafR3HvkwD4zrn53B
MVJN31OcjPnv+qzlD/jzp6XUKxhWKzag4991iwHykQMkQh1A3bGfKXR0zagd
mIdbwBeWajVu+Ar/y7Z+oduDKSqZlB/jyKrsRCSCD29QHwlqnEuYmd032yS8
OLXdkMtRd5fpRi27LVwjXKOXqQC5yRt/zQUEO6eXWzer9B8SybC2/tbyAnJt
QvRtA14XIPjEkITAaZT4/+jd1Amti3/TXIY8haus065Txj6yLr3LhhkRyYYX
+CNWrINHwH2oM5602hIqjw8iUfOTBCrJ4a9N1Lf1i9v4iS7tIHaW8rjfd/nW
FvWBzQgsbUpm2mkStRjz2d76ZiucuLnBaPsJDrWElhRtubY7dC5J9WFHUNdp
Bt89fyIRoXw+v8YLi19b+DjTWWgbl/Hvbwz+B0QIoNpHnBuVMnKfOeCNuZof
tfuAgtX/1hvJrKcu4JNQBz7nD2FccwWvLWk0E2h+VsXcDQYQYYXvts7Rf3ZE
hGFIYO1rBI4iKx8C5H4qRXh+Q0ZuUnDjuShUbqRGT26dMZdw2oGPqi+Mc/C2
07gmkcA++vN8e+6Wrl3p364gRCmawcRCxpd8NR7fxpvnUJGp3HDmk4Aaag1R
aAiUWfUL1zywuLGA0azvwkGGx1dF1gdN+eH0hC9MuqPZOgDOfYD9/7Yd+a8p
WGxPz/sgzJwH+yin60NS/Dsbbc9GhSCqQEgeRWHiuN2g3RZ1tr7ZIacrrIit
ilWFn/TKNHSu84IMz2lflYnpczoaIXSDWP5POeahbG0s1FYjg9fGb6zung/g
6op4fwuzGzwX+YtWypQ4dhheSgFaIjRZcjgi9O0Ue4GqHh5pVbDU1zfaDafh
V8aEvD+oaUirdmxcoYL/twbpKbMDEAZpw0rIHL/sBqedjekECWqvkxWvIAAo
9bQBbBUNIvnC0KAR8fUJRNscD9BZ3dwtyFfdnIU7Xyf7O/ssIjezF0HqQpw6
JjBYnI/eabmvLlT1dSf5bn/fhM9mtIGWlFCwnKGFXeIhthdyBEiiRNz9u7JN
GVNsVvHcG0yyffoyCOH9R1SiJmgcLtRqVXw/N29N0C+dyc8arCDO+GPiiv0O
haz5S2c22P/rD9QNRoZ6vbVkK1VcxIt1Rj3H9PtgBQxi1mgGJ1537ona0gLI
TI8/qwj9DJ5bQFE8x/4TjUyExAlyqmJVnk9dSgEC+L97MCBWKDl9oarad/B7
dk6daJeNx+4jiSVC//02n7aZNsu7H/6vOFkJCnCtXTBe8Vs6UDQnVo2QWRE3
eiTcMeZ8MFXyORa4321AlYS3jc1xBJjPP/uq+sJrzXOn7CcLcSMRk/NYQbOv
/Q//ykR/RfwJ34NNLPiBOpTVOo3KL/h0h6i0+/x6p18iSP0tSwOXmt+80Ajt
7qgCj0AVhIDcX33Whlud1d3AaNDYhwhEUKG34+ngGnCl9izZQ2WUKakySdS7
TPhUdkJT3/GepZZRPWZOpR9r8LkCGJBEcbLMZ4yHBnLDyr7ZOLFdNwJzbONJ
yyJQ4lXdCNMsRbfiQgxOf2L+3OqFFvYsKghunRxcDgZELLHKsW9QhsRM0nap
FdYXgSFk+3LKfNtUJZxtkVzeSnpYHTakNuRZ/AiN/BWsWrsvAca/58zybAlY
0/CqJoXnI2T/2/k/cqYIlRWbWSYHd5nePV9HwG+zqrtsnuFjS3d+/6EFOXk0
Ctkbtupo/K6cviDpfXRmCQAk4VwX/GnnCgK+O/1hZNwvdmmuHjXi+Vtp83cn
yxibLtMic6gRLf5HeRMFsixEtH8YYaEVhS86dhFhukHNv5/Z+uoN/4Pc/oyO
0HWohjUtN+6KYBbeZVTgtMhtGe+d3oNqC0xUTU/6NcKekt+dTgG7UA11zEhl
4HuEepVo55R6myGuXFf7w1EaQsFNi4OmoTAgOSbXMZGt6fEja4/od5LJbprg
owf6WowXSx2eGtEPvcgTvYoxFIRpsrZKz5OhcFm+BbEhStDfoZnGSo6M7qUi
Qz/NjhedxLTJAc6AbY0i7aSJt0Hih8Neh4ICnG1Ee3T0g28pazh4+Qbk1yXh
cUjdJ2lfelaDVdlABI8DQ6PuHJ8BbDqM6jFiHeCoGyhkFIS9DpbDTA6lKO/+
nYB7vnPuq9zw+gDhx4A84ZYoEr9+pcalH2rJYuEGAzOfzpZunpyFhXeX1rF+
5NA2PeW/viDWTmnqM8yOcMe7g8S6R1UqxSOsaT9ISDauVIpoSH1dEobJ60sO
8zkQx4sHcCaS7/goTQITyeQLLf7XOW2Fm71tBmABjG1R5R6coF2VouS2loFr
7Ymt0a10tCVyd5nVHclNT9HAvDOirp9p1KPitobBzG7xbzUkORKPG4yBQx/L
XbQgmg3dPwSz9K4dxiw/457ghZwKrX6JvapyCv+dpzWd+1FGe+z+3hr3cYBP
Jan5WaVvdokme23vz8oio+3ciNMt/pJGmxmlgsIPQzc47tTH5sUb1LlfHvAG
uYvlTt/qN093Ng2H9zgOr5bPu8FV+BXPozmoe/tAbJK27I/mldpPbaXDVgK2
v3UDhpo1JHg8LhJN1DnxILwlfX+sMe+4UtrckQOBG7esxpxwjXnZudINMGXU
DYRsg4mqo1G0z6nzzqzC+OH1pL5MwCHyu8OwSOgZu5XWcN6zZEsyNd0Xo34Q
5JzE7r6SykastYl5CDdULVHCJbn6rnD8Y7NSzjdMLvNiF+Zk8BWyyFBD1HwO
aFf5rTnSp3DIVGsEcIuPN2Utm+KNAjnUbxdSEISdn9wtCXpliu6Y72f8oAjt
m7TcU63abjwkzTfP2IAY5kINqJqz7crIzZtrEadrntNLf1dwDrL5ar7EBjd9
iE+oDqjX5VqqRAwJ83tJytX1B/1fMriSI0slMpaIvWMdboxG5rG4+pT28Gri
X3FE58y+/Cr6zhj+0uHg6aXmPMhZ55fMaq/CuJwUvXPcpPIyGlckfdR8Uouv
kR2lNCLLh3/QZVqm8TtDbQgsatN7qJCzvrpqCikO0cC80IcFMwvE/vEEQ89j
C2o/sDNa7v+RmTuq7tTTJjsZi4JIwJdDOOEKPzHA8a1a/G80ZQRYG96tm8Ez
h2++gsITHOZVlAcaGd2m/LDqDxdd+AAMKK4JATtP5sjv38kyd++WfirrFFjQ
eV845Hg26/z7JbaWA4n7ZHbjqw6pk4Py9ZNa8Aq/+wZdf5ISneg1N1J4K/NP
sMDAB91lWlxa5wSkzmmKn3ViYmprk8MNRbu2tkF4KgODnxHSmPZ/EYBwcbxM
Da5Pi2kTW24fun4Vc0Cx3Kzdj54I/CBLTVZzLJ9BQjU4qAL/d1qQULCSJESj
6PLTT0wOLpuIGGDRPmMGkdBpy1nY825exOTkNCy6wT+pgAJIywMxVtHsU8ot
wjjY512tMw3VrfWBcCW0PJnokGPxrJnBjXVTUBR/fOhEC8FAC5iSMgGqmKMg
gdU9X39KDyYii9RnyMjyu5A/TFHqEzw8nsuNlGTFX32p34LMoSnh7ESpMPye
xpQLeRk8tZuXabJ39fUW3HlbzJQQCmJw7EbjXL1F9SfNtZfy/C1AtvwnUvGS
8UXFMLq49hkoRDCPPmgq80cQTd5lYONY5i5OxwamodEoKB4PxOUcN/ipDDFo
1OgGniaSMl/hG4qIUVJnNo+29HxNdVCyisRKkOiKzPKmmofckGha/7SpSkEE
k0cmE6LLFEVo6wJn/Cm7JIuIQP2j8xGIskas3ls3B22iwELaPO4MBv5qwy97
DY8qb3R6XpI3rz/OOD82Cu4zHbLtLVKMfCQiWaRATiVSPHe5+liRDyrrepE8
vUZAs0Coks/T/oHAxowG4fnrZlWOvbk9cuVd4aE0WYZE0vXzXsqI0/Vq3ExR
HszzgthE+5m4ZCHiCsp6aht0DuEHmz1SxMyAflogpbRdImtiMMLASrg0qgwr
YGIXBkdvw8EPTDbGj/yNvxspauPbfAOYloNZ2h+c54zBdK/F2aM5kuo7YaLX
DrWIkPOjyJiadCQLI2GfXQCtE6g6da07Tq8GeyIeAjjFXcp4X16F3MKSqFfm
cb/nAho5oaOR+VkX3f0HKURu/NffQyweMFEqijCkg7OgRKouFkM+gSwAq4tf
q55RHHA7LF13nH7k4KIRpqeR6mjl7zkafAbvhPmPuLXiZ+OKgx3lywLycMTj
1s68FKqSMQttJCmNGl0YfOswoIpxiSfZa0FzUpOcSYI/6LzUdqh805l6Bbn3
Di0xzs2Ft5R8ZLux2ELjYU0J1bsvpZJ/XmQWp/HzW78jdBXNew2O3jwctu3j
c/xYDU38jD0MvAdfL8fJO7bj5/2+xdIeMPjlROWhhMehEiMJw+oLSaU67Gm+
pXHAO/oC02GzUqGcSeC1JTVwtO2pgsC3RFgIaxhXdezJz/qPeXsnrmh/pMOl
JcKVpveBb0pTY+WL0RwzoQaBfQI65htOMJ2nQfKM+Cc5gAMKyVPiJMv27sex
SaLFyRUovoL/k932JFhlNeFSx0dHJ0DscRByjdU4igWUg0Whmi8E2dMqhicb
3klf8JbLg4eM6s2E0Bie2YgzYBqLnolDR9PhAL0kxtCHgvnd4ZwPl5VsE8q/
qaXvF0ySTJgKilmT+nkLaXvkJp1EE66KO8Ys8ywybPK/wFnMQV4PIS0uOCyl
VBq64vUHCHvWz7MfbOt/EhleoX46MNt7l3ntEkDXm4YYx0iNF/NlHOBGHhMw
pjRBgIRJBZYIEtOBPZ8nliJS3LhEVMl6zp90Jy6lbEOUzX4LsVQflnXSUujt
v92BxvHTb9VkPdhYjQSsKxpb1RwS4lDNsKe3qB8EPzVHJWOu2a+GkISzn3BB
6h7JmNG0BGDKTM2gZnCSCrO5ZSpf4XxfVhg0+yxXwccT4a1FoIC0mfwPcnIL
UmowRWDUaDG952nkVehPWUjet1zGHjvYTSYzBbheFOMEe92lUCUDjeJxG8A+
RaknzXf0zDFVZppWk6rjAKFMj8TebHkFs6KHGTItjsuBZl30Kq+URM2K4M05
0OqZAJCg6Y+jWR3+uODWiVOxDBOE/9h08nlTwsy5CgMa5OfRyXTOqKE3Xrip
Uo7neiX6rMGsMPiY3ngNh7L4LLcVZCuMMiu1Mq1OMOUqJcuFa/UAciq1u9CI
9m7zOyyTi0W3Fi/xK7BIBuySzDpGse+8cwLg8/yN1/xEs6W6Qx3ErQfYq9d2
Ia83A1oT7Dhjia/S5WhTnKrsbT49r3s5E5L0Tc6rxAF/Ig8+L0pTOG7v5sAd
pmV2GJ4tBTIcr99DyF/DxSdisu+DDToUCFAzxlUSO5U4E04oMCfGsmrPRLmT
Z4BBBD/MNnXmcgz4ldna1KzonRP7rjIfFCJnz87CMael1GhGt+A+LTIPn6UK
vYe068ijVTQA7q6chVpCdk4EuQQIitB31weuEtnyum16XfBfa3P/HGIL0iHE
ipMBFl8wzV0K7v2/AXCl4oU9NdskQBYrB4qqEXZ7ncOAwH+PH/BF8BRebz62
VAYkR+nd+Wfes/ismKt8yY0yUGiWtQjYPrk927/l+ko75laHaxwuEOWLP83P
8h87l6JYOSXOr6cnECVzn8OrbMCkUdHZ1bizoH4QNNVB4LZZEC4Jb5hCoetg
rp3zIkGGMB38o6V/zeCFmFcPWMT+SCcaVWNMlG5SpviDBfiXcSvoH18vxGqA
zlVlVTXgPYVnPm59ujzYq7vNdoCyCEM01Ps5gIJiZbMF8Hidk44iZSj6T317
1q491ehMgMNc5QgdzFKmscemDsS/QfLTi4k5taK5HpZu1gG5giufrTeR/7wQ
l4RxLEU408F+yiPaZ70BVBvz1lK3ZTifJvuKPX5h6zStdW6aJwmNOwFZUqqT
w7LCqRwgedmXf4SA3Ho1Sr5ax/zvzQ8R0yenemovypj33YKnTalnUsw1xVUI
dVBqDDi1byLdzFPNIzPjg+22PHaOkkkKLKREK8P8YTACye1b6wFmCVqavFgh
EQXF7r7+mJfDLSoIAofSqYBTT/dPQyU4IE2c9dR6oKtST57pvHj6WV9olV6n
AlCf4lpo/EGQRSa975K7uXMuCkpwjUFgZ/NswjJ2QsD1Lg7U+F61tDgYujqC
3U16vogqGxmc5AbF6/MrohTYEbVt8m3KtMuwBRankDY5n0SqwvKxwOmKKSYf
yvRZit/QUS4VoyicZPi9qgNNd6Z/uuAsC5q7Az/FlVop5GlDTAjLQIm67ZDP
JahRYJ4wDDiHl8XGyvxLPjz8WSuCB6eXs/HIQEcVVr4iYDpIa919JFZtNZiL
q+HwXumDNZx6EalKdqGRkC65d5aqOn/ZQSltTP8aYLc70tcMWC7yl0iFzrV+
FkSJsoeszro20/xUAC1Z40AXmz/Lx1Ou1XCPQqVeFfrsas28fwjcUSzRdy/O
f9ih36dRQ9aXyE6Ic441lS55YPjoZaWlAjJ0NbtItKEK6zfUfc9EwsxJojIm
bmUZqdVf7KDBe6Xg7HFFnURUoI31AivcZFfmiKNrjTeQaOi73SEyldAcem/a
r/6noReqKFulp0SJ3gACIn2H1n39C8BBXQcvYeSDL2PKto85J2Xpm2BfETKK
n64ujP6vIJMQ6E7YKyrnx9qofv8VydyhNL9Q+gcCshUOd5xIVrAoP25n/gGW
PuiRPJicC9QNovqxmjxCuZS1q/Nw7gu9nrvwwSNTHB306VKnL5xSWfmXCgC/
NFPGwI+rXKfwAKtI4TTxzf3/NaJXQq5FRTDn7jw8ldzGplok7LMadMRik6ZZ
DEq4B8pn0x+Ni/slvaUfrhk2b0Le1W9khwaFvNMyLgVUoCA9PZV/PYMS3H9Y
WA0BolyZ9cdwLVQvP8gIzidco8A32YTQwDAkOiSUZxEIY+Lvi+gH+I7ON1a+
ai2XaP7ldYjrtXqmS3KnI8Vpfd/jPMULJTdHiAYrURfLiNEoiysslP8z95pc
J9uUkrMN9Fh16JqLE1Fxpgh8myf16gGz61WdSEzcnWTfBXqqmuHyRxF7kBio
deuu74Tx1KA6nfbx50gz7bLRg5J6hiVT8Uh7bN3hz0FyKl5kufO1eFGKcsUx
GAys211g6EN8HtWCilR+Ak4i6bD5BuScLVcVk6BQ2YA7OnDFRMsUOyn4rrJJ
GywTP6vMfRAMvHRWJj1fuskFiueJiMPba05AtB6weMnfKFvETJOYKs6+wgQn
Iwo8GfpXcu1TatRLuH6mo7QGIJ9VtG6OQMzgbv1KVKMW7hD45X3eoKJAmC4v
L4AJ0dTAXovVEmS9fKjYxk0ajl4e/grQ2J98YsiYgP6FG69rrNWyrsjKi9ug
cpcDltM79elIA3p3+xaDD46O8xo1ttMX1jDlBjmzTo1HQXmL2d5pR5NXLtMw
tBHit7/7gfiPAqtfZM43KcRg0IA1HGzug/gEEG9UMlNIoC1hSPbduerwWWbx
PtCmYio8rBgreLZGou056yb1gK6bdNG8Vpq1XwdLf3sd2gaReW7R2blufhWl
gpjxVnVrEFnTQZSI/cWJ3h7RYqKvbUgVxSOCM0r0npnvmOGDMvYV1FKp6vFe
UwJwisLDd5jfCE/93qirtgczfh3GP7M82HdKb4cZxvQdE7v4tZ6BH2NMnS5j
I72wlwjNFGp1qSKEd/bIPg0tKvowMfbceXtv9InLnnNZ4Sh26oLlwEb36s01
jYgnufKOOLX50m1eK4d3hAy2Fu2Tmm14K/UdlnASCmYpWrSZbESxwc/Q6n49
Hy2N473FucdLwtVdZHwdgpq8KFxnCAMNbd1WrMrAsaYc9Z5QZ1CJ1Z9E+U4r
sXTfb1Q+eh3DCGB6mXD1npCf+QBKgnPnCKaa+b600SpNQGHmjwezn9fNBP/x
Py/EyDsfxZTPAy2uMPcN8kx+spsdMa87ZtU9liQW8VgqAwk48c05e3uzygN4
EEw/ukiZwSRKZnQazqFPdCyf4hsMN/vCuhvatYp93IYEeudLZE9X8+EXNsgN
e0tmVnJ/Z7tbSRS1+UG2Z48Orzss8tL6h70o8Dy7rnnUysUD8Q3lLynzt94/
nVECre+kCVc3l7528FWC8+HQ6WgTdqsQhsqtw/jo8BRpy6vU3Di87vn/hAxO
nhnCS537b3wAfzRPCiwaLyju+gXWnI3OQwxf0jRgN9kBuXvwa1nzI6quJvTE
elIeRCVdeGjSZwTscW/MuJY7xmzh8TePn4pv6Z0KJYaI5QdyOHIjWWc+VMAk
vzxG3s4Hn0cxbjQrTHNz87Tm1fg0UMqVD0P1To0HNf7acF1Shg/7UFp/2jnK
Zn+2+yP0+Npu92R/DeJqni9i8Py0qIQF36Fwd5B2VAVluRJgGueIBdEL7X0R
Fb0BLZjPwEo6aqHHduWIYEhIrtT/3gCODNT2u21eE/g3T67x9DSD8PVM3lBp
Ko2ks44VOh0Mvgxvie1F9UMGXaviOfGj9TERA/JATM1ZvvcnFZvhCZAlIRl9
3Ii0YNQDJShQh3oB7R3vKl6coWNGkrrJb4RxTiEiHP/vqhwCkV9sBZBqxHdS
SxEj9Z7NX5vhAb3XB6rGPVs8qAXNch8e1Lrpr6ih6SNhm4rCfenyGtwcYDus
wTnaaeFkFZARnuqFAUXxGFLTpMJoqrEDqWrLvmVT79fC/f8ySi4xzGipsQRd
b2edrhbizb2KEEIgN5ptJI3hNMP5r57tmQ8zg9mEJfRMTIl577GBkOXe50lM
UWyHht2OBa3+824/83vOSJYBzgk496uPmFxZvtDYRxFDP8oGWcgiAjaHWIFP
LEJh3E0SoOXxQaO0o2a/lIwraxCJUnOIp6G3Py0lIgYO9rg5nZwF/ZarKu2Q
MyNLrfhtpyPobNEPQdlt4qOO0b4sJORI63XKe2RkZCxlpaXC1rZWXxoloAIz
sQrF3wpYbBh+ElhU5nt19BBOFwuB5dCfLvtEa3mBSiBquVHmZSB1Trfs81/R
ibc8VBBAJa+k0GcJMITFgNRqJSbZslJPmvvAmz5xBk4QXtRt8aBovK17r06d
gh/O53IaxBguOvw+i0lbX/3FMPF/xyJf1Bwm3DqY6UqdbMaI1rJUBY3V2Oki
s/fHK8Ih+c05m3ff7OUjH0kv+0XM0booGVRxwlkDTOaZ0lt+OKMzEUXVoCIf
sZGqbZNpfQQy7RHkVJzCzZi1eBtTi8oZgohyHWEjNgF95GN+iicfOO2bPgxu
BC6E2hjt7sYPH0UyESpYAxGv+GXCq/6T2cCVF68ORi2/tqeWgqp2sXgVGTRI
SexJKoKCGfe5Aw8DCNC2ctoklMlKp3DPMFksG+i6tfLzYD25cqH5oEKrlYSR
XRa5cxeTOE4p9u/IuKIxyLtv8hSd3xx6WOCtrvAg4jC+ZHCHCdefabXffyYS
xvhZ2XvfOoN7DG6Av0BDCqihf5EVTEMQxAYL8TpZ4DhpfR7UtU9fhXB2ze55
jOAAKZzESCmD5HJXlYIW3KaxKeEgWbQ6+b5SQoJfMaV/qafIPb0z3hGwM9j7
7WiyfnjEg25BRMcV680Iu2IM4ZgrfRkJRIBTmm0nHY5xAehmw0LodHwSQu+B
GaS6wrhQcjLK0dhnP9+Vtl65oid96zrVnTAURYH9W70+21Yx7M/mwYddhhfh
1/JiOVE2I2IkcSZeSIBX10buO84haFhjrQ8OSn7/wm/ER7tuQy+sp0G48a82
nY19G9nPgmPY6sjff6vmcaFkd4cuW1gnjpZwTvAw0U+MeLmm61tFJP174Msw
yiDon63o5pKNfb9S7Z8OAholva+ziCzsAFd2Vznp4d9/ruupvleHOtFk/o89
fsrZKjrAqDXazyZgYdEsjWlRTtGXlcVnIATWQKWHbfVgjROs0UaLmaivGgH7
A1TfFjOGty82e6pb2EzsUbWS81PHTlWFOEJq6LiKhHkq4jzPxsc17YjiIrGT
omlaypX4/sKwuTIqAN/A7JPyGMcc3q4FRGcQxmzLS2kAqclS1KkCM/kKI2CS
cSA+HFoI5ZroF6jkhbI+vlr6Rppov9pWwUr7e5MBBWHa5YMijCawd5bvtm4I
Hex9jXhIY7N2FSvkw4TRr8Rg3ZkN0t/2HS0maWR+IeUOFTX5kXNPvC/ByG6z
vn1JAHalui4qDzerPXt58sCcUTGF4CH3e1pM25V4igxn+QKjz7xpDcxPYI7/
blMwDbIrpElb9KAa2D/NqlEWRwXNZ+/gwveHhrRU/OXcne+o93kh5/+5B7IJ
hjRelhmEcAPxXxg9QdUlW4vITxv9ptnslYcGr4wrSfjKLLeleIa3SvBhD1o9
zlPNP7ZlFTF/6N0HxBMrK6j1QU0risv5ueMrRWmoJsegwDiS/EYpHYY4Fgik
XijwWPrJC53TQYzZWYetShP1T8Dz+R4UAWqAH6T8LVwjYPpciIoU0r6wj5Bc
tutZcNuWxaFaDfNtxt1pJmB+Zvil05mpEKKPTzJBA9djDx/HwfKJnzKrM5fm
2jyRLQn5uPoQQDS+BUy0/J21SiwbLopzRZxUFcjoELfftMR1TgkmsEY+9T5p
wntmgxgDoILc1CCfsRuTNtEZSpOmlm7kFpw3S4rcLh4oHPGTrDYrJOeH3eG5
oFyYGGO4o+jFumrHk+8b2PNFp87MNtwIhYFuLfUgwiXlA7aQloys5VJ++/7w
mD4h3KBsmzrMZEduaFkhY313nqjtUyhZASQEhHTB5jdhn9GK2QUH7KGjyp7C
4i4Rrvd1Y2fTwQhysm460fhjodxVHmW+CDGNPmk5oWSzHp1l1p7k8Etj/uAQ
87uaPeXLsKQNA1DwaD+yS2nFE0W7LT9ejOtSJopC9q+8XLY+h/kU4zLUH5Co
AIlaF+iB8LHIjoykCgk+LpMxGVTxipQfbH5gXToB9ALHVxinremHyvfahG+i
w9CXf99LDD6cIEFpdqNPdUGcnpfodG86KZ31e8o6ZG7LeH4o/Bq4SbXeut/0
57LeFheQJH16ljy3Hneo1+XksXz7V5g+kzVOQ/BACPrIh3RbZkFVHxDqej9a
HgAQtR/jfK5ekizLtbedRPmfWuINxqBBZncUvjgYP8DTFziChV6dvCteILdd
2eQXB5oKtz/aUgFRneJj59JbBlsLbPjVh4KafTCAn2tgIseCZIQmdA0c6slX
J5JaYm1cZY9+TpADnDEtnkaGMtaWFzKxYtu/IJtgQKN2wOweM21f0HXa1FgV
/yDwVkQT1LCJOOIXfgJFXD8LUb/9bInpuJokAyNuMx9mX5kpJqLnDXM0jK5h
1xhMJ9s7eWcunmCxyckkCQ5Xx73rUzBXVxfjQUQZrA+xs/V6nc4EPozoHPwu
yhJ5g03wHR3JZuTE+X/xnc5fE4wPdPuLm1wf/G0cpdUPmqCkFQYIdyaEQtPv
AMi3idFrKONfTxfzXZe8F6vGMtKs2AXzqXIbx+3LkRIHi1afNQFBesCiRwIY
rU6Ecz7wfDksTbu0BqMJ1jwmZuiCkeE/75VaWbV/8l1+syjmzqJmO3TyZ9Ws
B3nAhqVxZJnGZ88doy/UWC29xxnvATZifBHdKxa1OnfueXHfq7Q/Ml2Zl3rD
CTnydmijL0ZFgikZu5eUFxp2mDCf8xS7r5LECuydaESnTy4ZpJzxNycWNFTo
2MlBD9pj7YRLZeH9IGDgPBktMwWt8ZaZlyR6Tt+YcWgZlc/kmC7ajWWK8kO9
O3yGuA7bfzHsIPG7EibXHRtrv4gZ61OYbdpVq34SLtHoIEpIsrRUxjMtKEgg
2oc4RHYWoBC1pE7YNN4lDgWROKihLVdf7a8dEwS48JPwicKuYimMsgMd+uj9
XnI0P6ROYoGNpIxoNRO+bd4+H1XSInYaPMW+fIwNkexCqzoF71zbp4bENebR
/xf+K2zdpVP1xR///bKBGhzvkdwzzUJMHFpmMPxzIDQc3dCAlSDt303BAVGv
aRtWjXMST9ofI4ARqtlBRVJ3/xY9TYKywK3TLuAMo2JB5eyV/Ll2x/Npi/0m
VOKvcdF+s8M54fUoizUWQyqpcdf5vJFUTh9KbJuUuwCWw8uObCCXxqZprY0/
tRv+vxs+QQUW3nwa6JLd3fB42eJarxG6nxAB/PHx1K4rSqYjY8kDy+bk1xSD
SfVTG+4LZVaCGOFkYLmme9hfBMz8p0wawk9svHsCHG/7rXccv+y/hgz5xEJw
3Gy6cV9A7mlB70QqQJh1DDQx4WPn19p006dM2imhKE5ZagkAzlE0Z8IRCrt6
xvpFFNLDe+tI2G/vcAiHAnLbqWysbTVkjwSdbRU3eCeMLprZIFeShvO7Xxyv
EbkHMIdspYROB6Esu49oIHsuG3A69v5gngdpsabNtoSaBRSuH3P/a26qt/7y
/jQGGc/LNlYv1QqFcbC2d/d/rczooEz4FeuKG4JI2G3PCMY07evPqNpitxjE
IolobwJsPWZfPX9sCODnDDmWZMkL8KHj0sIxw/PDntLCj/fzThG+NFGAfDDW
0LOG5vf8eFrZoo6Qjpki3mhFxcCvsS0rjWI6jkL2kiJLBwwyJIoDhJ+Pem+g
en5URxgZAbCLywV7idSBc6lZRqoWqWhASs+JkuwpFM8YNVviiB0EL759VND2
Y+FCt4gcHN/G/mnl1XEK82sSdC/6zBEIdRNsBFtlmZ8XTH+iN5Af3wMvDFpi
tntzoEYV/r7Ck155H98lHM0FI84mjK7K6H7SjwaGGPeTmq/OCn11OdJUawv7
ya22J8tXBJ4PaDWmDBBlSFWhjfPMWftRuFB6XSVDxsDTdCesmNaRiNmsh22u
MpqKSwDaDVF6LxWWdx/ZsAHJ6V+8L97Ycr5h7AEMpTZ9Qd/iDo5jRDFdqn6m
6lwfe/zCA3jKtrbHdmZzzcBvOMABTeSI4hFBeSiCBF5Ff15jXk9eB84/X0M8
c/jXNZ0mt1LSN9q5/iP+A4IedxUiXLPQExG0h69wmMNYI8hHnxzSsO8rrsBK
pJvJu8PZTd761k15V8p6FRK2R14UQxLNT7V8sqUKRZLgV5vW8J6/KjcpQPS2
k9f+lLcI3k9dZoZLSnxtTj9UK99+r04rVBsikuvEFWiINzNbIqlCToPWtp1w
lWF/YciHgG4/X6rNcz3s9j6KjMcL9AtODDy1RS8Kxy40x3S47SUUfzSCXUkF
YhdZu1/KFIJpb0QA8TvvRREa2lx8UNZpQVegb2mLc4yC0TC2RSVCXpWpxStV
9wNaDyPXFcE2wFoWmb7p14KMJcRde0mnvJSdEyXZG5oV039+3mRgLkjhyBpy
lO+pu5LyCuhCQBmIRSKTr/U5iuGByRppaJOp4O7lOBy3G5Sb/UvmaDGq6wmE
lK4ibZPxY8PlGjIL+IgTmsrLWgZvKarZku8dWOyW9FxOWjfckC/5snXiNIu6
afhTdfG8NCpoW8vSNV4SwVgE1Tzf/7Zw80WUlNOsLT0OfOGrnoojqkqzZUYx
oGCFEfNZNYTvDQXuxzCs2bDAz2mzUnftqb21WNklzu0MXs/xMGLlVP+IFVgm
/HyujVPGHc1EJqSd6fQ8DfDkLf3zWFpeywFqbDO/M/P3mnECwGxob+44tJ+O
+yYu8zp7gLgWt1Yy0W5ePCGaHi1GS3TWYtiMC85Yv50pFWBhNYX/pEuoxRCE
QFywNVLB4K2uFjKhnoiH3/9FoQN9FSzGkXcJwi+9/jSWGfZtC4TQTO1NkOwM
agJm3S8BDzY0qrmsfSS8JxSFo5X+Jg0uC1u7Cp3xD6v8eFtKpawmPc64XTHt
H8XXcLhvsoAIirECkZSsbBHyC5HyR3tzvYDHOvw1rqb0Ba1tnZ8VrE936Mpq
iPfe+Ty4xb/Bdy4kVmTKVemVQBoofYWQtaD8pQRKEvylHoues+hug0R6vOrI
llqQWOzlJot48n8OzCKgKEUnVYpJrG4kJ/IwrJFJaelr5zTUVyQv4uUjRzIP
HW3FY/4w2DmQ0kKRsKh2XkXsEuT8PReJiZCwjxvrhgVzzbWZ1r8YM83QCQlt
/UNUi96m+4etYYNDtUmb+zdes0C9uoPT7FLk7bD+ewUv3yfR/XcS9wh59xBD
wDZWm0PVmJQY4lCuwURA/pA9prAgcGDVg+XfVgJa11EBAK0XX/OG2cdV3g12
2oJl/Pi939T0D7JKqluDfo716OrCl5LiPBbww8isVfHDcbuEwA/3gr+wrcRp
NXKgmGpGpRwdO/4DJ8rC+aiHtLUoXC4r/Gfo5seeuaSrF4L90d6rS21UyZDp
ZsGNdcl1CsKbrr3dI9MhO8L6ZoCoBKntQaiUxsP7yLSQjeObLptqBpk/xCSJ
8OPpGFaSJEeZweazJUBmM9fwlhaPszLMgiQMUi+6wgffsTlfAX+BGxahn+Wm
OLaBRk9v5NdaKlVUo5E77R7HhELwfBsZb2ln/yrUbRIwIwhSupK5sDSIOYOH
BNcb4Wx9O79Q03R+spTSWhjzYF0mDGxYgyZBf38m9Jd5WQ/oafRUt8Yy1Vkf
yrmzqWQN91bqoDxatsq4zH/2uR7X/RFXMjYqyA5MfncCwKIzt/0EX6WUzNtq
pq74u2QnFMgpl7FqsHcnp3+fDrSKx/SKVAb4onyJKyeyu1Rr0pJzDWMh4+o6
La3OPyImgYGH4Ihgv0LysdDKkd5p4hJLXQK+tuVS/kNdLsZxw1SKbRZSB4/5
iwrHGPVU+AB8xl0+dZ0iYOK3bPwlSmLe8EDr6CYfSna5MyCDaJ53fznpTCeA
hgnzI0npu14bsC+xDqzbB9OcKzO1k6aQUwEWM09dNXPegTDXmrJHmSA8vWei
K59bIMJ3x5B+K6TCORigruOxA1SVNkeyOmFnGFhoGJb2k6CNz1uH9S/eYdP+
yJlPvibMFAWfdcPdXyXAiED/BWOVZOwlE4FP5sU2fjtYsVIY02aQfpFFf79J
4v38igaBerfdKlB3kMFSnRFa3DXFhLOkpZ1tYr2AeCaQgOfzjeccbnnJgVsr
Qod0qagn682oSv3sPF58nMYtZGEd1KPsBGSoGAs1WqVVJGmowfEb2hNf1S2N
CCfXt7oGvb3CwV5e/9/63FQxROG69FwGas9RqtPPnBg7P+XqZDxE6gtR3Qfj
SQ6wrnWZm61bAcdovXzlOS+X+SrOw3+p4yL/mnbHfSBq2Bq2uEob2Se8h0Em
FiqY4ZdcKbsxeinOaciFUKOhnl36dYI7r0RsKRlKK/UHY8LysQU/nqptjomZ
tc3OjRJwl6MVfZAyxIzABCWb/pBvYATXHreARSRayaBb/hHwJu1Qa/4KYtLs
/X0A6NvquUwEzSGJ4sFeFZ0i/jRYf0LbQa99kesGR5uWxvzMdASqoNmeQ5u9
dojXTb9r0t1BCAmS7z8xaMacIeg6PELwaL3IbEAXAFX0fl/y43y/djaXx/ba
LnlYn93r1gD6Hk7lERBDiJ4GUFygHpbWkehANauF1tTAoNorHuQsNmcXZugm
4Da3rF4pItXZaahwwOXVcgjJuZ82wrNOHrdODHMKvpURnElfdsw8QtLQiPMg
wfxTh1HM2Af+G4tslhGF6d7FpbWNf2tBMY5muIRQnbo5HH9x7X7AX9impokv
4k32rVLpgNxakoY1Hyz31u5rGs4ZiesSAzHSC+Ogi6EucGqz2VtqjtNng4jz
QKg8tJV4Nxu83IXdQb2lYbbtSnh+1BlY2QnSx2Z3yCvus39m2PGsjnGbr0RL
PO6WkW2cbOKo687mms5wkA50mpnYXflwrvafkt/WJUgaZsg7Oi7Yb39NgWB3
NMKbwbmijdiPH4MbsDtjEHiFnjl4cBoxKWG2Ssn2P9LBekhX4fEQyK6eftyG
Ve4CdjU/asn4q1l8dnakQoPPSJTh6MqwGdv7wju1hgAQKpOtq61HtWoWwv+N
N3npiJTlDGBzcIqt85YeKuA9D/LWdcvXpCwjJ1LpTRXnCZAv5M39cwhYUTgd
BLnp3gBNS67SjqkOg+hJYesqNSVSJ5nZHZ+cH06rRjSNK9rSgd8kHC/jDWuz
wRQPQpK11WwdD8LPTyFhWcKrbeAzExxM/gG402s0GzTbw029x3fLug/EcLt+
v6uhYdkmSPJoBP/3pGwy2FAdzuo+OdXAgMCpfjGWfN9T8vdf5yum5yrGB2P6
kU38mQZA0weFPx5tlC0T/QPGB0NVW2UpnWF934X3aVaVb2jPvTvxaqFk92PB
9e+5jIapEi7Hft8Sj2y1xOvXaQikQSfhDoWzSewXE02n59rmTJ4AFE4Pt7iH
2CHDNP2oTxt22kun2FBUezySSTtZxmqcSvipRcKXqEZmj3ZbvkUfUHm/gObM
18lB2bOP5mcAnzawOfiDmrSTJzYjUgiRfB5RyppRJV5u1itTQy5/gFVKbq+T
bwTvuz8MbyUmaOI2f5JGT6EQhzKUOn7mt10iLYVfPjEka4qZI9j75AfT9wM4
N7WJ0Vj8jtDZefrrgqFQTi37gNlqooWVDTGrtymTCF4Ra+wTEvMJnhzeaQVl
3V/xoPG7UFNLxCGqosAjiDlYI4sPzDVX4MDn7s7FfLATgiasqJoWKTVeuu/E
ycaQvryoRy0JRDfvy0pXFhTJ+YwQJB9KyzXavJx20DgFq3X+amNTiFTRMIVu
s8mbDHr6+kMWO84bRlqC1IKQqG8u1YCWTYbcpVaLPVTVGNkW3ENcrgg+yvuJ
LComlDBZ6dzNxoq3Aj1CrVAmPNrsYRxUgNIjdJymdyNa/Kr2fMA+q5o4MPQO
XZ/oInN+1M9dL65I/EyeuftkDmTvvs102eVQjbXPnUhNDEHvf8uXhvVdXaiS
KB8ehVx97ag53lWaDZCRvsp5oEIlluPv/AZ3ZUxcXG0BjLoBnZIyyMaaxoTw
PQIq5nuyJO0JeFl5dtB751jHV3JiQ6S07fU9NnCnmbgk38cgMUQ2Tp7sQrSx
4XMprfzTUaArC9IDYw/e2rkMhhjcJwjRUgA96VHF9jxDAdSYJ83weeDIaiR7
fzsmoaJqayHWD/vfOs6ndoj1cKwZoIA/egojvpokrKgPbW4WfGuIDXnQ2btV
yulrm+UcwttLtwHaTA7s64I2b+3AqYCpDc2z34ZSNuPTIkp5FIK8G/OsQY7/
wKZTjA0j67sUwddrruIy/08nmVnUFLW39nRzkY+Uuo3a6kBPdP5WY52HtNKP
PljB0RhkIvY67ge7q85LeU7CfmpUnFq9BCma/iWDDEfzyjQuinN3Y4rW5EOs
59LcIsoYFlWH/8jL3QWfqVbX8nWjMysZ6SknSVaQ+cjoy3uo8/NgjHwTUGQY
bf7GoQ2XOi9iZGqG23mrzeVBQYdRJRkAYHEUlwjVFIV7Vp2ArXRU5rAlwmkC
ikN61MH8CLaI3d7icFKbr8HLqSYk1mXJKL4eRppY+bgwLIKEqWaRVV4WfL4X
h2O6zqSNx+t0u7DAEfgazkPw9tF47JR6TmPuPzg/EIFVIs2UTSHloFsKk3Je
jZhoBu/PIuw/oJuGt2PMHZef9dxBqUpe6Wjk7V5hIIFm1IKu0/myDhkllhBw
OXaOL3p0TDx44byZUlyKYxEhIEzpExAzHH8ICzz9Wgoh/lq0jB7g3i7k0hMl
C1+TswwkpK2jOIlbrZyrsZpSpPlFxe1cUE/NLAiOAHg+m6jF/+pSbAY/8EQE
kwuW4C79SlDXU9NNxUm+XcsybETLVpz2Ej/Zvgh4sY35vu5qMZnBu+H9WTJM
AQEUEXBo5SZqVnJYJHCsTLB2/2fOlRPcob8YQaxRxfjHBfreI09Ng3bZro0F
RRozF30H9hUr+E+8x3fmLlnvxQGPzQR4GgVgxl3qp8fdncChp7o5jnib5H+K
g8yM7i6lbutzAUZ3TJD8W4ivEBsuO4oChnCTwltVeO3C2oV/56k2q5aixqSM
vpcBj7+Do/b1IAArX4YPDMUDddORTj2FK8jMrMxuW4LW6IDGjURiVVcOVXFf
OlOKNLPzsydotGWhhZaR3fgOXZIBhbXouUEKguK1NVzfhC0AMcb33VFIemrY
apkMt9mrZKXLzEhENc1oPJG18Ie7ArEYZJjwJUM1fj4DO/WWrekP/Iaaq8Dn
JAwJC8PG4sZFaYAF+uGhTcOorHMyUg2TjvKE8p21mA9+cwlSQ3oKNnDXmIqT
9UOOvrcBYzoT86GEq0xqJLBlRaTorzI2gEdENouPxCnbvHODJkIBeFkb1Joh
nAsdz/xhT/xLUaPwiyvV3zR0v8XNDMrcT0VIC41kZVLmdvV4R0+85/XvZrgv
tb/drNs2mln0/A2OzG0HO3Nnm3dhsmZ2etKd60uHnN86ly/le6vlJuz5Mm3t
AnXXCHG9opQzs3FQUN0hAhGq+XAZDQzklq7DSqC8hLK/mO81pYytuk0VoTUS
++S6HDSbLUo/xqoC59rlFhfZCr7Ob6HyfKfTs/qUSPzHfTj6ucUJxxvgUDdS
u1NUfEOzUyisNlb7S1TtVb+VYPG9nubUVXW7Oyez/jGdbK8/axXFP6mufMGT
2uyG8sIy73Zlt8RaB2dPhhM3UvcJBz94wb9psV3KGH5no+a5dZ6uBUC/TlVZ
0/ZwhZb2w+EZPHb2/EiC04LTgZI+J7tgW7og4TheVQKQIZ1iTX9PQopYqumY
Fy6AecbhIGTe8euGucXEXo14QcFF4qMxbbtdNB4DhkQv/tCeSciaLSc7Cwv9
B/GTAONbkg0RUWeiofhOnuYr8iROvcdXd1xUHn+UHqycaAgHqaEtl7yhV5r0
erdd12nRyLHUUUJAn/IKhdvIneFmVeYi9aoYSs0tuUlldsXBiDHs/B7GsHQV
Kfl7Q7/+YJ8I6ty4gxxzAStYk3KXd/nR2JulLGeS3Zu23/AyqzVAkyXrRBX/
T4tHGZwVYgoXTbG4qRSNDwg4XYu5R4PJgpNNoWjBpwMpD4D7fT5dJ0OKzab3
dvF1iatZEMq/+GCA+N+4S+1jzr3EHI+CLE6WpqqtwkDXiI2ogOfeFTyikFso
6Ggpf1kBHma0bF38WwhF1cRikDj13bnl/grwTaLVPmVZFIhPMomrc0vneJpb
bgmMn+NI1c0QYYA78j1uhBZdY80QTX5S5C8u59jX2D3WdTwZB6DiPBnato7x
E87+j3JWpyHUs5qPXEcEvSZcxFBHNth8yWfK1i8soukSoh2BhjyL1z5B00vQ
SfCqY+uSTvbmKRGgqDS2lSu8Wu3liNngwT5jzDDkWb6fQXc5KmVOZ7pMlDtu
ZeavRsM+cAgSXpe7qzH0DXuSxyvsho2uj1bbFtOIEgX20yo2Q3pmkuy+ha/E
hI3fDm0G8eticHkkoxaFNBjSfzwWL4Jq7edz6Z1XKLQ4h2WNy8XzijODca5a
ivhZ5oOSPtUKUCB1pC4kZ7cK3VUsgskoznQkbPdBu0XsNwtNwqN0hg7gHHeP
X7n8I0TBB7Yh9dRVnYKo1ZvBUZerXz9fdconja3kmiqUaaS0TJeBt2KqmjKR
euKpWs2PBxLO9U+dwUZBdlA9pdNRr5ZQZJcPmzmV5UkDdRmUG0Fzlc8AcMsB
d88lZlnbjQljaTxmTDlDpVh8AsjQOxrrfWbEJFcfmHi7N3LRJc8RCdz6mrTD
oS9aY9pV9Bpxd/iC7wc75FuoSo3KrdfHgl2ZvttK5DaCYwoZZEKPXf2Hjkfg
ipFpomxdlf4y0Dnxp5zu/mfMenjPh3EzLfauCFrM+xF881db/p9by1AAsJDe
9UlR8Hz3VamJ0FrJrznNpfQMzlf/dkLzIGe3LGV3gmmhnL0kO3NJYTN6hnuF
N/6TD5492gzSgN6yXbrK7aEkuf24IQfQ7CH+995d0e5q6Jt6ZtDV5XQYI2l5
TkDborWTj6MR7oRvh8AizZ8L3UCN9djgZD9r29AUfidz/FivsWpXHolWnFMf
OQzl7qF5gJH2rblPfuM9FZcFGMH8lO8xRhv9y2Vb5ofM3BgmPjUxFnm2LdZa
ZGrhDsjnito5cAzayhMp5xydgS1NsprRPSkUMn68qs4lBrKcH22WhEx1fK6F
mfTovIH56rDaxA4k05N+0MAQe5EOnCLiy1Ym9fGEf0ZW93tvkFuzrj3TGQVs
KtitkRE67RMs3oz1UU9VLSQPAIsPZ2Z/o9hgnKuBgFLfdxM7QgxqxmqqlW0J
fXT6GpMAZlCZ/pgl9RRIscrrQjk7DVW6ZGi7KYw1xao/xdFPheeIKrPKr/VQ
WYmD7XO66LrCSvy4pBtRLDf+jLwEykMwe36HHkxjUpTxDObwEDySC3XYM4B5
48+Y4TKgeZySTLnHmUENv6pMwyT8wlFvvOuPMU//pm4y/MQyiO3dGynnce+6
zHJzw0EMRuqBn4nvibCu2xfbJOMeh+Deke58WSuopo3Tm2EgASqkgXzoQN1N
3bzt647PpqmPfGahz8eG+yoYkfpkWkkMAwzlxsM+gB+FWCFlrwP45RUdPgxo
+6VC7CRlbbzP/TU9IzQ/imgeJknlBv/b3xIlG8J5UguCORECIQHz9aded5dY
WTJTBUSXD+HCffrm2SLBMJSbdMjUutnhTWW0s56yp49lXT1VLZT/zBbcygmn
Bd3lgNQ0F4aHdJum1uI/efeWlofXKm0pWdOm9ldp4nA6wO0OGnpBj7yxRIR7
9djE3S6TfBi2SnJaizKQFz1M96ny7hV4nNz3y1nZuAcgh5emiyUZA9Tf/iX8
7x7C1RUYJ4JA3hDCYSXYixkvA40SrD8AhMFd/U03xSXcxFqs3dBGWJ5/M0eA
DFBquh40EI8dSdwa/CU4zsT8i/KtX0JQzBAXWjGjfbUjzZzuIlsn1K94iT9g
V5vyzNXCUS2D2DyKNG5+bT2rwkig80hRB0IDBtF2/90pqTlZKDHNoAn4UNDQ
oDbWG8UsdduHyks15NI+a8eFSIKvR3py5a1H6BW45mT4O7a0OhClffZ04Ckt
PKJkHA7oHWIFyM8Z1Yf3Eh/At99ZzI/weK+hXi3yCScLndRg5uDpyP8zh8W8
xhhvg1c/lc4YoMoi8jQUG5iyk9GtqCvrv4/4Nq6sfwaQ9mPLsMh9QdQjgo3R
Za2ZxQ4zT0DArNdnDXyRhHZZ2oOP001WygAXEIluGKRvPVUnqzUMJ8KQbGs6
j4NVRZ8hSwP4iVVFcbPD+MpbqMfWkWjGvI+mpJuKM8B5gnoIFrXUwx++N0Ak
BBjpzch5HEYQUznQpb9fXaPveC6/j7Hu5EamDvX1MtLM31Jb9a7GHflBBJoP
F/aK6dm4O7NJyNozS+r6gCx7C5cah2DbcbkfdNq2pcY8sA9aMv4oNt0jFlwi
jTu2Lww34Er2AqNG1LK0dYdJCLgjI6PHinHzzJvojW5sPSiUupc4kldjRJBl
0lzOrNdicnOMEHiiWHFuHpPg8XamgFDgYI2i28Wlw0/pMc+MuYJtocCFWLyf
GHE50yfObmL0eHOzfXEAghgmsqYiJgntV30CyoE9KSITUhchPCbyQOIPMASw
A6qtLMAaMC5Dg8mVjv8GyDeu0SexEaSIDr2Nb/u4U3miX//O93gnQFH4g/cT
1caTEMOw2VjBZPmuomo1i5HmRJ/tVJi2FMHIqLwm/O+wqW8d/Wr9GqF//Y5R
4QmyqhOrHbPQwannah8WFKPO2xGeOspCgKZQjPhi/Prgtt2mAtLMHWuZ2i3X
5m8/YRmCdr1bKcWcVnoGzvRzJfMzR2TOXE/DRzqfPHVsHUftMQWHHGrh3AeC
wXPLVD5aaQ2uECfJx+jMB0xhE3i5QxPp7xWwbafA/sMJYMwB9OM/jFpNfEwy
sIvP8MA6hlfHuVex195T1PPB04MS/uoggY1ZnpY2AFGUqeZB4PWofeCalrNw
fwRT/omEZhwJWvMvBAIx4qd5krXwYIqR7S0K8fEcxFjNgTDmT0zrcl/TJQnr
Xydk+jWV65074Wg0FyiTBkA7kJ3hh4nrg1lXjxsDt1RcB2XECd/0uTGlvWVe
VRwEjIB1WtsM9bJJr4PHWiNmNAUTAAfPl72KKWhT3eh6SZd+AczHdMrwIGYH
K+CVz0e1UaHkTFbY19MXjKRqZYXUmFIv+LQgc6G29IpIy2uTP9DOxjdw9Ti8
LOUp4fIZjzotO0Xro8klbxrEByg8e5Qr0wQM4AK7y7AmNzyMZnk3zgG34ul7
tisRnZf7G1IqYCunwF+4x8TI/mEVhu+xIH8ysG8aDhGodOcz9DrtgW2Hg5Gv
K5z6MaFo8DiGItmfrB36+4XyHXay3cK2SGbCNvq1YrZUB8u7EW8CKDmFzcK3
0U4LY5gNKSMl++JqQZY0AGR1hY5Su/aVVC2L/4GacNA/053qHN7bKdss2DAc
o+kk+vOdB4YcTSAvEYiA3mezguSbe+okfKtdLk6aWDtxMH/yv46YYLLrcYEa
VBfkXBzDibbSVt7tM/k4eSGkt6FRiWcXGHxZauehMaN1uBQUyqpZK/JGK2LP
7gDywdAJWC35Ye+B5u3iTRIzkcx7+JWO4eMf7WWuNsaFNwIpM9w60+Ns0GiT
NTRkcnf/Lvt7EybXYM7dUNl732Ojjbe3E3N29Vx3rhfHnbmgI1vAsGmPWOsy
Eyu2mHGShT/vmjQJ02vE17UeRlO+CKbMNiL6VBSAmDycjKP+l2QpWrEpXjP5
IfUQIxd4xIVjBunuVCtSnzUMYfO0bJO7FTGpBmoL+9T/H1l7iu+tQ89XYMtJ
EQJQW+A19Nc6/ZWOEjcHzat5Ib2SFXmeMq+Q9k82orRdg2/CLWQkAzZC8Gtt
oUaq3LRTbbqEQ3gfDPlgc6mlrOmmnKOMPGibgoD5d2hXYP9pRdAJ7we0oG5Q
3RwXtBTM/GZt51cMSeVt9qfQ2kYuskf17GlH+DyUOoPoqy6sVhErGUZOqY5Y
nAEH7PYJvpyS5L9DThISjuMtanXJv60lh4hSQrDuZYbrbVqfQmQMTHklhoDS
PpVjnS0iKXIRfU4ZX1vYGYsGUCTszm8i/Vi5TICHa73RL5JcPYVnw39MpDSH
bfARFHD4SfAjWRpso8bcJ0AZhU4jsHcREUsBCDjCg657h5I2qrLBW//XeRlx
xQVNcYgrlohQm94CBWdjvt69LXHGLUU1YqOuI0KTPfNF+PyBSIWKAIjircCU
mDL20TgyDsbi19g0kdqtyIBfE41HhAiA+p1y96yoZqm2qcU7VmXR0yS7H8CX
Q8v7l7uA6t7xuq6uLBMrsBwVkIOa8fF4evysQx4haXOcPkM1mMpSa9Be9ryI
9I2Ef6i3A+bjq7RydJn8MhUPqzWqXIkwCQdNfbYvfYndzR/jWNU7+4w2G5jU
1Q8drVmKHGblmmsqADrI64Zo2/PrAk17JHe/32OJWPPan8r2aOZhG8DyrOCL
FbqAH7phZazbc6gUIny2I5kzfMrRUJlflGO+Is2zjPBCJFExGJ3j/RYuH0FA
G403rhIqFrGPaBTu0AAsFdRCc0Gc1qF0xPjsoLv7Uf4qxTY+HOhLetbPzOVN
b6+hr2ZZ8XOZwqxVD4Q1pVSunB9RTAspRPxhtBceM7eALCdr8C+fkHzM02cS
ieH9t/9HhTHBqNVvOtZEzQLNFuWetONwrh8N2J/pt2wXVj5ydqLeYZKtlUpY
4plll5dK8vPzOj2vkrpxCZ2dbKxNDl/+NdnXMgF4hKl3NRrwflZMss/IWtgY
gUIgKF3TvYl44EWxH3tvgrLGoIOHdYxxxgU230bvcWdwPI59xW8kBa7r0jUU
eY/7gR0nyZd6hbCrm11y6CAwY3PWz0ibjPI32H+53rIBaxOqwo3t9PLHiFn9
M3kILoX0fibj/Cb49WGs0G94EZD6wsC5ca82B1Ixfz7tj3CQ9NOa8hXaNjgT
9r7RqUXT365KqUjrpZ0DSuCzLUHV/bIjKPI/LeviN4BoBMn+Ugcr3uieZ2X4
MQ7ELwnjZcn4L1kDoJbx4AP0ni2DM107b2N+kdbwO6RYk1uqP6Fb72ZR8wC9
0kTGxzlr2X8Q+fr5UXiIkoSkaU57IpvS9Bvm+NftxOlVgK3I7ygON4aJ3Z3K
tn3LgOZHiSz1udS5SgZkKBdooX3dNwp1eapmrV503YJES+Wp3W8wlMTd6tBT
J2V2nqfku+MUYgeO+hT58kpk8xbrno9B6OX9Oene12As8W6sVbWTcQW1/rpi
LR0jB3DIbgiVLRCuNnYZEMutje8RDk4Z/52DIcSRAweAjh1Bl2+CdT9ZFq+s
vhJKNzTToLq/ZSu8gMhHt61VfAfWb1Wq6dWbKNVVaiEc3wkfgJOFmhEnf9Us
85tE3EXQj8PD9V82RcMRH8L09vsYfpP5szubgIwU6i9mv1RYEdxhgaTfDB2M
v3Znt428xDoikpp5yXv1Xs3qFWzNUB5vbO1CokBawj6cwnjcoEkAVGk6oJtT
/shmx3rHVIdyqnUYyL/UYT6uXrOUVSZMndS8Yg/O6NRPfXiMG6C+U9/gJn9y
ok2Z3pkSxcsoFyHVLrSdjV9VlVeBTFOxm6ty+tygEsws16weBhyye18oQy2p
ML7DNs/CLO01sUyr4wZR1692+ZZbjQ0T4VQS8mFFqTWMTymd274B4m/48znS
NUBionLKV6OufTGBxH2yeTsoTblOtpBxumEAejqVeNkFFU4vbscbg96BZmRD
jF9cDVg1IpejlSMBQFgbFK8dhmkzXZiTspkqWPVbwSNN9ySEDpNg1FelQIlW
9QDo1rkSwPxvSvvumOX4dAAkLRlyp6b31K2tqpptm0Fyna/QzNMR631+nXzz
147qYw+SrR03yqu7DE0E3wEL8r1mhmyfKnVSoF9tSuJO2wlA0cpiPvx+kD65
RI2MRFZksA0s2MeAVQ1IpoIDQpaWR2qcTe5u3DSKDhfJNd6HO76QbIiWHnHu
0fYTIu8XQYErtmchqF1KwG0FlqU4qDV8PBadnpXPnxylYVnoX+82EQ1Sdo5i
k2tjObjx6DThHuRiYAgJvGZSKiFTRLOdEKsWatohPl9adqi+rHnXwpxBxJPl
EqrpPkw7vSfN/kMMrLBZAWqnhNMlZMchCwl3iLEFrV3uaeTLdOC3v52VkkxB
OtvgFbmlEo2/EkklDv3ZCl7mPZhIMhcSNnmcw/b4kkBT/zgoeTT3copHkplp
2H7WkESlzCjjGtgG6bZNQWym7CgkjHQdjuVJF6n62eB58eOkkxmaHZBHmILy
bF6oMmE2REHRcWRrHej9+AefKMmnYR6f/S2vT+P3bpCmai4JSyJkS56+5x3v
Z5XjuynMAzSxZnUlym9rxLhXVLBx72WO1zYAVCXO7jCoRQgY93YfdwgpxBSa
mbe76lozVGaUqy2yYqvQPbMFPaS1GDzFGOaWmmTXOAf46fbWH2bKzfacSD3x
d0aeGZZFV6JNJTzeZxlrpCqaoavMNVbROpNJba+y7stqsXlglW+CaJR/4k/2
GWibM2vihDjr3tLJNmxojRlvpfzg3MIZ5qhHvZhmeBLjUB4nP5PHuzgjv3kW
y3h+EYWbJi5AVdkzZcB8uYLwe/pcm1LTXAaB6pQjP8+V1/pOgagJ1Lebv4iv
prx09HcSI0ck0oEnPRc2cQ/LvUzeUgcLu4A4cFqbsFyHRY/dDQYU850VpGHg
FIwBm+SQH68hEH0ZhdoxuFRXQtLkXDv+zRevdya9e2F0UiNYK+tlDjxGwWrE
pJZxNFz4w9tl06bc6q3ejPLaXB3htSQlh0RaCX8rMBWR+lqs0kPGarqpq2cK
NvX+50DBN89ZXMHs+9BgSZl6d2tC0rHjGJfeJSI2+PivhOtvMz0OxOk0KWKq
8LaTs6u+saF5UnxnzYaLnYX6zuXu8Kda7qMrebiw8PB80MdrlAPsmylyg3yB
5SXxQru0ua9uhvgKE27WwRVblFGIO4/9MQWvcxeTeuExrmEElbYMoLnMx+ok
m4dDkGUDKQmxDaNE1KCEoTf6jFEWkm+bp6I90j4N1IQXL0WT6foreKMKxS52
gZM5R8+28dM0PTWWyfVNUYjykfU/SR6MGOzpezKF8LEU9Ck2Hd4PxujiMR8T
tp6raQiknJ+WvMMtYz9EgZweizR05OlgbbHELH5wcgbqbNWTZK+WkeZG6qRi
FmycIYOZtBaizr8Iz3NXDSgBmc7iNHHkTrASebR4waKFdjv80LebkO3Yh24V
cnzLss/aW3T8QBapISvCiaGgBu1XEXkyGGrka07VYP8rYyR7uSQ8zppDs63t
Hy8dTvv/NRnkQg+iHnM2JfL0TPKYFpk6nnRaMm1yLeZwIASZmYzSq+aOuysh
vT3du2tEdhkF3AAQWGAsbitadxIfQmC8Zd/qviMbkp1LKKGYvzNzVUdOqk3d
Omj6afhud5x9lc34F0n1nyKixfn1K1LsOgoNK7yXEN7RvDIAMc3BciI18+5A
Joyxf5rCAPYUV/CW5cygXjCBh9WG5VgxXdpQe16dQZ+qn0RrY1jVLCbZNMFL
L1wPnB4duLREk/C1BRiCPRecmeGSD9MdiY5WNU8P0bhOpL7fLF1TfzcrCi7/
t/ApHBnbGy3AzTIzJaj97y0ncyYF8sBbn2wM73E8lq1J1zRW+bM9WrqWoDX7
UCPzJ05qSmYKaEAWcocVixfUxVMTZ2HEcVQI+tJQuXHlli5FKZApm5CSK2H1
cncYrGi0Ils95wkn25NLtqC5nwWs3U4gtKmc13QlvJbDhmdNqstxYXQ/CQgO
8LIebmU9SX+ImjSh5kPaGDCoW96TBPiCCgsMn8FZeUUeFLY76PoSOtaJ0YXz
HtFJlN3ybXktpV/iX/3Dbim0H5Vdk9xUUwTNRD4932ihAEWlX7Ro7UGjpFM4
cXuamXut8MLyijQ4CDMaaleo0gPwv4My7SsGNdGyS/xo07LzNfv9bUpTX9QP
Cy8xV97NIaxn2TqR4LI50Bz0NqVH8nu5P0z04JlazSc1G1gjBeS11T3I/L0s
g0a4vPPsYA1vH+MLJqAnHUtKuMRPKOWFOeO3jo3DNMRft+osA+UHDINCCEJU
pvPtWl08ohiS0ovd+RU2xv9MamRqItY1AxRzUZXom7u7Oc6UKwvJjKe1Uyli
WB/SxfjOoPDHkQlr58ycJJ44/YX7XLsjOum0LaT3qaeJe6v71iKhYL3csdkG
wcBgEK3xkdVip/7iB+Oxekmxpz78xVfsEsgbMBd/F+WurCV3q8jR1DuxuFyW
EIMWzTHKd5D4bsZjgH++1TiEYO3CjT5zf0vi5vElQD4RNGSXWEo+a5gynJ4G
I/jmTDpGtrFojGSE75dar4AnR0Jjm3UEU3UvWy2E1dqCe7n77r6UT22tSp6Y
WKpwxw5b79xPhR1GG/c3SA5rHhsTTPyqYeyAKxl1yIzuCxy3+NhskADnF2wM
yk9FQLFR8ovBC3fJTgHGA6iYV8jCbYZNKb5T51QxkE5+xLY5eAfgv39hnCFc
jWJWWY86uClwEQ8EUNFktX8bQbHIE6uXs4PpSuQYjv9y001iddeXyrLti0ks
mfRnGhZJbDNwYmtfaWDJN7gxGre677RYK7bZncGIA+cNCsHH1trUOuEUVSZf
ucqjwD+L3jnNuUEGIyclRD220KsaaNLjPK1VJ+/P3vOg/mAnKnNy6PUH7/Hp
tUjqBqFwk9QsTdxKfrUxIcijtRhscNcLK6h8ZEY/dgrE6kzWThP14OWbhSu3
4YsJOoEbOORK0a/vMRUhDaN/4nw4+S5YfXczMzaG0HT2cm9FcfWJVf+cKgrV
33XHSFKcKZqvtqrIwiwEJalWmKZuztUdPXrGFHee8qnY82PHe1J13WlmlY+Q
w53/sUbcVLICFZMWM8ZhfBrnFHmWOTl5GKczsMtovLnKdWJEGIJ3AymvdpyW
R2ajMsqUlZ6BSiA6dvI9oYaIbIvZCMAo5rgRfpwVU9Hz1+Uwe2RJLnEbgakV
6DWabzZeFtSxS/2l4VsZceVkCkxJX+69mHzXJP2oMCYEnGo7NpQA4//HjQmB
HfnOvWjQqNosQuygFd4ngogwKCFBVJPqD0Pp1YU+FqjDIZ3TSAP8ajbSULeM
HewfnvN/junt02MQsTCRUyT+TgE7AQzaX6ET+VQVfWP8Yl+PSPh/coree6Q3
oQi+RSWx6dDXrB3E8nnVWY7Y19sDSmPcamPQdDMdBlJK34JhKoO3QQ5g9V8q
HBF47b6oLbxD+1yiPNDbfZP2iRononkw4UlhEAPEiOmlkwT6nJ+GluG6s6Ow
qcf82a4hPELE8lYmtvtFaLLe2rd7yyQTNgtRvFJQsXrK/b3G7vWlzjGhY74o
3p+mIdS9Iwe3BG3X4EO7LOtCpUt6ahaqK8ano9D3iTQCa6DaK2/BpGBwtzdr
q6gtQIFnN/UOgjP/2iyORPRyU8jmKm4LlBuwMX7Chw/bHg/81TzPARjD2Jy8
vrDPL0e2Zg7OtnovFkYKmaI7VCiHRGIgHp4jcL+GvDaYZ0e2dGo3gkHogL4i
QE2/yABN7IwQwJ+dfFSNLpC/bFm3pn4CssHaSXTcVXVXdlu6RHhnk9ykYcN6
KN9aQZvbuuGyYV/i20ULLbkr2iP/8kp2xdbW/uFQvSFzZGsQ1UR/ikpymjVN
hr+qIuASNR+Ny7CxFN/Xb2kktlBJl2g+YvduzV6Q47Zyz5YiPMLVRFGLnhjr
HMElun1IzqBr6xEN3j+Bc0WGGT+wR0s/PpfiYorPo5RYiH0VuIeSHE3OpF4h
V4ee5+WXof+VPYWURab50OtOnj6MSV5+oxykJ41Ld5AGxGcYTs+JXw2vlhdN
MFemEHolU6F6Z7MChal3AymTPs9pUroCxsxUIERc00hLWuSk0kHbfgc2Yr9d
lbqA5w9QCrZb2rXSAipfJ1zuh0FbTp1RjiglMGcMENO+mtMJNHASqTNBo1HX
c7KK4WhxCqaBxreC1SJd2NTpFDjfCWX/JeTYsRfOLD7m5jJ/IjLGN+ToMCmh
6UeYWBNjGxoAiDPq7HVqo2h5WnfgoLTHXOeY6LXbnjPzWnBQ5iO/bpfZocnX
32hyKshR0ZuQgfTy5l5ihHS2NZuaUHSrduVzLalFU3Yz8UAVuImFrRv0Gc0l
zeVxnht5tb3DEnZxOEyxT1bLNAnd+qXZAWqpXldCRMDEbPgX4hEUU9tW0C99
0Y/5xw7qYHJwCmrnJHkthny+I0sqEEzrQmRQQDBjUhtvtNLnh2N4vw0w/rpt
nk9w/+OaZmG0YGPt+W0lb3gesSvcfIpzZ/SvSSgNF/fYAjWi6bpHGHgLm70i
176yX/uVrX5byupQlphbxdEdJeEgRMHmaMhSz9MyvdD9jJiTO0uQNH92F/XZ
UwaB1ZNqi3ziIT0FdfVdtekQbbHUTxpP3789RvVG1PJRVGWHxSeX7nOAHjFT
twO4wuSjbK8q06IL4QQMoARD2B6HqkwIIbI4IXrUgnKnUCDn3rl5hRh3xXUr
Sxagqh511a+1vLGXaWJyC3hNgQQ8D3SrQihJbog1L/hASqYCmE+c1Wzmd0ra
kYWGO7svmScPOSIn0i/KugEhcgx5i3ns8uhKN8mkXfe2HL7e53zWeIANJxWK
eFjrjLB0DoW4lHua5UT4iwU5WFmjop5MFxCw8TSNlKMt0FbSURzAZlzf4QLr
feBcyU40LIH4syVnjrz3AAl4liE2n4G9D17aSe53MtYH81btfYS7SSV/CcPd
HuemeCJHl9G3Ca6UcUJMIW2X2uC3OiZ0ob6Ufe8NFzMtxLs4oBd0YyWkTHR9
G+ZD6a8TRSqAXMXYLFV7XjwWZzH5CnxPuPc/D+Lowh9QTFxEi3HUT8VGTdAc
imkBkIHXF+2br9cZh4qQOv8/XrwEYu5Xy1jW+QfIzD5OXiBGgc46Mz7MtyJ9
e96qRTev97JBaHredLbyRkMQtyVbdIdhc9bq4X/8ttTkmzln+Q887bl4Gtfv
O/zLwMpqmkAfVDnTvqlE3DyoBr4f6M8s9SpWcjlI+Ly5vsTFWOSkW1+mN6OR
c2LVmhAgQ3oUzMCwqpVYqpUKjodOM2dVlTmwDo2cyvty8WSv4bWqoqXqRi7c
V0j1SNssWyK0MOYdQAPmInn9X4YGlJlkehMed9HbE0fPOb7lA3krz8bJ/CkW
anbdce7pHhs1XtCJHJs2ryfrC3Iic27ZibbJBQTSUHiWL8LFxaLYfWCH3ck9
HMV0FUASOLuaATia7g486+LYAEjUjMJeQmI3p738y53a1czZ+sF6qSkXKNXm
wFxS2Tm6JDM93Q4Ukf66X/C9eqXqPadRkVXFQPQD7/z9t0hiv4qlYPwlnrSo
xRrH/+XqQalzIe1/iUTnfyfJyYJKB6nlcG2pTVBGKDnOcobTR1W9vLuECyPZ
Ih6Zg2x5BmQiKYlRRHYFjO5VtkgHa3PcgGXHpiZpLiFP5xdv09sQ/wcbemvs
a1EJTSJjALZM9f4JDLOE23Zv/Y9qs/DqQKe7ZqtVbRfjggo3u6UFQMEj6tT8
OH2ZuSzjIHw44LCx404dRpMSPopuH+rIDYNZHteUsGcDirDBNSL0l2NKoTHe
vnTa5L/r0rTa91k9aqB6rcFjpiAHhndM2ktaJyLM+xrf4T4fUlpROSdNdRUa
6qr9Gc8laCXCPQoD6h/Y4QL/ZVS/4H3XSKYVQwhaf8j6EFt9+Xgz1DhR7lOk
lTp4e/PKvTkNKzB7bg08+l8kKXWluJ8d7mcKdCCyJeHUMuXfXzT/Gukdp/k+
t7iXlLeE0AkiNWShN9ASn53VAaCRvqBITe54UBVER9V1xfWyEORs6a4aCO40
xwTfu5fPH4K/YCVcyA97xItbytPiXvBtJqgxkTTChM13rksfpKYffo9/3QGz
TDinFW/BN6+RUdRhh7PtBzU8Xpuj0GWZiNIdQ0D910XDQXAA82gcFngA52Hq
dnhzv881qygBiEYRfsE2C0rXaY8Ic0TUFSy5Rv5403E8z4Q5+XbMDuxltDzK
50nFKZNDhKj8+mPqT9YEiG0uAOFlDYhKXYJYqT9CCJNTPuEW5GGwIsGX4xXp
dJ5Em8VqRKbZbND8PNEhXelvmWsrJFh7mAVbH+6HBRh2aG/TwT+J1OZBcggU
CFcwtnzLd07QAzwzt2JYoM8rL6Lco/58ZSeyDOc5OMGr/z7OA8t2oLu+kVuu
k9gWRkDy2FalAB8kKeolstBcNHDC7Ufx0MLUCtjhY7csfqDbI0TfEtD/kBE8
fYEnMIYgd5v0GypMcumVik820ZIWDF/AIV0XjlvwRRWUdBwj/GwpoNZ9vl5L
vXECBE1Ah2CX2+Un5XSXStm4yrbr0aBg0aVNbGFvjKBtnibSPEnc2wazKhJd
4tY9z7qeE0M1sfw4lz08YRjdAr2R0tJuMGipx7v2ALRDlbNpLBxHMbP5jct4
pJx13wFKT4RHRphNHqX3Cb8S4+5kp0/t+z2yoJhJCenMFfJ+jNMPWmCHK8Of
h5IB9n6tqNi/WP9MDzwwOJ4W5yfVCcKScgVQ7VuN8UVZrHzLQznO0Ds5xa6u
J+M0/8oewoYYjooYPXgbeOMFAKNRnYXawF2Awgd7d+o02j5XbcAComtT54ql
Cm1zynXIKZGsZIuzXIIBRDMNXXbSVUk4h4/N3ddBOhuirT6240zYZz5EAftF
FZsGDesHOCBZCFZ7u5jC9MHGOS7TtaNCczLfz8SpJAH6WfGF/S3Gbl+Uvnlt
wXryzADhThav41nO4n58FkCRVjtvdiW9JiGCYACB873rvSDE89gOQYHDYa+o
B23UORlVLsTaABQn62EmeZr0K0rI6ceUQwgZHpp8j4ynyj0flJ067Ptmte6J
OjkMxPQo49TJ2fyqK8/OKFBWqBxtbzDmfyr1Wq9IOIwYMTGXXFX+vhaFV4Ct
CP5mB8zWYDR8KCv+VFuxdwipT3XyPzXX3Rm52oK/ktkjBp+RuMXJ0G7l5UQR
HhO5HYlgJ5AVekbn1K9Z7jISNRk4durCwYB8LjQLZNAcWXeNaUA9v7+ShOrU
W8OEN3E5o2xh6utZPxO9HIAydTRjDBJkA5xLRt+a4VgrnDSQM5Spv1oNq+8S
TvHh5k8jlWdg2+6zk5dF7CLEXj6dGgAZ+5/mjlehDocY/faG44fDRdlw8iYE
N40PfKyPywakV0S/KwWJSbq6fxamc7N3yEaSRiQYZyqengWC9VZQNeNaX96a
qJKF7fs4/7itrhCooJUbaqlj6a8oOwMRo35xxVnFvLiLGPxXYbmGULTta22T
pgbFoxY5pi7uxfTg+BUdOwH45eszazwD6Zyvx6dq12y6LI1ggde8WAG4Fv4Q
XivA1Ak1xBd/Ic46Dca5SQMR0rAtzxOOlkW9xHclwixz8u0p8N3nVHCWipxg
0jxqBAZ9ctORCe4rhialAbdlwrjFFHSdvmYmI6/teYBqBcn4IwEAvgZ6skGa
hBkHmNJ7oszT3kre1SKZ4sy9PZWY0hCXqcI1BFTnYJpuok13KFb2FD4oCtAW
ctrIdkZ6A9Ald423Db5wFI7G1L1vyJIAtH6PfAaGzvOumQQP9cEO4MrkqvMP
yJGCvA5zPruGt2mJe6pWGFspuzUORitRgchbB6waIWDdPd4/Y4BPcWe8P13t
lV2KqwgodTx5SXXUQAn3OLzicLYO6xbJOI685oW1zYnOTsW5Nyng5U0t46hf
SoUGTNha3FsWFakXGLahW67gmBiqpWuJX7Sm+gQFOdSZeAMZMkUctjtL12cM
waa61GlvAL80hDVsMzUiXgGt9d4cRFMJLxW0tf3N0ZL9rAXGvqxzkrv3JfjM
OlrDxZnRGTutupCOjz+cWzmU17HeAdFGOtZtjjaywwo/t3bI3y5Gbl3zmPcr
yzZtskcb6orWQukdKws9owRlWxOt0+D/k+3cxLOXLxVije5PRPR3FCp5XlWJ
G7BAvjunOQaM2qgGpDFvcBo0nqEb+Ag6wIVu409m2xp5KkiV+CQtwSJVSTHV
byHI6I99IBJdOmz3pDQ4uc0ZyjNplVplWs4qGl9WEqKKt/zTUAbtJC9B2inj
FRWe2c88iXB4IFwf7NvWLJBjwwKxsxJjiXc15Ibh+tPVbwqgnbwGtMcC+qUb
ebaEgEsq19BeFzOzO7k/Fd/Ad7HC5WdI0jtcwh80XXVjfhzBk8WuwXPwNJ8z
NCbdajs4JaD67LT61KdkRoukFU6JU1U8EyoQQYetB2jouitjSgOneTVcONBu
vvE66un9FnEDwhwLWtI2KClQgpq+xrTeklwhVK1ctYLiqchxA/KaJBEIYLyu
LGoP0flgF669I/DhpevAyEXeikh1F+KhxNxVa30ZnXlsDym8Sp6ZdULZGf8N
/Nrrwr3+W2GL3UwrWF79Jdr6TyksX4bA4h0oW2Z6XeRF8XKh9y+mUOmTfNRR
4tgRVWIznWYoBHXzLuS83VDuBLhUxVuF5pGi29YvDMOUs2nXAXEwAo9pvpTj
y4Lbrmg8QkhF73bvNMUw8ZLFoz7AkRLVCOwjCmkQ3pjXNxuHZx4+AG3GLMWg
YnXYUCobd+IyyCJygNJObZMCriA/2XYZ8uWcxOSVwgHrrppVYxh6MaxUcuY1
fzkmHurfrW+kF2ByFsLJ/5KfmmQwUt/bi9s0t5HIU+DxrY2QIv51wjJLM2eb
lebwiLmvT3QINUry7y6KWLtV8ZYMeKMy21seChN6r7xcPjCRstFE1lfpzAhn
HNaiUf8g5DuNi2h6LYMbq59DLyHFxaHwSV4fR42oLHp0CKIUPCyM4SVgH/q/
rbF96h0CG5RVgWBOPDASou0Gn9+001CO1TtFa55colGItave6OA7jq2432dR
/W8X6VamOC8CX3EEZrRkxdLcZtM2TD0DtknPdtF27HLl4ievC2L0E6eVCIRh
y4t/px1E4fKG2JmtBu1tBqxqCrP0QKK4vw53jPD6WmlDy8rxi8BoNvG755tV
HjfaSrxniX8okIm957guT95x0akJej+MarD/JhB3w95r3hMCOx341lAdZ/qz
g5A3g5DL+DU92LjwSk5uCnDi1KqjFfWPTsXdoO3txYJsTI0V6VrjDRhs6GOu
TLVbqZl87y+HS8/zzNmJMhFTJ3Xz3eLgduBEQydIEyJ0L/CNgF6aXhSfwuGy
Ako2O6B+f2zkztJJhBkM6/dxinTZpN/vctrLIWMRL1YQKgJL8f9BQnucsdFc
PsQcsGpD/LJSkvyoQx1T+pamcYvQBi7BvtwNF++yj6pSGYCiO0Q6POKLYeN1
SOHaskKl9gchPS3D7jt2XBmROzEBd+otGlzGUVdaPQH65Qk5766WMjG+3aJP
BeLgdJoLa6EtUeOQ6+Xvaj4qBJOb+dutUf++R+sPUZb2w/6tedZXt+wIiFzp
6JxywzEVwc2SkTQldVqu88MfIdCFImPqgmkQC0BOJxaiWjf+23GhecSsi0dE
iqdYmNLO51tA44ghamfSadvkJrwx0606rlWaWBLcJOz4CwNM1u7S1J8QvaG1
xj2XiQEuKWHGn/lXqH0/a6zKEkZlRxZPl5lYHjcNvf7o51g11qDfXt1VXnZU
NXCIrls2udFyY4+UGZXWZKAGkF5jtzGB8Em10cOMrT0YnRa4zTvi2Efv9Pxw
FBlcMEVvqlnJ1CtbwhYVGLJiqmMMg1BVhFVKMfrkQuVe/0bvkMYBRVqlqToE
stg6EG/2kisDbv8XBccjl8GlPaeXjfW7BVvt+idsjO6Gi2eKnh4IGnqwrh4l
iPQ5DHhACr4FzFBm5fq+u0IsPy7oFGhZzhw3wFCyyJNYGh1hEpMsFRbfEjLl
WJbQCkfI6C7nHJYfpGVnSyAgw1t8Bhqh/05J+Yl4BfUda2CkuPkPBK+HHe80
5rUIj5BJPmmTkSZxBdWqCw/3PcuqOXSyVypYCKHHDljCB6KvY3ocJYQGCN1l
lGaIUm4CqNb9IH+/t15drriREDLgpYFiZMjFDIrR9int0hqmwBy3sxL6sRYw
CEr+AAlk2Skm8bIW9tLWETIjmdE0xtrV6UGCL/AsfQzhMX9aADmJbE5VVub/
lEb57lzffx8MTB+y+ODNkrLik35g076gWTtNGyNYplPFTsx8RESf0vaR5+Va
myjw6RbE5hs2dgrTgj+qB5T54tr5c0bgzcRYaaXBUdC6KYW2vUbWgR24sTFm
uLV3+mpyVvqf67L+pInexie+uThOGBWgzzcqRZE040aunBjKxRzgzyNaEloZ
ngAdynKggakp/XHhFlhfQ5Tp5p69OjfU0JHEDaPs6ABYoWxacBDpNjX4Jf0A
y2Rbn6YNWxsLLq7ObdLTvsh+39QBiqc1SimeAzrkhP6FDRORAoAQCB9n5vh5
vKwqIvitHfGsX72QzKEKg3gOFxFiArDDHGO59+RJXEaKqcHKeWmqiCcDDuQu
Tg44/aHDoV/8CKyT6z5ZNUyYlRFIEX45P9rVDe1R5Y5pn2GFo8tGQUt5xHwE
SXtFc2gM4FkGsy/eLRaRWsc3lYYrqC/agBc0bCW9ylLcKekaUOoOdKw2gegt
xLo83RsxFtVkjGx1D3UyzDF5nXB6tetun0GOwc8RiMtFHlRt08y3kQvULjDU
KJhD3+xNiwHpD1aaqWppJZzJt6fbf9uwddXnq6iL+LnxS+vRipGN6x1s7k04
/AA4iyFAyDKUeG6Mp8BWtIb9zzq9dHfO3v2+HUpsD3pIwthdtoSBELII3jHF
2KnzZdTZqAwadonztxZgI0ze619F40Fdq4lr9PwK1BIWm4IvAfnUjVEnLzKx
pVXzRRPHcdobs0NfG0ZkDFPnUtmMKIfq+r7GJb8Aph5El+gSf074yHGFJmFU
Q4TxpdMW3qzeMULduXk4g/9VpKDVcmc5tcNNrL+ToRlTQ6//ke8JbXtLhMMV
vT31DvpebgAN6rbcKdtpF1Ncqe2RmUgAzOt5m0ZT5LdDrobs84WPUaojMFBw
JlQEE7YyKPZLLfo4+H8Bwrqrf9MHxbewGRzZ356nEkmCsQB3R2EMrAArs+6O
TpL1AyUb2q8TBw7durYpw7CIulp+V5OazYA2Xx2Zda/78cZWWRPlFFvSLB0g
NMVUX66YPMN5FgoyHMY2N/dQEUArmKd6VDICKcBuBJ3koKXerq1hiTtpQ8QO
shR/1dGizVNuvJh6c142xzPKj7K4MWvBPVLcxMr3Y7E6pDqHABeGKkaBOoBp
RnQYXol5HZAv4ZZIouh+7AZkd5VDPiUJ7hGRZ3NdrB0ezbHXPWW00d6NrgWQ
h/FLnuyc1yolvVQMX3sD9LgsUZI67EbhP9cFHWkKq0ygv8WiPG7Gm7SjNcnu
hIleKOvRXofkqO8/lh03cy+c4yjdLTM0OI4AB/kEPa28O1JZv/iFbClOfqC5
x3d+eyzT9M5GOLEMQALGqB8qffosjp0qyE7607RKgcTVNrenYwvXOE6EIRTf
5p2JXDAre48n50OScfkxtv4PWQeTsOTbi8JTSRcuSGwh2BK265pRzC8YdYRq
dV7siIj+1poahyBzEBWaqks2B+jVkxldc3JkIDQ2M51YMI8iT8+MzdCz9PzI
S7DU2PmqTrdMTiz7qs8oZSykbnKfgeoE0L2BPQnrG1rYSgyWorjpLPDBira3
WqBOkMmYTlEgkpaLfhkS9XA5hQT/FKHPYvhPe9S86p3dLX4HzDyZE+ovyJSs
4CbOIvgcDgQ5cbP5QsP1KQdxPbib5T+sIFHCG5oNhAkmQ+dQ2Cv7BjiqdW+J
cCsCIoAZ9PN5MXQ+7CICKHS15I6z6kQNS1n5DuLNOx2ZWqj7s3Mun1dZZwQ6
HoIlO8Ff3bvzPWn9+FNMDpzNpjkxzJo5HrIRcGK3kq5SlKjB9xL5f1Y3+/wM
kslJS7kvbHIMMBMsumqorY4wqO6ilWPNk3kj4vLi/LmQM1qXq9aFypacL3uf
MTOERXogGG8bhv0j0SJPAQtZFUcjORfNkS1ROTM2w7zcbYMBuv+DwEmcDlHk
sROZLUnmgQJrhXMErFzgFHA+04rXhmsCEPADqngDP4RrKsexiLvTxikEoCWH
iLep4853mtgsfnosOhoTZ7tJr5YwlGDZH9EHaUu7FV0mEWkPpZ6110Fm/8ir
l8+Kre/CXWclZFA0BrwfihvWpeGQioMrq16iOVS+sYM6S+fCWDbLktIgeOXi
ARc/XBt7ernvNnkOJe+i5BoCuBqw62ER8UXgwJdMWPXo5d8QyKFD3M6QPJmG
J6xVIcqTo/epGgSYRqhtZwzMTLW2xugV+cEmFTsOXiLqhN26Ni2xPR7zg13i
8+1uwzAdHFnntb7h3qRoLK3LdVvKMqDJkDFNG50lmAA+sZ2nq3VzKA591xsD
+H7IrKniqJpAg+iSZaqXdlIB1v+G7ZHIc5eyNWnh5L49zeJe54gddBiikYJ0
aGdNJRymna0ZQ3iBpqTgqSwfhS8+p3eZvJJ9kAsJrPCEQuHsg0j2vbIyXKYb
Zzba5pa8daClG00vIZoaocqaV3DAHrfI91+xUwW4wNWT+MmfTTcWtT0AXkFi
0oAlzV0S8otQ8vfgVy7goTTePAu9uHfgNUGM7GOqvITpM2KItsghYZYPKmIB
VUXblbyV3nFfThJwp/jpkylCTwhnmd6BaL8FHh5Ux/qLt4hIntlG92DeFU8a
9r6nMQV2j0WrYYNSImSSNYMjpMxxh+ch5mZyKE3RlUDzBDJmRSUH9Slei45B
iR5ojVryaXgCIUsUhqZgDL4pc1xFG/52AJUUJlc8HzXy3rgcN0Dzd8l4cqy0
wCci17YYJ9XfeRnX+OPDWAeVd+9kfVmZEPFCoxWKqLICNj4auVFGFb2yMxci
MQ/PP0WIulV8AiMh4sHCz+MEc6Xn4/j1kPsZqY+Mr8smTDq/nB0cnjtA9M5M
HRm7cRmYKAFGw8w1DaYrSdN7SfJhA1qSvf9Kor+3nhWVUuslcP5q9NqzBotb
jNI8jr03o9ace1FBiKFu2yXxZOxLHdkNJhWJRuB5RxgXR5UdXPuvKtEe7gE0
PKz4L+4Tkos/PIsgnwIYGB+8wxppMpBb6EwsBNTFai+pHb4oUCIkeKjJ6oza
YOkZteFE4QuDuqDYIV6yxErXa+hOV2gqnkcDE5E0oap7Y36V33/cyOk7sOFF
br15fTOZOyaClXFR0xW7pG6ZGuYELAbfOMX9oa4rFBWDqH3PNyaMpiWNXIqr
NHj40C53iOnVa9YtdR7s4hs/vgKUKjHOBfRAU4qv3aKK7CyRM4oSp0NHrETV
AxkdgtNtMVHOxfeB72Gzeo8uHj5YE9NrQu3Q1t38Pw4+73/BLEdUzrbu5Tl4
VKVrJgekrvL/0oOM1zFPWkKg7e4WzM9Za+lmliXwpag8h7j8MZT7YblERPqd
qrexK2M2PbE7cRCwHEDDfWfzFMGbCyl4vksaYztmlpQeWMwG3utc/IfPyZkQ
XvXEJzTbS5aH1/I2BQmKh8w/yPMUKYiBckR+LK87O791M7hhl7GbHAMGf42J
jpn/tBdwad6y/7ZboFM6fo+n7ydZ8+timhCax8CCQh80l78g5AhPOQocKqlL
9KRF5x6SKgYPELM46biGjBronxZv0H/+fr3e7ztq0AIYvlUeCGYoltzBu98x
I2nSYcPdPVKqBqdZyErCOzR3BPi6BAKZkGAOR2rH3YbsF/7kAv/7TZ3pegzj
0QU0aTXV3xNmr34NlldsnomYbT0Xj4d55n+hztKnRl9ntsRZ1oNAAl5c7pYJ
RASmI85dCGJX/Xi3zD8bOMnTvdkwmLo9jAfd2thGHSgtG97gWrXLiAWlgFG1
HVxOQDlS7KPSDl+2yF5EExzLlS2hSW2AUwVRWQ9xt/fIGDrMHcp+yP52DPdS
EgRlkFkOvwjv1vAQZsyYXGkQOgHWaUdFi/ixE8bFR138dbGfWZJY5OjykAuL
yThaH4kK3asglrV/SNDa0xZgJZl7Jt0VuJ954d/vXTj+4e5Au0kGiPUTj3jt
OsuetQ72Ns/GOlx+wOl4rlTkQxk8BvIC7EGkfNMXr/x5KV334fIilTjB7cgC
d5siCYTYqBuBD1/i7bspAiI1G05iE2OufJF/bogWncAYYV7yzDFQ5kEmxx/7
1mUWSuhzAh1ABYcCdQJ14B8/uKKyiKHo2MpnOy+k75oS8oHrKIlKjNs9Xqly
O8UKZLZ5VmNcSRmqMm8mwc9QR3BF6vK9Idizy6L59pRJinPlBboWEx6v8huz
eXB3aeezbSWHSJyDcCGWoHyyb+/TSMOxz0Q68tFl053VP5LoI8kEGOh5PBhJ
YmcHbMHFfpl5HD1g/BydnFV2USQoYt/nT5RHeCUwjl7bpTBz8X2SC7rxBYXn
1ay2nPSdRbKZy/qtznewHYveUX1GJ48qLdKaJudU+nNyFHPpg0h5s9Z0by78
O5vGVIo+9jmo10oB2dwjnHddsciXi7EVmsm7RtpBrUqr5k6RlWFdvlo7CAgV
W/utwsFYTFlwygIYVx9NPtnp2JiCprTQgKNJrB+fqtWhur76/9g1L0S6KHIM
KhWY/3Es1RdMRleqbraC4UZW3ky5yW8Q0oCwBZoumR9g6UHdO5dL1kvZWNh2
QhCc7QHcCnp+nfJKIi8e/ss2dBYUD+WYJpXUjTot4a6lO8tPc88oZQrHI++/
VbMOws8SclYUT3wACO4bxpXKZUxtgV243iMnwhGsXNz5GCSkzL35/cflkFmE
ShGioVY9FNKF2cUHMAV7r7PWYfHA3sozUj1FMKoGV6vmY63ENn+6YaO8QI45
O0M0AgEUHnlzhO+YkBNc1hnQgZnGB3XCxtKb6n9zjU+z+3i84Zuu4xI3X1sh
qJjXK979+8W/w5AuRbl8/mQy1T22BRTjHp+BC19YoVp+E0cRl4CfKEAlsJc/
8IkgBCPJCIPHiN1Cy1xuA+40K4GPcC3DypbB5IFGuas4FmEQ9wXLkM3vnve4
v3+wv1b4VhdvdMUg66HMJIZtImSusTItzrIjrPDEUgS23/5PY6hBJ64BQiyT
XxWGl2tK4ge/cyfLWjxlyZn25ptyq+Lo6BlBYVLEqTUrPCTVIlkMzeDvLXpB
mkPv6RUY6CDny4682ds3dLs9kPKIkbVy71bUfPA/iXjZY0yOJmruT2Srrobe
gdq8j6R6+ISd7cySFO1WCeLzNM/BTPCmeq3BHNjrQQrtz8oCg/qFUGDn96dw
ikyvaeF2MQp+3r7E7pgjCvYjS0Fh5FC9d5xdTWRKbba6JY39A5hRXGQHD4XQ
vvS+vHRmWJVmmQ0PRXB2KaGYzWQCqIkpCRJdUfpmtvM24vcCKMxMPVg3D99Q
biwSNWGjlhzdxhjrB+5zd+mCuo/pVhyFrQbitaLJYKbI3E80dH5iE+v0qFlx
6cGYsTbfYMxwl/Dp5HDkLZAy5t025dcOHWdqCiEWYJO/AIpRJ8p8KxSK914X
o+oRXYb4yp76Oqcu5U8zmo3DUUxi2gMMDG4OtOdr7aN5nNwryA8QWajBljxH
vJtC40isVLtYsDa8l/FY62WmCuKOAYjrCX/qoWhyMT12EjN9boQiqs47uyOO
SJdvAy+nBjKaxsymGH7veSVZ1nb5rYDLqPrds4yCDVex+WI3CdSpgk2NkUQC
JhNjqSm2cO8KHLnoTrjgKca+jMXsJ2+8pQ+PtIvYDdLQTWHtEQKLlDU3YciZ
DRYdzopLywSxf1MdGGyHiDnE/WpbuFxrV5Q1rWkfuoL28ejw+w6waFF/iuFg
HvycSixKS3e4RsnIk1Fs1bxquCdV4+KYp4r7sJGJgaqShM9lm0+Vm+7tE3Im
rF8mlx2Z9JeUp1fHQXkxqAF1E/HcuXqKcoJPBPSd3eT/fKR05fkUdTnnMQkf
PCUS8aNr+5Kwa499kE0ZsBsMlungUCWNf2aipV5gJOfFp0kzqZWccGgrwjke
atSpU+KGpNXtQFPLJlGWt8N5Vgpj5wY833I1npmUsa4HFtX/j4x5+cb6WOVV
t0znBRP6GtGlTDDqNDZLAIUiTaR10Y+kdJwh8cwf03sEyBoBZL+ag/xfs/Ph
jZa4jGcosUbIs+UPZ7jYmAavSZ0sFXld4nW/NNs0lLHDdhbkg/TPMifxXe5m
uN7aRn6R7i9COA7uSKjVwakU0wEuLXhJUv8QxLQAAfTErk+WH0Lr2Q7FWJpi
2Zn6QIALDZbk6qhd2HKHzQMyVAulCKKJ5gm+3qIxC/5hivzi+sUiAOst3I9m
LtuNUfKqSHB7TOMTyrDRTSGSHmLYk/niVsDopDBNjeVVEE9GL8Jt0/T8F+AE
sZll78knLykc7KEwx6sfxjah+GVTdiqkigN86+sogyyrpJ6uCVwTcSD6xqxn
zx/kY/gKo/9y42bwzlSHrIRI+CFro+EueruHIwWcBc1F2stlBKytf9TOUZg9
2rrFARO7JtZInSVU7PQjoKCUtz+4oJEDaXbl8vnpRlT0vo75s2xGRvWFoaXj
nujJclQt8kdCoV8rsy64KQXpRphLzgKmNqbEACXggfwBvduetT8R0GtzIYMR
JuBggFZ+JwGKqVAwyYa/AxyjYTI+K8JCdYCU8JMT5SCG9NhKz5u4g1o6179o
B2MqFDEpE0wFizUmzJfOUPSg2upwo5jgrf13e/M8PQgkvQBAuQK1eB8DLb9y
5JXrO2uBCwqWcXTJb+8ZtdEYG9w3afjU3hu61IJsrkf1jJubMHJ5v8/tjKVz
FUmpMbdEZbiiUrdypRNCbr9GCXEKvgMMsOp3SFzsixVTtINEUqwA26AaTs+N
b/zYgave8bYggH56cokDJWRLYM3rHkBm5iSTD7lNOLOOUE+HOotWgnse50Gj
VPv1AtDmO35rpM9gGCmhvXwklToAjtdP2PGbPZ1DzVN/pJu6lzDjQ+SL2zUC
BXCoagjB21xVP2be5LFdL7vSSVey36JMiCWfaRskBytnJWewrmB+IdnivTna
1c866sJ8N6TLxs2FMtnr+UcMbQCGRtDd5E0rPd+ZKnaBTXay7syJDxAmB07p
uV0LTcyt2Ve7v0QLl/006e6LeBYgc53u4Nx3WpaGd/DmjuEr5PbZgMeXeDcs
ay/5t0o59vzZAMCsR5WPDRDGPcznGPAtCH44Kk6YwUTRiOyluTlNsB6mdbtr
txPrJgxmVHWyps+C8QF0cUyLYi9wgRm7A5tjLB6OvBaiezfFTL0Tpmi0NrEC
Xdjiw9TmAWrJ1ofiYSGeDVqzoREa6SaokRhr/vak5Fe35HWDwx11fxrSyozj
j7MaxmZgsZWGCSc+tDIAndUEJN0MZTTV68MWF8pxmKb+zy0/yzS2oFPQH/iP
BBZhY7smfOkX3dkChB5gBL+/d4FeDBb1wNr0sc5ES6U5kJqbYYo8+3AY7eN8
8STVumjTIqJwfGTWnpPHk/cBsZ5eSg0JJJoxy+WhVllODIOL2FADuiSadk6C
db1p1utZ7lN8S1T2+rJgtnYCwKAmHl79sDuyHph0D32cFJVkCdaXVUWQKc65
LsC2eFweZcR9xG4Zt5lg8ET/RPmJ/UrzkJ0zAc458gv9X0OGVXlibzpBgZDJ
9gAWtVnF7e+5d+JKEZlqCmr9efp+bB8SJGFok3bTkd76ji7cFOGStsRMdXs8
uPIpHynddp940YrEydEV+YnX1dylMvRmno26RncEn+puSGzObo5yzvi0t1rM
xhGrLxoOeFkIoh9usw02L4hIjzeWoHXw3pNELjBE1JEANkNdiuRWDQgG+5iD
FM0cOKRPwQ2Y0GjXFQ97RCgEJYwUIwEfXNmq8M+W4fC3DejDXswKtG2UT04h
bKrOK1uH/ebovz2v3U57yY5sB0CELrm18vAa0HhQ5ncIjhakUIVYhK1F+QkP
N8J6TTCTtp8gttmqqRGKqFS2YK1Fyg36hk/heT27BqSjg0wOK9Yro3f9Fltj
SytWzezIDPz+2xC4sHrIUxO3TFcWQY2tt9/urKRk0JSxbxMr40pLioqPUMd2
3py/cVrUCLQkgZiKkNQpDF1MhqN9LSTMBTODMQNZvylk08PSW7wA9nXHlM0N
jYjagb7JHmwbKwllV2qnCxg8+X1HcdQrLprzW7H9Q/U/IDVgjKw3kmCM6MP4
cmTO3NgrfEu96EV9JF+n0QLlugW19FotWGbYI3pxXpXkHlb16/+yzXLPMcN5
B4jIQXmK9KiUusIwHPnmlaFWBBxJeQKWtBNaN5QGG3dY0ZXCsrBq31iWNUg3
F/uMhROotg1dHmhphFNUxvU2UkNf46p52iRs/bCT/jbP44y9marlYlNr2iD1
LiSZ3+enz5OpxwrZAtIKtxCn53l4kmm8vFtXjC0fxPmnFr/czEOgDsH6yF/E
0nNMOs1osW14t3u1nEtY/R7k6nJvmRwscWlCIiGPDyso3A14TUKx/H53/k8r
ti/SlSQiomIGQHRPOXZ6rIiQ6LLbjwj5wJWRa9Aj5seV+Wm93wRL8yE/LJ1x
EFDAI30mgzm6xllEDDHD919Zn0UWzpYnCIv40mgQMM8Wf/nW6FkkRhs+NY3z
LRsHLY8MWeWMwdNneVexE2EzXDAvS3G7HFLmZbkBoCpDG2e8UCJqTHWdExue
rW79W99/EsYQyhzacNQS8T+IgMRwXYvzeAzBXDivhfXqfdSSGj45x4mNReqT
vLHhuW2JW7u8R4JCLXhXIpoimk09Lz4Q0ZvZ3k/uMj4Cn9HLKXC6Rzi9GdRa
5/ca9d1wI01BT3QDW8zsnjzL7/iDhzAeekjPDNE1lI82uwa25njbPFcFK2K0
0Vg9xIgMLLnLhOr08PgVF3MLtqBEEDUUKIZPC6lH9vvLGIsDJ/W+NGfYA+zY
lqLI7vbHKaqFJW/oELp9TikIjvk4cHJbPjceZorUuibKeVHxFzW6SXyGr3Tz
XOoWXbDTSjn02JkkMvlr5SD71uA8O6FgCMO6TLQaFgKCNwwu2FBm7Y3bcbpa
HXz+r6MM+WrNBxmU+0JIJ75GpHjXJuq+5vYVtA8ZHDZqfiRfN4aqIZxNZen2
iLrcs8lRLLyWNqumUCeYrQFYZgTdRg6K6ySJNvqE9gQ1moMkFfxJf5mxTGQ0
RZ0+1hnvEGq0dirYFJi1r/tgA5iKcVjluV9ZwEXETF1rS4R6BL29ZYlBq7yn
QptQAWZQvKGRbtK9VuSF1LfpwdGVy9CJad3ox+/cOsXxUzTFnW5n+m365fVV
eHwk2lIGvYxcooSwqWKuDgrGtTdOEOsmONiVKXDOe2dKbFWWbjXlf/mo1u0R
PWzJ0+yHnP8gKaG1HpdvceFdrj8+iImjj7aRs/+J0SrfsC1rl8nNXr45B2sJ
sPBYOKC0xTQth3YlE5G5SkKJEUI8/IlSdK3MnnIPZEzY99LYkKl+Yvv8mSNn
tdIlCxg8GomiY2lR90h/HHiFgxa5asgCXNwqcSoOGxQPBihH+wjAZ46CnC3/
oIZ4UeTHBcBqf+bI+3hy5c5CtZZteDEs6JSpsD0n8G/84u8P7ibnFw0KkOFl
I5JAwl8yyBi0KSc9JRKgmmfwL+FOXQrS+wLJFtqEF30RsEvNhkcpPZ4FBs7J
Frw8PZijiG9cxwlvUySvA8FQ1K+YF2k5NfHKMGRI2VCYDCqaXDHQTgZHPec7
pA8JWY2Q/Fox8ApjfTz52fU8RBJixQQnjd1wqSHoHc5577xAgD0/mDolhefz
atBvZUcXUziJo/IM76I6rE61eKH9Yn7C5osNo1MQWAxzFr6R0IT7noKSXc9D
ggvULiA50QlPeuizhFHyQcv+FjomYXApLIklNtK+ymR8pOoFuvidyMKjT1A2
CgYRUhSKVq21eUPEEptbi4icmHjAJIkQb8osHm3wfiKrPTR99GHvdCagAjpI
6BXjWS77MF/m1JgteLOyUkidJA3RO0xexQRkGvIBn3FxwAvlEIpB4Uef2MGh
QiTf6cc+MMPexSeRr9lj6SWZwVb3PIvNIiU8YGwpJgiCyehKYMN+FEZYzL9e
AfuGuvqkvOCoYe31TO50yHte1zFoZbRXxac3E9dE2G5e0klesH1ge5UgSD6n
GxabGR8CYfeesUFuPr2xsHVGjNE0o6x/ryResBj59HBPSAdmdBCadBIPVzW7
ITZqmgvHjEq4k8Ja/fkdw2FiLoe4wIyl2TSdt0OSdBkUds2lkqyd+SpiwrNn
dyRj5VnjZtJ35+7RAt9FisVL03WATa3JgwiFngSxZIT2ylXkmfDQb0BrF15t
7GHyxznE7Mw+wrJ06YK/lPJKigmS7KLikuQcFU4meTK+UDve2UROdJM7sfNh
77a3LwCMC+ywnUcTAzMw10LEiQ/bR3w5Q0ak2QJ5+f2kbBi1mA6eY0IYuHZx
U3RNQnWViTHQA08L6SVeA1EWI9+wi8h+HRt3jvYflGZRaDqxqCh8ithhUtnw
3cAeJrp+BflgFUVWBY1Ajqs1bRwxtlS5bCbbWd8wKdE5gr8qipTXWqQbsE6a
Vq7trYM4xDrl9yP3rMergQud9YBag2jxHcfGh+Zjn7SXxld7/7k6few6wi7h
bY/ECZSIdTcLGMCyXlqz/JyzahD6zo2ADc5G7TikzsYsYNdmKoQtGxXP2zHI
kV/bP4wg6Cqju2PTlqxSpNrbPwpihXSJYyTULpiy2oE23luBuxl2exxc6tOq
Akp/Tk0DpLROPMAiiHlvUiZ1vJKb72HMF7AT/m50haDKjUikeY4HSRfG0lvi
38YYERVg9gW/KMxT18xpirz2C1qqavQVTxLchJJMsBrr1Ahu/vg2nOlSltUg
RULz3i1p4cZC5PYqPQO0a0325beOdNL/AO4fRBHHuU9TQMvCOPwnC6id445M
/6RTYP11y/7wd37MrXfKT8pZTMip57FP9xCncBPtKE7kGRqkJ01L0MD7iMCG
R2XfrBjOxD/uJoPzk7lkVWY0o7YWtWqNveVsbKKMjb4/L5WpO3j8+mKt+2W2
eT6dw2QvXNqjjNTIzG6qTTvz4y6/b7s177hG+Nqydq69lfnl/xma5FtdbofN
YD3uwWrFRc1bpfM3C39Fqu1Ji8KYotm9Od8qQHKnkmJmoiCz0tCxwwku2aAk
y/2KedNfYB032Jn83DKUR6BkkoL3eatCfKnA2xJ24EyUJbCtUyOYUyg+tImp
kSmccMTc38yY+D01qFDrs3l75m8YohTBCzEcHAWAHZLF/g+JKZ8LScrESpGw
Bv+g0wDRgzQBH9hpy/iFOh1Q6r1j/HvEP2veprtiG/C1r9RNAggJ+r8n3D9g
TN+1/nJHZ+GtEU8Xf1AisFWrE4FAJgW+90beZQK4jMrH1/hCqyt0qpLLfw3v
DFwXdz1DxeyqXPsyG68X38Pas0K4XqUD1NBkoF3N1ijAsUdWNlwgNkrOIVbb
Hew9yDVB5Kt7DZGFjm3Fd3ydBzwccnE/WEjncjlCu9RJbhlzalxJGWWGJ7B8
L57cG8ejafVh7XNeFh07Z1jE+h1ALhaAM+DuZvn0Z2Ttz/4cpE4FFtHDb+iU
1GR8gr1Hga3ywZR392FddRVHUV2c2q72k1NzC5fAsLsxqMFErdYZ9JnReRhB
lpYW9m1cPAj0tjrRKbs6DTdDRfKHCbJp2Xzs1gF6eaYh/+PWN2+B1P5aNM+k
eqlLP790Im1oJLojiT7yEPbXpI3fknaU8HIndThBtwVSvteVQ32Rtor+Uo0W
agN9ypGMg+pBb9Y37Zx5YT/zbJGABHFZT3pkywdOmwSmO9yQ3U2QyiBcfQQv
aRC+2JMsnq5h1i1gp+MDqySsJrc4UYUlnMjlgMxkSreWkjqwqDmevJOsS+5v
yJ+pE+4xqetqS9YGF0NeJ3Lu9r7E2ZaRyfjku7GG7Fbgak8qrcovG05updoQ
yQlgEn/lh1nUgeyU8oh0saOgQIxwFkToKAIdx+YMvD4nIlcny3ir7VOCpHek
wT2RInVBZPY+wamtgzZ3WqaBEx6yjVJ4ClbYxiUttaAYyeGFZ3IB9JjC9M1i
qbXkd9dEIb3AhNI0mgJjpK2e7zRtny1OKXLrxMCHdeh95i6ftW90WXF1weXh
EzzJJGgSX8RPczjPC3ATNgNE+Rm/KUluwFgJFsAEiDEAOxYcFnI0i9XN/d/z
ARmO3E798ZkO2RWDIp5T4Wl9TeCqOFic8dJfLRa2khECJmSTJbpuuzE8NCU7
K65HpS6hWTOgKzKbmkPys/UDzE3NTnnn3mrfmXzrDuQpYJE4V5n3Bi+UJLI3
VHRv0ndVn8DqOC/GjOrkJf8oP+cpo7kg1Q0XOzQmoRug3BXMNj47G8OrTqcy
de84g8F56TcpFiYzjcta7R0PDau1uepnBU8TTPB4+8laQwaksbd2/EaKjpSj
fRI7+R4upcNV4jkcxUO0XAObignypSx2YcD3M5BUBRx6BopGdQMOyJv/yJew
qR+vk/3odDON9qXb60VyllLHDj2xH6Z76Ram0ziMbe6jtPATJoofKKAEGP+z
KqTzBt0cF5IxUdYYurAT56dcOmC9E+K1ko2Ok+QYakpmSftjj5r4NMb/fOPH
DLQ+aFMnVz6ZNopVJdAjj1HN0m4rkihHnlq1TNQD0WFyl1FWyWAy6TFhNZzn
WCQTesWC3CZdu+aXmS+7sq7sl58eH8OkM6H3tfzk3hHwaMYzMVdQNPr4hY40
K8/j+aJsLus8vBLhAcvkvnkWTNxVBMl5ZtoA/BxVfktDSvvdExrZmK2Yt12/
0AkVMYsTdO8xYCg3ATbmCoz0DAj0EwqaVtwEFyqU36+aCFQi6BQAaeZsQ+7B
G7JpuwG0/88wG1cZHPoTwwIHyvcLmdO/rjGavedegf6Z4ZnwID2OXmu6cfZs
2ipKUk55sDFueoPVFFhgbl7oTVxIzwxtlukcevtfUTV+l7hzxvVIWIuerQCp
4I6cnfNpQaxmp6vbVPyXE5nqGiepDYdENkJpHT1xBYkZNuWAOgYq5rLJDH9t
tWGhk38WuoMHuNtXF+/bYAwlfQHpXpDzewtOXycKpwmTPEO0vWHmJUo+krb3
UuMSsBYoGYYoOVHO/fUMK5YdD1fYPFr33YfWKOa0mTyTpi8FBEtufQiQvyI5
fjRds8Aynv6RQ/BEXIgySMepYt7BrgvfGAYaxFobvBhLsBi0hnn5q3trhyos
/X+4CpucoxtrchJOz3nAycXDtVPNXnN3SeXAVxnh1vDrMDKpOzQMXWnhhMsY
EWId7rUs/E6ijECdPHwoqY1LwEAKyJAllyi/ljzyeLmt/wrss+s4hbaG11u4
Hsu6AX9nMmUc9FaAI9act7vGIwE8edRw9hd0nt+eckcNU5Ej1URtFjUjInD7
i/E/uXrBV0aKW+w/pSQG1wrWxtmAywVy4BMIiScQcLw4txc+gJ25Obwx1SD0
oXv4vyeAlY0xIZ8F3y7Q4k0TN1/FDcVVo9yXtIo4wwxSR1N+QzXWhPgBoNGx
kMPguuz0xhCB+8b1N6w3EdDag7BtDJFFwoYBBl71HcTpOZhn6/UezV6DbOIS
kh6EQrhXOy/cmuNEU4z94t8hCEyFlPmjQqzq/a3TP51mNhwB2fcN12O2s0DY
xpX6EVDwgczaxTbMqn2XbHiKls66j2zIdDwOViXgDAkFv0EkjuXmihuIpyDk
uPFyFIV286lXR9JNT2nOMjalRr8SU2OuqZ3G8c3Ya/d3x4DECDCrUwbtZi2m
mwFngNabilRVnNAUlmIvFByXg/ymxfeaLCilrNq9bb/wAtz62OIUMxOD4/sk
i01PF/DLAYw4WjkkZua16C0OYOJHdpIwPPa/sjGEQgdtCdmCXi3pGmmTlzt+
sDWCnciIScTHZjGhLHIiMjGYClPu2h+sdUxP9Tm7GYXttAFWLFPB980rtD3R
nk6HI4BBQNnK7bWX3UStH54Ew8YKKh/ZL+3nOE+vY8itpmiJXzmSkEAm0a8j
e6TB+ZOIUgzJZFHf/zGTCLOCSkycyEQ8+YTMKw0UATUO8eLSEKo/JHOfb5sw
jS3HlDRdsHMY0BQ07koamrpv0/AaVOR1L2F2UDpBzgKnTukiQPHQ5d6ys0+5
a5baeEnYad257thiNCG+Wtl+FaesCyDzjQ1BAmkCUQBvS6umf4OEMerRp8//
tKZxJz7bCnekIC1WGTBsZ4nZ3D5kaQJIMQXg3UZ7Rp9zd4NPAuEmkZPGJLRZ
/bE3KLRX66MmBIyn8UKl2d/phoP02m74XHCY56l76Vkff1h7mo0AV4KcXJKJ
NehXcu4GiqQLxe/vuFdnTjufythw5s4CDvOvecq3J+B9tujOjpZ2d+oeeSlY
41Kc766UMu/zH1Z2E5PkUO/p7LXNTaAl9psO/99tFWAQjOjhYKHOhm/PmrqX
HuWVuUaGvd1Z3X+jP+8Pl9TFU01FJ6VD2yhIKa86qnz2qTVVNdz56UFy+1Oz
LB/D0ZSCVHMDXJOSYdFR+2y4TQ7bViiAnGfSttO1Tmud7cCzcYgFAVPnhaT5
DyS3cruyAwZTkrno8IY8zOVK/zVWn5TWCttYu9GogtiXmQX9Jg1nzH7xBk2k
RD+svJ5uUXFNIN5T+cnIOGChYPPegZrXuEl0ku7drmhEbF7Mp4xdb7hTBJTY
+719aX39ds2AodY32t0U6o6IUcM3KkOwesFJSoWaOa1qmAYf0gyDqoBbW6XN
JcDC2YpYT32jNARKYdkeZ98qRhqZPv9nOEaqZdXbvKibfgfRyl2OuTPWlE/O
Y+LfAJdTFRB/CcYkPtDsZYm33FPmTLWFc9Gf47uglA4iGIPiF+lLk4is8KgO
oIefSIJ1zE+7FoUhpRtWBRITwyxhQZ/UxJ9YdcxVESelp4om/xe+Py3ZNaki
1yWZTehyGI0FGRimrGzvOCGIhUnAcinsSm5wVseb+ffNnHC/Gk9ba5duwzPq
FkceDkREDCyw06Yv+Ywfti84QrqugBPqoIIsMnl6m/dAwVSoLMkG/zi6vdnK
vaiLG1Bll7twUoFL+kJM5VfPOOO7m9R+O1ZNWPng9mDXCgSTxEdgxTk1V0b/
9Wb7SEofA7NDpQ3eH+ykY5wcOXrhiYFdm1Dibea6mXur07nefpBmDGDTxs5z
9I04ib0jj5rDdMFjjZE+ucXnpHfW84rQ4wBlt1zkvOS6xwEWfkUsaGQSi8wD
aABi1yg4rNvuJUTwNirH2RxpSlL4RTgFpk0RmA8Nk9Hf1AL1zhkv9Is5I9rZ
XJINKwLL66iiDpyCkgwekwfKji/TLaZrM60F9JBp5ZQnfPoJWu76q48l1tio
cUOO00aGYI72XNQLgvsxVz7MgWRF1KeLNYq44iCIm53oc6KkcwqXp4gRAiDl
OLbZAHHsqxDnqsIuLStAllk+d3loKAefIElctBxQxZ4rtqHJPxGUjLxgPvSL
mX95pJaUDBp43132OXRwKhEjm5ih1ND+5u6iMwte7Hjylv7Svs0Rs6duWL/F
qWEeR2azujBPcdQRlrqB4dQdlUYc0H+iODsQ+WhOOQ/EW3aJmAt/oOolodkR
b/nBd/TSGfVlSHKdKmreQ8RlesNI3I8PWdoh/xjY580o5GSrD/m0d2VqQ/hD
mqFPobTz5KC5vWoJlEIR75bowx6U9Bjq9FifJvg1d3B6YKrO50HwO+COf9di
Q+k/N3SlgWJvzZUDBBKWil/qQtCdf7DnS89y+qGF/t8plX52Ag8O/Q41sJn3
lxeccqUG7tcVsiL26hbvinml42epFwV0ig/Bo4ipKjrtbcN+d4u9f3VK/sf3
1e2clTI0YyAkxtkbBTNfXb2Z9kF1qUiu3UeTsposxj5vh6HI1CWIe/zf7si4
A9jkDwTSb3p+LkUdAJGKJsdl0A+j1YCaPILt1xIGl+1wZpu0/cSZmF+Ywia9
U7C3CptYSk31rhTmlAnrYSXVnU9twhAxWJqt+FO1uXYayduV4NauJsuCjNZp
8ibFUwZsBqk/NR8U1YY78zZslmBT6yi7/CPQyN6cmnqzR6FWw9sZu5yqudpI
qHaWGCZMni17yKYxlTUN8ZTBukxEB+TNXZdg30ogVr7Ad0P2nEgTen7jAhoH
atGHCmLIlczRKSfmIZySnv999NUCnBJIQN4YHgi4cu0caS4FYVxEFvmKQCmG
sHgkmEPiXKqwoX9KDwaBPPbaqnFpwydFZ6hpdIQYRVSqUscKSBLGEXCEMbS3
b8sx6yCZqWXu8rNz+fkPPkEwLVT/zzom8SikW6l4urX+ThahfhKSIt9E2wJw
H72Z7uuiWTs0AejE5BoMRc24r/D7c9myMjov6ZGOTC+x+kK5ynQm13TxNh1Q
elef7c/5xxNiZAh8YL810oihQUmkzGHUxSPa4U906xGOANMggk6qCaqgnZkY
c1WlTWtmHFdjKwXm9kxEgY1B4Wca+MtRngq62HofFjMB0uByEjCtQQom3VD7
bYkq+N8IOg02P9thmV326BulBoopnQUuRgpzREYKA0yPMwhGOpJSTAqgo3Z7
JOv/s2ER5mPjpE7UbmfLW0pVHM1NWoQYFjVGpSm0DUWtebVM7M1/okoiWsgW
RIEj2R2jrCPSb1jRtmlKvNhDvWupuNiCgLVzLhyQouJkTSMXJBeEzenj2Ccw
+5f6v6Gz91wk3/wEM1yuPwX/LOo5cagwZoBZvw+CY1zFlsvaRabAMtq4agAs
Vm3l1zttJP1dg/XnvgGfOou9B8uQMpMpeC/ZDPEKGHhhILSxdonzcpGjyvjE
LKLpSWoIG25m9jqPTGRakzn1lEkOD2+DNqCb/f0SkTwso8lGrGXmCgvF1hfG
hvThUjmvEKXJwWsZNrEoLQ3NXEPnlOAx/jyl/p2JolepMAKnliJ7z+bVgmp8
I0vnyguoJYoKdIAdjfMH0is6BPiNODwOLILhSB4w4DvpcMf4Ot3EMllXzuPE
t2qSU5lgyAYkkpTc/Q7e1mM9SUCoL0dozIjiVg4l0jjGGMh3IdM+L2I34G//
wfWruNrXepy4YhvoVFU5NZHHmo3Zk5YpxJAspEO1Un0KkbnxmdFUc4a1LSTX
GVWp2gjxmFgdZTe8/b3sZjHShPhPxGcG/OiUTXJDpEX2dzgUfqMYJi3Ebl35
ZQXSUJVWn77nb4kFuIjrHzRsim8oZQEIdIzevxY2Goeho8faAqc89btUiP+3
STbwZ9v6q7xpD712pzObMpnd1Sfu+uT5aO8lrG4BpR0SHTrJvmSnS+ge8A3W
rR/TIlkugUgPlaMH7Cacp3LT9vfbfRyLpSNAcuWoT8IbzJmfNeUIAO830jiG
RDPMt/wr/yd2yWw1cjnINPKEY+qJ81tT7qZhAxOlfYM8FNem+cwMYKd/rl+2
i65+Ky80CsMfNPxRnv0gAqdtiq6pbmRFWWqvf/P1Hda5mdozskMBGSZYwXrF
p3f0QCK3fTvCB75YEn46l+GDRS0q/JWijWVeNBtJ55IZddxMW6XwpOTE67aA
EVMKKNVLPE332R5XhdPa6en5YHycex+4r6S5Ia71gsuto3V2shVxKYhaGzm4
w82d997iIwEykWaYFCXhqrWgsd8L+yCi9tAl9wsQi5SpAisDUfH1A4biDXJD
0h/PYGQMJiFpRcK8sCAUTzcl6qZ4u0+BRMnsjk4yokfJhOY28SWnzZLgiIaK
Fg1qZZv7u9syZ+V42FJZZ0sKnlQi0dAW0Aujua/4BgMJpGkIM2iRuzqJ9SJT
dwT6MXvrMarjYomasxhHgH0jsrwStlYyee3W3KNXI1O1gbqRhoos+cHdTajg
5fwgXbtxU0LARr7A5ZeXSnunuTgB7AlfnNMEnIv7bq0vMtpsj9aqrUsYG2sK
Atg8VvosnYm9cVcaBitUnAR4bDoNRsi3LnxHOS9Vwp8gx0eBV/kpWC+8jf0y
ix7fmY70TLeCSLoNgigt7v8ljgLP06QR8inxvAL5fqaFZbdrMu2C49/5WzC/
SKBEVMBYEDVLRAUejYpw0GBv010e1cwngaYZBJP48m3XEkBPWW1vY2Z2gwho
rwo60ivxDFwAxMrREGL5cIRbqhscPw8hjhkZsgLwTC+37Z3vELQrstaEmA6a
32nHJuviKqbne2VqlPy/IPg6VazUAWVHYz8EK0oRCZTKmTFGMZBxUP6UCwog
9jMCvETvF0hLzr3mE/P15p6tIoM7DDhAS2IQQy2IdVpdzjs5Kzv9lsH7Zpbf
6z2zGG4BdSv2pMwwJSKWELpthrCh8KK2JoaHBLxcXgrurY5G0m+BV9HaXq/J
lx1bimLV/ABBVymSPS/0xy6cX0eW+ciP9b5Y2KyxIdMxiWBkXJSYw8atAtc/
/dMfV5oLaXmej9oTqtsslIL6MGpO2Td2sOnfpJIejm7FEb6BMkMuX7yFxQAz
1V1NtfAdglVgs5cyKkGmXAqNQu/sI17i9UuabRxLUZ08GbqXtW8sV/g66Fil
WZcsfydn9HRXKNsJ6r1qG+hJ/HH+rb0k1nFkfhaeIDWNYArYPzkK7T5w7zgw
+SJKWpBFzGRMH9l81KPFEtoVLV/fghUnOrdYv5FqPXBCu463seVDbsjrtkiX
fXtSHOTSCtCYJReBM8GAtAA9Jh/RbPZYtiiFHaR5E+KIO72vSWl3P33Qwsiq
m2wEZGV5diNmSdhp60ZRbNcvpczb5RZUDqRa6jreBN3oCwKeVRd/lmukl/w4
z/A8Ei9cdNsR4nCgkNwDlylwEeJHkqzOStPbzdT+eKmSE5ML58hp8LumltLh
ed/XqICP5+6cRXya9hZH3tMmV6Nr+lXBHVjXM7Si89MmhxQXdNtOS4pKNiLl
RTr1G6FzS4CYPWqMtnOl366GkskTDd1IgXqwZQ29qgYYlSnBFNw7O6MpN7ck
bZ1eruWpN/gwTovnhQo4+X8v841EFCSz7QWFK1YnDNzLjmp+UghzmHykSIBz
HcDWUhoXYauG6fu63EElgKIQCpHwnSJslGjAgNiTW+srM1qZUPAPP2k7cqrI
yvE1zZReRQXtCdJf5bTmpBTBaNdQSf5B6xB3VPrsBSycNNljw29Trw6moups
nLmDuTEd9fmbEKJ0VWrJ/SRJiz+4Ojx8fITThvHLi6reEUasRkWMnQGp+zD1
oANEXQ5CQolwrRvzpMr1ozIB/rH8dpJfAYH4UXsbIx695n2WiSHgPbeYJSZa
urN2YftVUxqo+XrsZxl7v8q/cChVI/G0e59fpn+86vqY7GE1dexYKwhXOvfY
0/DK3vHzQo0UpstxlHz7ANH50hpz2VtZwlCqimY6Mrdmxsny2DaD/UR49BF1
GZAK1K28w+JcSW5vrqraBEercEjvbrsFPkxKxJtVX/cu8MRYvCJEkOVCDSEn
8KmFRGGktNbcxVOevxEp+XLIuGwyCQ0CJMJvr0iUgNeFbsZvH4c8AZrbyddc
84PAzlMh+ImQQrYzrlblHIdcyoyVMbfIn/oad7FHPRuGM+F1qL+NbxGr2JCe
MAqzkATBdJV/rnodZE9bjpD0P47n9exKnvIwdGDOSi813sYzsZja8YTwewUx
ScLEga0op4vNqNJHVQT4Z9dgSswR1C5rkKN2PkZMP4+DkVuFLy5TNQQ3IXTo
E0UE5pFd2/K+RIyI21I4eE5/2o8wA2cn3uupCKGwyagdF848n0puIrb34bRh
TA590t3hPHwNKk013PzuPkp1vVruzZuTDALrHvIqUzBhck6se09QtI85pF/l
q22/Xp5GJ3wrgC+YXPqXiYuBusf2+CBzcL5iQ66qq97S95sdkWsW5K98byvg
W9+/OqYfDN66CyTfW0+KO/sQtKBd0abDQPbIecjqa1+BpgsRs2OizNYJciki
iFMQCBfsRM8tktOA99sca2YGLYK1ivb6Qij6tjI0KCSpFqG1OphBF6+zFzDm
N+FDfTEfBPNTKTdiMlGkja8tTicPpk62yOx3eRUIlOcaUYiZzBCS4XV6wZNf
FrO9SeOXZqcRZmdASVcAUonZHZrjlDCotPaNxy4UuuTnIM3FgJXvpS8eqGbq
MYzx24nnrKCgX2zaJHCg5CA0RAuzmdKZweFifKeR4ExxNJH4y7uMyfYZf0ss
OA0aHIlkoFVz+ViPPnqlXCnp66IjKkqMqHOleokW2S2z0vgvbEcw07n+cNBZ
FaIb9RddLEvF6Ue/HztaGXic02e1zbaSBQY1r+Q5DVqlP/vOIR5yN+B4ZeD+
sEOlLjCQ86Xult4JDkCBX1OWCtXoxl0MofNbqiCflG6qV3jFtP3TOajZRHR2
qi72XtS9kPLLTKHqsE09xHZ9W4CbJzlSCO1OkZ8eBn6GfEVxLNYwLS/DTznT
mxFYi2BIlqd7v7phN7RXgtdIBh55ILeQZP+2s1Z45CGPungiEfzm3YWtfPiI
9rymzEUVXAU2PA0SHKLHu+XBLgVAqYELjYcmerSD4gF1hWe03yvHtIhTZRm8
45kRpDZaD4GoRBpd2Sx74W9gByt+I9KIKSaGf/aZCMua9AJhoSDcEy4NvkaF
XD7eIVCYpbjVrs6Plr3tv/AlC3yZIPNV/jlMA6Wjw+IR4iomCCVlvrBswPff
1QDFgtbeYkSHedelMgSTJ2+/IB6/rC/MmFk0G7ixsjvLG2k3Hhg3ElTVwcMy
JGnSNVm1MeHrOByra19wMgWJK7Rh4h7DFMgCBVHUPs+aVxjLcVKuNjMwcvQB
xAoz3S8D/se0fxBT1cXY4d6GmzkL/H/CZCUqmk6K/hn+Yu8DYe6DQK64BWCw
LO0qdLxXp+kprXCcPjAEp4FXX6Ief6GF2ky6FAFdQmuI9k9q6w1a6E/aQIG/
dANuKcZIDASfePQonzn9trtxi1nY6i2FXJW0mYzKLS+m6D2e+INcJUZJQPxJ
sUsiKCf4a/TrUsOJ63VQsCSEXyywzg0qMSVNaWR4eu37rQ3DjuWd+xYesoOJ
04mgvlytWDDyZ7sGprkG/yoIAhGD2QMQCpzLOYzaXYlC+wtYLRlLMWcxAYCw
Lu2xSnynpooPs3ME14ohrEm20+uMa+qqYx1Rzle1G7vEurnNv/hQh7aTAjYs
RAvr30AwCkr3ztFcxDdTZhiSwpkoJ5SkHjFWcJhWQoA2l2DBFoaKvf8EnSP1
R529KFmbOOXNkqqvpPCfiTalcjtekQ5NX/A2r/HbfLwSaC7R8ddSHxWRTq+x
M2AkcDq7Zv79JSSHWqxS+18HA+JXIf0F+th/9UJVd7/AF0bzKuahf3p8tkPQ
1hBnfnAm4I1UUmYbySamvFmKczeoDaDvenh1jnqMgsefRR/MgarxnKwYce/E
UtdjwddWxcg16LjtLGvWBf5P16hwvEXxBG+n5wS6Cpe1+xF3NFszu/mJ/dgS
7EZdvgJS2o8URhMc8SIiBSbGHCgqyUB1Ru1KZK5iT0rlrH5oCQi/BfRpBlDg
uRGrDhrwJlc17Ec/3S9tPX35up9J0kNQZmJjc8pHYreoxmQE0dABR9EhlMVR
opTBlvJ6d5dEANCj8xr8JJt4oFx7nNCtZtuecDQujJwzUMwWteduqE3l3Sl0
blVsNlARyk5PXOcD4LL7H7VTXDy7/CQZuDXirQz6P+Qr2PGGC2I7GYGQ92Wp
I+YqVaRBinqcQtuQD3cCKrLsKfGSYBV3Rj972g5cbLXcEqKJaooY1znQpYTQ
OSeJTtCbz9QUNRrp8GrO8LlKDqxXyKlW0Oub/smbcl1wEIAdoEjEFo8PSkyZ
L6V318Fd7uiea7Ki18nAWdxnHGYRhaH9wHyGov6LoO98OZ8UZX/J5YS9gPxs
os58f9d727R94nWMrA93k4yhgtMMFZ1Gwus8vEXas+Qoeh77eCoAiJhVn2Zk
/idiULH40gqgPREveg5GMTd1G82u54coBbWuMEOKRM8BwN6eWn/WlSxajOG+
QB75RZTcHU0CrYqH4rmxiO67/dGJrIzyz+yt+yoU6yiMjFIOOpjyqmotUUEJ
Y1hn6Z9RVa42O7SNYS5+H+33TdhtcRvq0uLOkLxrAIFbj91RSAc7RN0s97EM
YzQ/XEsjHNPAaCZs/xvNkn+rkd72XKkzMH6oXwfSqLTtHzfllQdH7K+urzdl
6EVr+kVLFwDoemVyjFeCka79uwwkWPT4ArMXOj1aKLFLGXy/C5r2KShETTvw
6UGWa/YDP/NAebshsWtGH2K8L2C10CG1waloMS2ErGAJ/NTlDIAgPgAMmzHR
s5PVV/z1Z/I8VEYJTVdQij5xjufng6zeoabVDdAzriPWUOyJd8nqOjySIKkL
AdhdukF4Y4BcS1Oe6hRr5OZgi1R9ol/ir1O32n9nr83dLgKfZBfzzZVM8+n1
Lz+jRM8DFWtTWjhx3fB7cNKNAPQgxLAR8qruDrJGnPIMjgKjusSJ3gW6GXZo
0MmTQEP1bnLhu14CfbUvgwYcMyFoccvsWMkGz+d9EXgvudkIUm9Opm4bxc50
Y/PHOMScA0riGiXKPJuajfoXPz0+C2JsGR2mMq37/iXgAX+IXzBMTRZowzJm
MhRJ/DB369VK22FonkNWnCLvrprVTXxsB9A3tgai6VYmecwlWCqkDA67fMpQ
9UVYg3aLbce8DAjcnPvkwW8V4Ic+LuXXoGETFV07yw9Jf4q7N73gzB6YiVfL
chPYaX6qiYkB2THe5iwth6BnmtALZeZIDEWz/JKRRub9Z8loFI1Xy7iDAKmC
kUBQhFiaq2pZp0lTWdqAghM+exBW3li8cJjmKVjcSRyyGe70tUB61nH7K5bF
9eMDbqbxvQhhy87lTMQGJMZR9sGMsnOBvzaVTioziTdWXgQiHxpMpskGrj0x
yY7CDOiQOo4ZLVfOESrOMgQVo86mDA1Mg3Vc5bpCH8dzmp7y46u09vbGtx1m
xtlZ/DLNv2W9HZUDc+uSVG2G8agUo5QFNJo03mJ+AH+ZsNu2lPRiUUdCCgfz
er0w8TrZk7XxTJ/XrTaJkk4PyVGk6ZtWB2V5emxdHioy6FFXYoGPO9Rg/b1V
YoYwKsj76etjseQ+esHV3cInwfx73kTwSl5AtRXjgeHwWPs4FDclWhTyqhf0
XWfm5ZT8DBzlG5VyeCaWGMxhMAkTU7o5LdA/o9P5woLzSkXUrBNqFt2HuN+I
J5C7U+Pk4iqZL7nvZDoZEvcvU6iBM9s6CT+tw1uCiHjz5lwzst47lTydjme2
YIsWbEOqrFC8affYuj+5dBzssV2ea7jPJtsiA9nmtpCstOHeacHFLHfBcB0I
y3hJ5HZojF/m36R3u/dFQ4M7a9YiKgI6SzIZfpIZUHCSTKh3DKbbsztFHU82
B6VX7bijnRLjusx8yalQWxVNAPFhXmFT4ct/G8x/mmkdWpvF0er202uhD3nO
3ida+AUglu1bMugvsW83wQDpK1QeGhjCxC702CkL0EQTlxp0gT0/9UfC7T67
ifZJ1NY6xQ0lS/OpSSyQ5QsKvoCGLDJjbrmxER95Xj2sdtLR93wAVSQIpCul
odWsZ9TK/tAu4ZdJ99bTTDNaisP+iUYGf9cx8TW8lLKPVo3XD4vsfCqPI0mb
n4VpC+3iy05fOugy/dAewcCtVm7tOpR46//8+jGa0ovttCjE29XZ9h2S8tu0
1YPSXvxgXKv7EYmImTKBOYXM9LOh9M3S1/h/uYQN0a8WzEwT2gkgzKClZMRJ
CVmmO7EiUPNiT5p8R5Iu+i+nQIkj6FS3j/3h1CnfRdWe0qBBOc2ipgYY3FAP
C6uAUWiWmF1TQ7+zj3z4GOeG3KuMfbFP50R/LR65cUVGrAxhVocfZE0ouwho
FK7AIJs+laAs9qq4o46WuJPTGVe6ATmz5BEzEUPzi5nR2iGWTawJ5lYdicaV
8yjdqgelVFwgmeBDy0nR1bV+tOfWGHkm6AfysHdYVwjjpODtUR/aglpDH0Pz
aBNgzHgpEso13s6gUolRCvObvGeTkHoodwLDubE2H5LuxAhrKE799MAJ5fX9
P5S/y+l9Jri1nqO2dT5+1QjSwkWGjNYehRUf8nK0We6OJ12J41Nve1D1Q1hd
t5Bd3yp9VvTywNBajYNi4dGjG93FQBWrNNpJvJJ+T1AM1smZwxbCedCjlG3W
dxptUt8mlkAU1HPd/qtkQKN7/CyA1vVjs+W7tVa7WjDAa90E83YEDVvRs1F5
ix2HQW1NjW3cyE7amanBo5n3or7Z8F4L2856obmTkiy0/c5Nvg10pj0nWGFT
CfKEqeF7rZRfZJjNecYp2XAoMSP3nM09JE/fqu+mwUIqFxYxsinANND93EbX
Nr866uVFYXOyN7puvU9dqCcbkgEBvpTJzRPli9xYNzz5mTQUj4t96RZg8/nS
xclhc+19wN5ZEgMXwzMW85dyj5OCbIz0rHeBddokiQg0+fAQkSqzutlJce0H
u5GA1wo8lWRr/koDvrXOokC41z8cVQaICRR+k20iwDS7xx/OIkohZEzzchER
3JO0LrzU6v0T2jTeKUESVimkBMaYlfA9tdFBi7gfB6hS1eueYSzPInX9vjhY
kbFP1rvXl4y4Lhmi1u/znbnlslmuUr7W4XeCPQQgyI/63MdhVuU/tfYh9Lsy
yp3xDC9oxOs+CBZfPS4t9h06yzHIvHKSgQBbtsE/NKelA1WQWIQ1BrEKqL73
umm3/8AmvKw/bCi+KAYJuAhO78lO8+hQ2Rh+UtrmjVv26SChZhuGcEn4fnrB
Bgj9LmDJGwsECvAofc5O1Z8f4PXiVJINtNYjOMwFtES5J6GC7Vc+nLZJZnaH
Gvr2wHCWkJhgyrLvnGhkrVyM+SMbB4B53dwzFusB3b+juZJtCIqUCnl3AR5w
4q9nfteGHQDw750Wz+NOfLTjcU0wLFWHsxLy1vV3KPNMG1FCEE/S+AFrrUNV
SLM+L8MizZ0868r6rHUlxP2cNci3aiZnCLquVmZV+fJi4EEEcnh57Td0qTnQ
aKjRj+rLrrSTRoP78fELi4r+WSIzSWi4YQbLIJgaf/G+Hfv147x3ILdVvei0
Zq1sLjoaFqOspHSq4jq1pBc171MEiNXCZcq9aQb2iZzrD9n1G0QZ4PKIcge3
pdG3gfzMSG5tFiIsXTSTtvcdWwL7YL9+4DhKEXbFKQRlKT0C7DSyjup1nCRo
zqh+mcTHpQ+/TZSEiXo08aQKk0hpCFvumZSmvi9J1axS10GTM5CO3nc/xHZL
0pyGCFHM/9wgEPQSeGELByI0xNxyF1DvqPqlwbOm9G4vNSN3HKMv9+rHKoQ6
zeiTzh8DgBuGUARiCk4K25HzbUxFcNJjvaYQ9GxgHBFRuQdg4o6pGAdiNagN
86zRQ3w7EJSuAP0SrHsAWCfv+ICwyN3CrgV3ZlGWKClPA7T+VO4xBvCrO1ab
N5qcd6YmdZsw1YlZi9YwyO9JbsYNx6ScMZPN8pQNSlxqLy5160dABZy8QsAX
hSCP/pDL9Ihw12RwH7WHYAPcwsGkEwKd9G+4GAS8GflgsPXN+kVa9AqxIDW5
wGNLw3aYq2JrA3btt+iLei3vwd1TdlHqXzTTaqJTzLmjh3q6PK7FfA6yT0hv
polNzLfDp13i91nN1uwr8cW0N5mAHCNEc8ReBIUk4uc0/+At5WtFSZ6O+hi7
0oE9KLENpQF/Z91wukVfiDFtvM/QEc7KSe6ZAIWGD0jl0hFDTkBbMLXY5mki
HjCjuXrI2a01ANd3Y9ppLYKlEnoCF9vN8wlElf9kG+OyVsQOeBSMYrKn0j6d
WNljvHWARPwM87UEPbKrSGg0hg8qMkYhfsCJM5gzlhnSGiEjkX7a7WeeyVDJ
mrS5PAu7uGKHGpX7g4hBJukJHP5r/hCGDizwOuOvY8SHFQc8CtrQxotmLtlA
7Yz5VMz/LK+EXHww4t6emC4cFBTTlmrQCeoEIrfXLIPjd4yTnRKM9NgL9AOI
TSl+xzNDrf2l66FMNta/YnyVmu6LUY6R79QxOAAVEvxYsKiOKOo2RrOHz5wa
OAq5B7j5hhoAspxxOVKfFXz1zk0m/Maye3Q4Yp3C1LqX4CIJeav7hmJHplBV
vsgwPkOTvY1WN+INeeXBl5Lq1An+XKxOUiHCDAJP6bc95zpjEj37zSVKK3Yg
FlAUI0EOFylgKLgDtRUAO8t/aXRbKQgiVo7zTaSKwaV+dxminn6yXTDduAA1
pFxxHDzI1Xdlen8NgtQ9VUb6oM/UlKVI9WXny3JVlO7xXDTblyApfgC5lX9K
mveBgT2D5+uxKK6aUsbK2+gckFE/2UlWommdohKZLFgUGCj+AGpH1E1yzViH
RSEV6zjcNz7aM9IIRHihFn5TNVSZlcift17hfBS4/qwmCkb2SrAtMihE/hfy
EWADPSj2n94MHkKgltDBUH8SV/+72ANRsTZcNWhajRxntk7UIGglBwUN2a/k
c8+by7sIlG0xDDMKMKRHjT0azIWh7s/5Qcn1XcMJHymI/hB56AQCpl7727W6
b1fnkawzJGnu0lnfzMuJkOkMRPVVtMfSv8HAPBVz+Bfvj9LLV73P2qaksAxx
c+NX6S4h5xfN+392M8TliDWQHCSQpgY6EGWWzvHss3iDcxXs7dKew+XIOePz
nlylwOJNDC5vrzl2otnZBwi02eVb1I2m0jqvgLpPRZY0SERh56/1fZliH5pe
4YbTKk50zCpx6JL8hRrOb722lfT3wOTAHwkgB9ssDqqURygogsSPeOnjM9Ll
L4YJ3I+gqeNEYbyFdweT4Yx0cIDK+7/aSK3zNqcn1yFZ6qj+Ui/tBWhPI6oQ
X6DpHv71nf50138KI59KlM6RM+D4KBWW5D6rdkGdXUGSLUWG6nso3M3KSljT
t9EGxxVn6QKKFub0/ns/1/l7ETgsXXvwKEnurogmGrIR2IlHg67AVeWX1NYI
TMpXGBaoSKnNYVBT8kzFtRdmPXnXNiPg0VH09BhXHSv1Jg8vNgxcDi56UoWz
enDczn3evAFAbB+uQHYWHJbqA8byTIxByD9/LudPVIT6jUZhTvMKmx6iNvlu
UaEtT1Fer7Ax/bzjw8bArcXF3rBXviSacMu/+++E7lmio0RZdm29GB1vBLPK
V2IE2/J96372pBij10aJ2hMKdbls/zIS3VnhD0hEkJoIdwb2EbA85zByx5cR
+HrW2xHR2g5fBNNtQagZ8sl0Jrlco0a//4Sb2CbnASgB0kJ8bUeEjh1tMwND
RFAnBpHSReHhC6gg15Mzz8yc5Q9Crg7+lf70jRY00k0fBLllx1zZE9REbJTI
hEnKhbf+QRMfHGf2OK5L95VyWxcOLJxhzTGVzkqxxypfduZyUL3cfWWGdhol
nnp++/h+NvhL3Zni5+rFJhoW440NngXBzWPTvhAah7VfvHt7akZyxkMAY7pY
IN5vxnrbjqeto+0d+x3K/OpJP9rxfNSDL6zwfQbMkUiRPj18QwoEGVFOZoyA
JjUDcX42dkXWMN8UU9FetQA22grSl7Iog1fm4WicW9ifZqDf2VQ29ZwnZr7h
diy3Hs/5hhDpZZ7hLrpLIctLKK+jmAiu8Bhkz4sm8m6LfCMZHqurWCF55+p/
Z8kNy8HLgTFQpIlA5zeN+p2gSlmx5t6Lu+0o2U1bUL7vshV1Dseljel1lOCw
KNqcvPq7sMq9qBBrdh4jCRVMInRYi6I088bxG4dib0MgBxAuYLlOHVkmVdmz
18UOICZmApIn1gyHLNTEAGndZt95fLeSSXZEXLISAtntTdG5iCGshdS+sLe8
90JGscWgaofOmqlQAYS1uirHr787D3UXucKe5qTtvKsAYn2ClTu1QtKVUctn
vr7Fwu3ImGPfxibhvnBnsZzKvRp/Ch54vES8NhZgMDwuQ8En8jVdQyd2zhl4
A6q5czCUFT+ZOgsQ9fTXfsstfHIqigKOAeP2nLpe3oJfAv4ipbZZQsXZ8vZm
bD4YJd3EJkM8EvoTSOFU2vgJ6sBurd+Q6Ztp84ZVIxwgJCuj4AEyBSerQZPO
XGYqjg93VMOtMie9TkTPYoM52NDbxYYOBlWjo8Dt3/gjfbDkKEiwvHdqKGeE
ew1yZ1Gsx3d1zRvwnoAzVTvO/HoHqOjVbo7Cz8OAYjPpyz5+CglpDdRFb67T
AhzggcC1I693a1eRgSeNhVRjBhkw/thSDA+6Sp+SW5eUVhLqVvxQ97dd87li
pu2GqTuElSMB/cQSKcek05G2ovrmnf+4q+xelydJPzA84+znaJtNCTGPZ9Uw
bSUKxFDVv0SkDGypUn3pTKMBBCPYcKyISCBkQjvYBLwzCW2IRQQrDD2jFUc0
iA1Ee2JaOkDAZkYHFMptRpSWhHoXvxhpvp7ppEju9Sk381sOnRxgZvWRwglp
/o3q7EzAGcEMLCsQATexTr31KeqgLR6sgCazRD4Z5rnxlgVOLTuG/j0UIeTB
EcUdW4fo8SUx4etUxvwGE+R79SXYKKjJHk9goPhmiR7z0+JMRSIBY7GQV0eQ
sFR8SuiwNsuPgYZcpzbHye+c9eNvsImdStFdRXAgNeSgGr5xYkEJhF5Cm9Gh
NMJ49A+YAwiJflBmh/EZafJdNERUANX8nAcS7c1jseaqJgbeSSAwfDcQCYWy
nwQl6JDP1Ao9NYBurwljVpsuETCtkzvOVgEK9V5LFfgXRQtnyaobFEEUK5Np
phSNoRRuxKf+hFK75XeqN6EYlVXhR/UfASDQDD8TDUr+Nq9Vv1B3rL0iek6B
wNZrzW7dk5sPLgrFGEKtYUKo/HiAe6HOxz9W2kRcB8VXFvjgRCZLfmmGEF7s
zGV4mGgztQ3udl2e6QNDajDFl4ctM4ag3e4UXYQjnQ00ISNpJGqSARwne9CP
TZ41e1FGA8/rnZP2Dc+1EUV/Ze9DTj3TJ8nuo2ClhDYwc9RnOoGMC2clqauv
2oo+fxTwk+Hv0liV6VCF9JimEkntYR1lsgSMQ+5Kw9zjhI/XqJw80bxIDND8
keuZt783uVb9pLferzN6JGukW8Hk51eF1MPRa7Bu8AME3QTUFRtAgtCqfZ2J
Jm78qpTu3Uy0C2TEwtNgKyG8FC609bQPXStyp6DpNmWrOho6H6km5Mpq/QYh
vY5vTydnafcCgGEso6MF+xvAu8CdULrW4v3mOhjqUHuujdfhas16tMrObB+d
maksWbty6FuIx6XBNKmM1bF9ssvySPqbpa2xE0Le0iEkFt7aTiFQTjSHS5Ys
qsTcKzAO6JGkpdoEpF2NZsuBSYZeEtqH/meIz5iggb8462rold74rz2VKbiL
/MEkT8P1IJ7gVo02ua/4B30pWgOKz5Ntbwuie7P/VRFgrlPqTe8ZP7NPZAzT
iofrtQUh7R8ivCj4LFzocoJzwvmmHTSMlxCwXMKWm6rjH4VOGXve+hZ0h3Ty
l68UXktWEIdQIA+SFcRbpAvAPb4AFb8uB3xsb+R/UlPgoFhXM0r12Cl8t7Jw
3J8Fe91O7bYUBjpfOBDCEwfh1qpHFfHR8pZHtPHK+U5V52/rk/6LOu05zDQR
WcGLQWq2/+PuXDIBilgj11PTBg+I73Q2Ah5MX7TfmJh/UedHrosCPr25w75r
R4t8KDaxcVJMk/kFHk5wVlKuwmSqu3WteOaXWmAzj51dKjj3zjnyperL0Juq
tYRtH7qza9HiRWChEKr26Dnm6PucXfQae8rxaPe+n4oczvZowMdwClnkKQBU
1eO9sGLP+fperBfWdEKi7ZTsps2+GyLZQFu8CiBKh9VTtpuhFcNd+Rn8NvKt
zAe7Nb7xNKq/dGmXNXzZjwwN9d15d9QuQZiKKOAN3pys/lFU05h3hxzMdZH6
IwXvdQv1Nx7DxYaWTGu223YkEZx17rVFSyTPmjH8/BypVd9Tq+nRrm+ztjGC
zS4dWSBF63hbsWYzcOHXaFkFtCllu8lZOBavnxvrGYA2fXo3Ikqqj2PQjg30
RHeVnu6dGeBG6UKI0iK2w/wATKD6lrUcPU5/88RWLIpP78afApL2t+NbE+6r
ujcHgKG+zBSeUt+iCZ9UHreFCUVN2jTxu2HQEN/bcfxP46MVNwrWMjaDPeIb
a6fj6pE9N7nzuYcTlorTZADAJ7oc7NX7glDM8DKWRjkbOrbvfexFZwJL5shv
bS97bvJcudR5uU5zmb5Bvq3Fb7YzYONjdXVDUo0R9fPTxh4dyw35XBMJjeq+
CTj2L3eAScx28W8OxlQpImRurMKmO5MPXlgiKpW4zzHQhU2c//strPq3nhVo
W2QntYSKg/knFHSwaoZC32oqHDsW7PsWwstCnJqcpdDCt7ddQO9eCiO4/Ahw
ayR7DREZHTwTUywFg5PGusQkAGdb8DKj9I3G4hrCwBAheTYivw1rKTbiRCRZ
Pi24GHgRdPpMdExdDAL1QPFMMqV/irPyRb1tDED12a1P4VRON4gklSPpWNxR
ufq2vimI13LQlfjhDauq/VYPZq5GC6iucUvSScL7VZ8y9gTIyUMsq0CX6TU2
yRHj6WmG5kkY60Lh8H/MGZ31U4AJLgWJKaitGrkHGfWsBje95JU9JzWX9AVr
N9AhkjSHKAB/Z5lI+CRPASMwnlc7Tyag2R5k5UfTDHBYbLSZgbxnkyaYiS97
QuVDt1+OPbJIjE+i4xCvIVaI0GuOLH7kUUVk9booeCSNOV1oIBftA+aK3Rp+
qzoU0EYRsg59WGVMjtP8x9kI98fAPoF1ombfqlcS8LWYqQwCko68PWFV3AMa
7WpkdpoO2+7XW64fQpFFJeE79Sfu9mkmgnlWWdNstxHg2iUsSSzD8iKRTNxd
0M8zgs79M71hOMC92Jzn+FNmlj3dkFAoSmoGr9WmQYb0UAjLcHAzzNBVWRLN
xCtbbJ1VQLRfUlQHuPm9h7+wx5JMG1PAQM05zqHsWHfW5aFpw0oU3RTCzItF
1o4iM3Kw21dt9JnRx2L0zxTVEM5erv9tolB8Q/xRuyprH7cHf7+tmEv57CKt
popFg/Y1LbAN98Lclmqe1r51jDttlB1mtyzK7Cv9MbgPxr53bC0vJ+RyJ7Cs
ynwlwAydyI5PKg9rNE4N/AfqrrOz8ZI1mvS5FD4Zc4y4/Br2vO7DdT3XABgM
mbW8rhR5mqPySHdvLSUipcJMVawGsnyTruxkL4FUAhtTyv16EoMaCM6Uh3mc
3g5shWBtk4iL8BtsMikKvZHXbdfneDWvuVZ5XW0NiKBVcsIa+MtW/61Fq2b9
UjVGG+WfQPD14x+cBUfGS0BjX3RnDUfzASKAtRADMOfXkSyD12FU54NKg9Mn
GcRK4F+1gpFwFtqxXKeEIbxitmf4u3syfDHQcAz+w0I2XYv7ny7Q0Q7TZlnp
gTZjpZ73R5BXOyvsZA18FX03VQ58qXP/Ts3Vy8ztYcHbrOYsNvT1Nmx/hFs0
uaDaJVOWNCRdCNvtS+PviKNR3XOyB9zl+ZrHUREfGczTBgibAp4U8gF+ThpH
rR7csW9U5YmjnzdF9xdEqW/YjVcxCIH/BVYx+3zqtsF5itG8o6vMAwiCWEQ8
diPnFYzxMzQGWmMXkC8qDKics8claItt/WJc+sudHOPfyesCp44Luudb+5gz
DWvu53CPGf7H29lCLrmTiiELt7eAkrAogXZ16wwwsD+xdK2cv5/qLflmzJvo
CLo5DTV5RNQMCfIhqxaqZNgwQ3TwPr4eL64fLXavHY43NXh6I8GBvLObjABy
YWPchnNjZM0KPzjgf7b0PFkHUDtITSvs3WQfliHkLHBdur7twpldZzlS7Psu
mh/UEQ3U49/jRHgsBtSAJ5Gerf+9imbTuSg7wFP15cCfx6tXD32t1Fh3e+I/
ysHqct862KeyKzIsQYFCT0c7hyaE/KLFIU89oGFYSPB+b73yMk4NKffYv4LL
XQRfSpV8HZbq1eBO9PJBcpE96f9KDijBpxmnaao80+BtJKrfhpSoA6Rv7WFc
VtOgQlbR+nXcZUDjVO4OE3fUjbSPdLPRgrVXSsxVynEHNQv0Ve1qz9acebeJ
XUr2+PLyjuP6+QADnL1UFVrjAGeot3WYgk5rcY+w7i0EbjVCXCMenwPt3Vzr
kg/n3uADqw177ZarI7kXA5KQcQWfBro2i4bo49zqzCdhJDM5/3HPUUfvw0j3
foLqGWJWXaSsGclETWBiVwGt6lVNOVFknoSwouUA3uor4YwFOqs0CLya+Z9K
QcKcSNpvg5yCPsauDTgZm2h0Oq4E4RWcHjuHrPPm5greqSRgQGs892WEndsS
eTco7XFreTXurDWbUod6wWw2wGk46rtx2UCwJq54Z/yR0oGTUWcD6fnvzyjL
mYdhX4SaITCNVusirxaRsjQCj9QazaIDVwohlEiA3voCVswGqgyxr23auldt
y8oInouv6o0zVITd8Aw+PnI7DuH3cxyhCf7o5iqQn9vyGvJHtEIgLQo87QuS
dlHlhvQsVOZ4zXc+NNjfWdw1IYSmc/srClwC3eCt1PFyQUr3SV8+4jjrIVBU
zD0bqzppKJeQTDT5fZLPkFEcbuL1m6tcchRTLThkE//rcSwMGfBm1aG7pZd0
lAqCnjpIlc/UbOgjGVfCpsTZITxc0KOGaNnvyfiauR0uk2ZYCQE8d4x6/rdB
xD64lxjYLMHHfwwNJlv8sp4dTGt6id96lSwCH0bZohOfy/IO7+K2FQvkgLm9
D5stDrtmvU8VZ/wdeB+nXBPEgDgsN9bSMkY80TPrSxN0LGjgZXABXn8PCdn0
EKxyALfiuGB+OHKXNAbpt8SVXZ4OBzkrQE0X1vl3Q103sWV0odWRAk/0CcUx
JEefWW11YnKie8MPatnLTsGxE9RhNN3lL735vP1z70nl0H2gdK+OLGS7NgEe
c38Zx6hYBuXSPSx53JJJ6oX1mpkfQY5qMTWNGtYbCGAcHTXX8n0qWVgYus9Y
fJHF04A7MG09VcX0KaY8qAn6rMj0vm5yWisfLyYEeNVY2pSlE9/f6dWLrLZF
EaL0uZsVqdHdBuiuznsYIZNYhz1YbL+/x6wBZrOlwSL9m4u8v2k/CKuVCOEy
YjAnGNji3OT2Errp6H0e+RwTC49fbOyVZFeJLW8M0DDtE+Wk39hIb/UEfiFm
1cG+V8arFzKSo1y3IGxzxK50crfvp5QfNgPLGzcFW04QWB1dVhJkDTUMjzYK
9dDPyg1s0/NjgfyFJSb1ZI/xkIkub4vX8H/btwBHTHKo9K4szLle9tfWF5Lc
j79EtCXAsrH69gvFSMSMxGiMxLs2YJWGpXx9liS7N/5QYrGRxEAdjxO6sK3u
F4eqirIrBCP3wAFCAcXRE13Wtq4iTPDMEbk6lRw7GXazSlErbo8B7sTcxp8h
pgvQd9BwarnpO0XxruP2Y5eMPX/HVxSOfZWAxt5YGYSJxgl2d4ZF1RNXZHWv
eEPVOCPQg8k0rodtg4tahxku/Orj8T4+b1kHZ8uAMglo8Dj6xE7Ul2VAsfT/
d5Ap2fOo2df3P1b1bEV+z8TjjKti4FgNyvE19trYpdoCUoe8xjQAxDVzYOSc
gV31T9qRZXpAA+9aa8nicriJ4vXp85bsNqtLm4g3TmmpUGU7huyL/VdhI9h9
fLc/coObImd0tlQoV9QkErWVAPciTfeTPwpz+g5AXtIBpAFmlHhEAPFQhLaK
dKdYF2BdJzYTThu/wmlCuru1jlmcrqW8TayKXF0VngKO0YvcOktzZ0uHPkVJ
pt08kpWlAq6LGdy+B2GXr0KL7prMg7Ks0Dps9tQYTQ7XrdRDQsC9Q71aR0TS
lWFCwA0pNZYJtpqOsteobQw/QvgeutBT74sWQd1El46gXnOhGC8W48aocwZi
ROGae2HlhvjwVTtwIwsttmPqbPsXntoPsLcO+JoSDgr1VqzgpZgHriJorV++
v7h3/3XQmJwJoa9IEDYQTFmfb0OylWp0/AQ8iX1B3uCqTwLiF44oMq/GM2Sp
V6IHwgA2lvTLaV7KNgqk4U008VRHjzJipOft4MWTULopq0xoX1vGyuZXKtkw
JM02J35+mKQFfHsfkcEeWx/J5VG/cFytN9Dpy3SNYqSIJXNhuu3mLKopclDr
dCG/90y5IZEeDDdm8+CCOdwstHFBKf6LO2ebpiCo5evYLdTpdmwLTb0qxR8Q
XB+XNdHmqiqHhjG+zpDjcdrSaWlS3uMTzGCtKraS9DFrsF4VlzbjpeO7lZPT
hQ78WnU56CbGP8mWLnGXG+3TWqeRL8iPqOK7M2uGmGfX7qZnTS3srivR8LFX
OER6ddR0kwKqhZ18aHYafkZanmmwBn8yiNrIINdvz1oBjt58P8CzOBhdlYIZ
55UZKbL30iXF/I4k071OL28vXkmfrT1u2wOwFibSDHeLCccSdXKdwOvU0+7Y
I8P9sYCiQoXwTFosNxq01kD2JVSbOSjNwNuPT5otHz0gY6WI8IpKp58AHsX2
iuMoBrw8MOyWvnMS3INs+NViWZcTpnPrU3l01hKmiIhgqAbYhiEdy/twwUNK
9oA4vZayBoOuPTG1hXSRotgttO1y2OGh6EdUn7iHAQMp0ZKjCamDvQcnctuC
breEZrVOT+aLrpLk/GClAnnWCxlH4CUqjqq+OB2JEKrs5tICpi8PrxyTn6hA
GG7ZqSUB9d0IfWXZEj+BxbUjjiyb+W2MY1rO74H6C5JEBxg49cw8LLUDAmND
HSW9gFNn3W0oFc8Xb5WLTIsNYF79Nrwb29QewnpyDys3fNEDIKHwaikt0frJ
GSw8bhuLW1jzvZpxxrLy4Q7f6XVIIViqSDDVs2VquS4TZb4RBuap4iayN5f6
55LKJFmG7nWIJCHF4bRrH1Iy8EfsDt4ddDcCJ8cMmGtj+8NWhwaWL8jW5Btl
RZAB3Py+jG6RxuOG1a14O73lMWoikB1xiYaJg9B2+FHQSTa14MdNC3bI8qEz
qDKX1YHMTk5sg9MR69Ui2rwcgd+BGJS6SHjDNuvREgDdhLWD4vTjKL0Dqy2o
Ny3+b+s7Obtfu90bdgVpg26eoweeIY7PWG5+7azNg5L2fxZf7QMXhgbKiEu0
tdcSzGWv0gGUfy3aFtldjU8VcDQyVOgoSemuK2o9ZKtxagz9DfIsvj1N0nBs
8iWkc6wSWIhomU3jA8pnvHU2KsEgnRHqb0dPSs11ixKPeMB1dYiAopS6it0n
/C3vG+561lSk6BEtx+xO6O3/iX1sdL2qD+kLfaH5kABU/QcqF9b0bcXAX8P7
m1wZeP+OmUA/W7AVJxtb/ocP5Fw8hT7sl/DciLMfnHxbfYVo+Nrd2wEsRoZu
8WOlYV4srZbVeCVMkMH6HjWebOR7xpdtUrvfZJm+tNZxkXP2nyWZRdttN8Lu
bvNO5YxtR967EZgNrsd3zEi2uua/4nkTB0v1d080qZhXMp7c0NKD+WiRLIzH
Hd+xCa8/Udjt8xBXwbnQL1K5reIQVGRxH3uGQLa5zptDpJzGd6eHbKPdHPf/
upTsUCqx8GRhMUyp9x47V3SgrHNQLH0AaFqkx6R0Vjz44lX773NcMLD7BdvP
Svt7lvfz/R8Tvy3GrBTAt3OhuQ+jNuFR0E9mfgyCP4IPiMUgb0SPQfr1BSfw
oCVhwFqXAkyCNTSr+El2kZxWVr0at9oDBQn421/+A8jOM3b/MbdmB5nCG5GN
sNo01gUVFIqzd76yVROamzx2CC0nR//jZUH95L3lWa66GSQYBTasPa8rmehi
JyPJwOZ5Sq5W/DzAYLazkUwV3xS/MFFeKhOoydk00Si5Eq1HIMuLOsKqCi5t
7n/31krRufs1dgbw6aBhkl3nJWzD/iwqXlbuZ4uXLpiGfHhQKmYuq7S0uRa0
WTrfN/o2En/MbBO6ctcSr8leOLxmDNzNoupbUcXcIqxVFGfR7h1mM+YacgzD
b9+M8flZw9UFrJ9zujZCletRZllHQBfrJgGi4DWDd8PDXeqxsntIqw0VG4Ho
HcU6Bv3A9aqaRN2CKSbFCfcbvj2qlNOPAD4r/ld5V4nYNMAvVhMbEN65DCze
VSvexcZ0fyvEOVHDNVx32T3FEmmfj7tUheOzndP6eqjTdrmyKk4PBVVLAnV5
WjF7oEh4xscGJ5yHrks4bA2v7NrKcZfnP72U2resOKWKeH+GvBXkJAlSBDMG
m4chafXR9IPuICm9DehoMf25K+Owbx2AiZ6xRn/lwuzxrs0rXHwlZEsDMvNT
DIbhzCWlpUF/aFW2Sjn8d0YqhcToZxgNFv+qYGMAnyyqHcFXv6t02eEYFqhE
j0vcL4Oy0PSiwPYsF5bBF4d57ocVQ+VhCMqsfk2ElYZRL6ejBcX0LHj1kVCD
OwxRoJ49BV5s5bKVTre8kFGdQ63FOjdPv0YS+QPCJ9pH9LuCgLbQ133GKsWx
hHn3nFpSElwZbglqVDHUCscA1PMlcyiOzQPHvQk007RsRGM+0XfjsDXVuFIB
MGxd2oZ+MfNAKfGOR19BQC75N3hU+soN2Dt6PmSHm5eVGTk8/4728RxwSh11
gEnec7vw4jNWeKe9ybHb/ZQ1OZGsoaYuMu4NnHe4CbPE6GwIwITqCAj9gRPN
gktJOdFWls12ksP/X9kmy1na5QsFM9uKm7iMcAputxmuvJx4bM12FsAgyEL2
pDU6dowsqEUvhxfbGvhvOWIXGo6MnJnM7Q8qc65OxTp5H1scOrDexbRntNZi
1Zwy4RIVTudFxT5aXvGZvNrXhmn//+UNJkilsLgljg6l0cssPGrHDS7ZOJ4A
ccQJc9mQ79aDEGIO/LzfoLNbpcGfPyfkEYSUbmokviEaqn1+Yf3ew37HIMVK
kc4WoSN+UfmSx8UIluJ4whF2V8sn0wPe1/5OAZqNiLAerOdmdJeHAaCg4X8n
5/I/QyD/TYG+btJsrcKr96aic59G4Puk7P9Qp4N8nemDp7lih3sLMCnLGrfe
zSL5uXA5Js55DNl0BKiDrQUyo8sIuysr1DY/iDtzwk7rw5QSVKj/L1JkdbVG
6DEw+5MO5A+jbWSp6UJ+vZyAd6ZOmcItjglNMxl9bxubo4hJi/Hy9rxM3nLI
K8rApwh95BTWzrKVX0MN0WnruxkDLs+asBqpKjKLPNwcKDHy8TWh1E1FNZCm
2j+VQxFCu0SHPOwUXCcxJM0yHhQ8p4cxxQjWOiNymFQu+jt2pDYXdZZMZtta
iHJiYlYvNjB2EIlx7EK8yJ7wOdFglSOjWkNoNA2LgMSwHsnzYFjnzV+wnM+V
A6NEOq69CF+J+ni18IvUpcq4TkzMX612V4JlSs221qVum6Nbyr/x4ulGLk5v
GpXad3JjAiictNkV5EjqFGdt58plK3sLORtGgueuqTJohrCQzPvakQYa6gtm
Vm3rbUrzUPmjsYQ6jvGIWr/2CO5DODABkhDIIPfyBwfsuQdWhVsm4GMAECLK
sDGOIF2ZAVuCh6IN1cFsU4F5i2m5dRYsGop2B4D4QbdP0jHmrJigWyiYeoKy
kTWDcOuZHUnJk6NH21tgUZtBGyJYOX95/4oOEMGFcr+xkfww9jhNKAFTXuvH
o8CWN/aeF1+hH1QNTQtbu5M8fzfzMw12ru69wJKsGzGX8VVFwxueZTtVtnHA
4kOfOAt074qE/DLw0POe0AfcPJt7YRolxX/nYJ8mQ4xfjryRirU+DUqZ2kBJ
gmgFS2jXCmToCXRMiMZbujNqDWaQl3DzbGQEkIHTaL3HloJIy7mUFyQWlZCF
gQT5xNMbUaAXIQbPHOmaKhs0Doc7W/+hcsl8JIZWizEOxUypwmoDo2WjOYJ5
R01xrLqObOGxyEu5ryJW6gXatq/vzwIHHZSZvc5THAa/qn7BL/Ui4OVIN38e
fk13axkrV5DtN0m8z83ps200RFRP9HSHDBl93OWv6JYn6zqdaY8HURhgx+gF
t/9gxDS4h+F1kvHy2zfC8I8t/qvETw42oRciDmFYCCUaJ+r08OIhoSPVxoxD
ex30HhVG/OkiQnaamL9EtK3JNTgqQn6CXiclGMGv7L2bI7v1Sjz9uEdTpywK
VBfKemKbCNFgEHDFJk5zWwS6fjWBFAR+GYarOjMX2eJ0LSlMPtm2CtRN2qDh
uL3CX+I0LvwfT2p/2ODWBlyGV3jIpQGaWTzN8jnwGWoIflGqw6h/CJ0hLsSK
1+uB0L6YnVwYmB4VrQylsVCv3Erolgxc2WlVbCMyrD11gWlbhkfClbRmJgf7
yMkcON1uVtSVNJD3NtxnlCUHt8FqTKHPwl/QG3I7fus5poKPKXUfDoVAsLny
5Dxy86rJmR+5AsYlBRDRCdgXhU884XkPiwuBBUNnJRPf1rpxbxH5uPz8Ky7H
Unp0FedgMTiWMnS7nqX6LJUUubf647y76BnfjQOyWCaq/xI78ebSA6XL6iHR
wqlrr4NZD96OU794HhtOT3zk8koIwhkS/mfKI8PZXHVw+dYI01qAcIocDemk
MovJB5zUUksbip2111kJC+ZXJgo2gXqR0dkGOZm+OM40FpbtmtCFTNeU8o6F
N2gP5bcgplArj0hIzpd6DLCrF5HzyDjcEW5UcNlM3lxSO9x+t2sTnRKXiIwB
lLJ1KanT17Apy6MLIMjzJtNZipeOqH8T1zkrR98625ZVU7FsYTVKH+G8OpyU
VmkV8eUCHbktl+N32DCLauI6MKw4aHL04EZAd+stuL8YipMKStRgd8MQbKNE
Xm8Ezrw/Au7FZOxJa/yF64koIaP17p6Lukw110q3Sd/T2Z5jgAoRYHS78kfz
/tlf3tbmaxArXXoXa8hGWc47pXGqIQxGAooLb/2pDzuJkJJ+y9DdrZmQ/Q1+
N4WdkOBRWHagyjrHZQ3LPuRJnWAnG+cNUaAoljsm5Dnd/nmPrS0b13KnMLz+
7JhbQFCyn6WZ72SKVivLwfQIX2kPsqAzvQbBpJLGPVG8ipirzV/HSVaThNCt
YqMLZqCn8EPfKiBSqYQ8LAL3/tqw/T/edwsocsoDN9BpJyzH1jSF9x+R+osf
kSXIgiTfTDRQUBlJAF/MGbLE08tEruABTBWnFRnoF3pF/pLTX8nLyYkwBfCq
0gmAAyKe/4QOBviBPVuMH3w3qxu4ELlwSnKAyHIwsKaRd1Btus2WsvFtIhgQ
kd8JKDHHqon7hS877488jJIg8q52B/n1v2px9prVyI0bgXGnNFS8TJGEbGkM
0TBGuoyTEMwv323fi7oLi4+B7qdGB628TM0bWsbr3Q8GJgklpeDmE+9BET0K
t+yhYmGlxPnU0I5qxOqIGGj1xz7NrHspgVYdBOCB2oeTN78xAvseN36dlFV/
v7dgwjg7q/Qv1Z4XqQYmT5DFYH5WPrYcadUSfDUeK/GQU8k1i0p0UzFKIFi2
1sRnkIVFPXjRi6Tve39iVa8Z5latTSf5pgkEh4qnxvlcj5ZnAS3Oyu0JRsYv
dz+gCLYtfoZ42e/e5S+Z6j0p5obVbQOE4fTlMuOcFq8e8TRIhBad3WkVuHAg
jHVByjaXUAuNK33C0px4a+Rm8fQ0TZFfeB1biVI+q33l6mtkXPDG4hBroZzA
X0RnvLiW9yQaVOGiuj5RqJ5elnHxdQnUrcVWyv7bSJhXDl6vY3+FLChdtz9o
eU4EnYQOuxGaY6Qj6sAjt48T2nOsSGhqDE2S1um4psyGoydcykbbHwnpGjLm
TkgZfyy0Ba+9/NX9gie15ZdiAh3vBDBIbuoTol/R49FoIs0e/cf53vd2Oz86
UEIOtKfLltKd+5hNmpn/E6i4r5L1rExvtrsDAYj20gcKAZCyRcjaIG6e6UY0
wvjLwxNV+VJJsLmi6OnURQWHHA2wiA8FVT8jIxSwqRzRkNdEomzODZeycdXv
OKgcZOsqtN6tTcLmSczKgo6mGy/LChlvbsSbFowK/eTDwL8vIIDuR3dgfuB5
Yv9tCjrFua4TStwXB80/xgiLJmnFIZxol8DczY78HkJz2j5hGFjkKNXGT0LX
BS3gaSZjF0cNFMjgWZsLFgfU/nyANamnEJd1KQwrU7xSu4UYbbrO5sySwYmh
2rdoxOK8vdNLZIggpM+xwEHPwDb0tThEtIpuVSsOvk//3iLkv35NATF3GbNm
dgvw4Ha5beCGCzoy5HyJVYXGbS9E3xBh1uJ77vyr0gEWycL7wR8RPg1On/0P
UguhMyVRENYzquvvgCmdLmjDc3RrZMAdjgrNze1U2NBfznPy+dj6hIm4/PYj
caMP9RVCJPqZM8MPxG3ZiahBO05mkGh09maNBa571aAZAmwPxQlsBqPvkhDY
/ElkGZmUSrFLTwctXuxJ+bWmY6yT+dRiGK3NmYBiYCXz1WP4iHVeDTP56qOt
4EwUn9jLS40ul9x5C5GMKT+S/nIccV1R0J9UhVwBiNGwbWyR4kpGcxObfcQp
CTEQz7t8ZhVq0eEHEySjLediFoHQ1uluvz7XkyzZ+5TmhnadGIdzURAvJOhG
E8NvZFUkr+yRIJUeyNAbXvUBcDN33H8TQTfO2KC40fg4qKBj8ZDKxuwlpZwL
4qGzMxcRLmkdMWVXvjEFdclNGvF3TYaXOiWStylUZRfvHi7YQQiV//EbRg28
u5K0fzpmQMJx4+sBuEfJapXDb+wGeIxLrcsYZ9XL/U28lZm9N0co7OsDocUX
V2Eicb1czs68kxukEvwzMnmd53/x+y6eS+XE9Mo4fe8jD0/iw5w2E9KMb87W
S4Ru5hPAdKgJnf0wyrAMe6L/7ULjwSYDBsppyUdo6KXupHdnGaAJwA804IU0
RPvWWQ/XdMtavTSdiQMxdu60dS/4FMzt6aCEMHtypOXNUV5LrtUUmMDyVYFf
KMoAV9tKfL/z7YU/icQIiqjNkWhSzs/zgOxbnqlF1huEMm6yxpFsuPvsusnH
OLPUnBNHqcwsBgpbNPfhSeK2aQg4Do7Cq0+jZC9U2UlIsur4/WmDQsFC3Ca/
CELrYwEx96pFQSEXxlrWOmRquUhKubv1q+UvsBmmrwXQutrz+/hJZhzc1N7V
ew2jItZyoTst2FIgsjtB3DqTJVqDmnIRsjQ4VvXvDvlhONqOcH0kcTvzUUGn
li5tfxqwxpJ1zldfqYK8GrBPj87ex9OPgWWoBSWzJaLhKrKJqsXW24X4fuwu
t2w1a+eKO1++gswa08eevkaotQ4xsHHLVnUcYHEQDkK+i3Fe3PEl7aRC52p3
Ip637yeMHVrwxHeUd3KwdRty79gzR0kqy7I/SQMcRYlSZhyNZs6NvQZ7Yg1J
SvY6RBqpTGQ6RvRxAzBB4s7L19XPB4dVy4dVfHuO1lZibL3g+oSls75c1l+P
Ny12x6m4Bg5rZbFY+BN/xy+ECsJ1lCrBSE3zhzPpDLEYFzZPiwIVR0ccWyak
ciE6hU/vpMxyETxx23uurYpxdLo007Odbaj1En2q3Ixv/JAz2MfiZUXzibQo
yHFHTr4Mbbj6SDcw1OkLR9Q6iEjKeprot2fOfWeFGnI+upCgXl4zLloGm1RZ
6d8Vmu/gd04/2z2FVH9p1Z2I5z9QzL+HEDHHC3As48ac4lUjKoPLipP2U+7M
FJSenMaBPz63dqh5oA8hulSiaH18DFlFs1aQKClBrN5NIKkDFLS43UehFNwH
qJtIClIRoAzwqaiPLIJQVAzOBFoCmuLUsmGcQpqx7eDoBcSKhatZBuSVHMNP
AqWeyL630a0i6COOc3JOrKKqmU17p7SaFOa9UimvVmOJAEymCE8iwpG3dtwa
7aI+Ldtx+rI5uAfhHTvX8nbGolCuG+YLSAbU2ORh9mof8A9SmhkY1SJZsF5S
elkwVKos6qO/WebL5KCZ8CABOIWBZH8kHZDUN8EDW1h2a5+6ANTvHOLFRWDD
X6zD0A6YVduZGivp3N7iubtGtacZbxLoT37HSzjwtJZZg6LWq4zibdvKO0AF
RsWCOcU/H3MltcJ0jHYC2XkZg+Qk5L9mKcwHXxTzZn9f4vZ/B+0jFUBo20Gd
96B6lmW2OD+YDer2Qiqx+tUXQ4m260g1tlFP5gQom1bUgRf3LZNn3kwbmApe
sabY4KaDmSpwfrBNccgkNDPlc8KCddRCqgJfrt2Yx0CnkGzKfuAjepSH1od9
1EytEcYLnrNkK2XaK1eWPWL30Dk7SDCZiMbC7Eq8l05DpHbGFDnaUIvcUi9d
PQfjbLz3LVXD4pry1N3eMqSadaZRIlJZmY/x3piaJUpq7VLYoREy+1JrjIMN
yo2KX+03fN8sFgmmet5yAbUOXkhao9zPdOWS2773Ez97QgQ3S7rSynv4YgUJ
rFy7AEKNVkKCIQwqDLFY0jVVQnxQHBema1lQUOhyqkd9xDsBg/8SQGHeFHp6
5ZcMdFox452mW1+oTOiKx05ytkxTss2jjxpswaQs/qZZvYk1mkCzy/N9mdvt
tgnGBC/xxWkcsHi/jbfR9jyE7l10HllwZDK4amLanDrsb+yeHGGoK3+JfBD4
YT0miQ6+9oXXCjdtIwCl8RgRKcltfk7eA8DITyQtrr9wAy7UTEcWCzipRogD
Y/fI7hcBI/2/JH0wyxodI9n9wq6dF49pP8ws7kCUSeiUCuorgt5OKDeAhHAW
4eTnzFGN2i2G+EVOWNkor7Mi3hLecj64jYIqA/xtsMh6C/ogh9N+nr0jlcOH
iFEoIE9K4SQBWMw4Q6U0v2ughcTJlCGc6xn5LXHdPVYMU+r4YDv+/xV8/dwg
HjUMNuh+46Gr+4jR6TEl5sDRFbiGmBijWjEj+nmQfd++orgYo8pZOry7MXzD
c8xUUw76pVmOrYoZ5JA1omWToXGR4atX/RfW332wectOAoXvLHCya1NbIxf7
8ONBCKV6fB1NjbaXck1OkNg9r6JVobZJIGd47gIQCYjyVNwHn0GOFkYtvHSq
cxq2qvyRxuyx2g/x3uGy5hTY7vxdkaa6rMMCNZMbCek764CAJrCXcaDYdc7L
Ac+nLBz1fOuToCudLqrQEAy+BVgby6xutsRb9TYNKRYPdJo2R2UafdJhOitG
wUeu+VM7KBIJ7ErRXAyqpnt7/01S5ay4PXzyMUiR5tvyJZpULO/U5pcjTWZW
yvySVt9VhCJQO78gTE/ZhTv7jS8T9gJ9e0DGSR83yCb64Wfz/ByGUyNk0n6v
qTITBysJ+8y9Q3UuJ1lO+0kErE3gubTQM2hw7mAcftb7g79DxwZsqIw/PKoH
7sh07lq/7aRDwT8iihzQFzJ9UaneVN0jINX4smzK6OBGmXnEzsVBpgv6o6Lk
KMV0iKuRpY0f/+DVkeMJe9qi7XzAiGQJwnU7738SYyCG2dCp8ky7edUuMWqi
IwFNPC4HWO7e+Yd+ejRgPXS6w39QREBJq5OGcrqa+msj/L8OHl0cmWzYDtgA
+z25LmF7OF1gQfhMOKjKt9vcplcPoGE+OCYbk0iiBZeWz0PALoPAbhT2Ewkb
oCZk7EsqEsNlnEJNNOctwxIbk12AjaDiZknwnHMafZbUBDI1QD++Ottkr1ij
8FUXIWwJq3aP5TgfvBr+6iQ1RL82bRXflr5lOwHbEGZUFsiECh0H8jZA6u49
ZB8bVg7pDWbLh4Kuq6kSdYZkj7ZPdXnPSBL/cttrmML9jLOCHSZgJ0zME4N/
9x4kh1STTYXgRrQII1XkFaVdXzoo+EI2M9VONQYl5zU6px3PXQak/d/PuGV3
/cu5HACwmN5UiqTgQlyduhSRQByphkufSsDj+uN2QnvPJ2V3Veb+3vM5yqyn
HFZ3AfH9jT5CMCI/JTM0Za0GDIIWIkn8OGgnWxLZekRATlR1cklpjg9iVCCk
w12x39i8gL+C4je+k9qYhcb2rDtKna49Vyli8swF59nVFd2ZXEuyVA34JaEM
/jY2TOuHK0/PzYed1r/1o4GqV76XlgMhldmXXK4vgjknd4bL1grnVeauwSrD
qn1NN9mbd49KrKETjg3s2XlFM4Nc5b+fbT47dW+KEOxR5nLPYpCjijHVLCcO
+IopocVaIIi/fKjZ/Hap/ueJpg+hPT+fkGkNrZaD3ietxVIq/vHim6lRyjLj
bAlk5HIKBFsYZDkJBOAXEa28l3TCOulogxz7UQ1lPVOB8/hdok+SFqysl2zq
xoNDRIPm/4AV/Zs/6ooxb0Pmjwy08POSjEa5qVFT3qS0z80gXhw3ubcpSSFS
VTF73Jj3Pj+v7Cw1it31WxaNyuRfqOKmJ7zQNbTg2E9+fJh82L4QDmhVZO9Y
vbGpB+p5LjNGd4dA/wsoTTL+MqfBQU4X3rhM3jzTSislLmVTkKop2Kd/1NYl
KuzaGnYrZhehdbc3sBZyDGqCQ57/HuXzDD/NKx2cqy7FtFqkcRo9NTBhr+F4
qGuAUQT299x+tmE7wFeRakzEDTNAInsPoUlxoPxtKuSI26J2gsFtoXnH0fgv
Np0sdj/ad2WC4I/8/zcocjnygjwK0rr8j1+cutUKUxTNsEWm3xUGfxObKhsz
qWSyp+A8V3SUSo3I2CkU1idcFcMputcptEVbXbvhuvKnCTzU6vPzDyrL/hf3
GHdSqJkBlhjTjn0rBREPBdA8iwpMN4tc8y6J8vG23xX/E5d7eh9SY/+AUSuy
3Am4xpQ9j1KoNPrkVvBiqLy56kpTZwA5UB419HLlWK1ifVTU+BFUNb3kZO3b
YL6e+HJUzQfE9QK+sttiWBHDqoBFm0L8s3W26kWdfTRSqMRNvxlofjNopGfm
5RS91F7ksblVl+HLNoKxv3i9CevNDEn2F3YLJWsRTjms9QcLyW6ylfHRYzid
PXUSurVkXv5efZTONFOP1Qan5ihF8FWHRbISqxyXD/vapVDO/M0SIZM4g2F8
MoSt4qmryPcH1qXwoaP7POaojJqH9poEK6vAk7lnAEOUsLyaOFKnvX+rmHwZ
WGnq7Apd0Aje0DgitN4cUYfhG/Hj9o3C61AQFFaX/eZ+Bgsna1WMpUFCIdJ1
FzZ72ELvAqNQQIa2PcPXx7gi735kBfZ+nNQGl77svOCUgOTANETWcmI7LEMc
x04YvIxxTAyPYJV27/y8JefUqgIxc5UN5NPAWT6EtC1t5M3oUKpYz5KXj60C
Ik+8TP0SY9/5k3vfXAlyof22vujNTvXTajsdUEWQI4TjrWgWi+R9f/ZDeHrb
X3W4BlqC06uUUUiFes4UgGRfVvmvYF4j/xcZ297fSlz35/bY64jvXhgXNJoJ
6SDPe+Oyl2iT2DDN3h2oPfDA32PW8XCuGfGczXExHaXSBK54irtQ7NjQQW1O
l9yeNciP+K/Rydo92rn5BraxOoAGBWpoHWt7GP3bHGnSX9p1Szf24MPlN17U
Mw4rWtRFE3+uis3yitIaGVg91u+BHjX/Ci0LOfQsoM1t5H6LtdWqx/hEUDdC
/bay5nIaUlkKOxvSYcRqziFRWIvKYsLIrhuoC6fhJVbrsqv+u3lqVP3eUBhg
xoYN5sbwtspEndh4C99lZaeACqPFgVtysNfmzv6t3q7wwbNh0fGShYkvIxke
rOCMY13hOG5TLlu8Pdyq25jVxcFNPvdCOxwqlBiiXiiCRB/vCrrGYSqnCQ6K
8dSX6L2qD82PfyESXTZbdy6AYa9o2ZeFMXr6gEbZMK46LRDNdGAJ636egRYJ
NlSEIe4iqGYwHT5iDxnKHpWEVZEh7FZ0WEO+61/x4qWPrWteCfkjytOzdsOi
2I4ZKNtzE0Gyhu8Ro4n1c3Ima+FWaCtPhiliELYmAGYhy9KVd2WcsCrXQiqq
wFHEeMPqW2U/f/djETPR8Hf8CryI9r/o5q9ULZ//MIxrcs5jGMH6htslPsTo
MAgFD08/ZVcaVrE0CsPR0arctX1IAZIamfyWG4mHFj8bAmkHMMrCGUK2+oHR
CE00EslfnUePWpzMSEwjn+FcqU4hRUA33drSh3f717E5SvZieOYE5IQPyWsp
EP9Cu79FuyrCusuP328j+3lRBl6hm7nW3Nhy8PAwASh3glEZDgsesbm2nWc3
DarR2OG2UgTKl/JaRLDotRrxSBfsqhABd1hmkwQFpMQPqi3OJlnmdKldn6pr
4f8Heq7UN0YN6p+w6Px0oUh7AlBKn9uHhuAMjF3Q1DPR3F5tiBq/waDZ91VQ
1Eg9OXgje8OLKG9QI/S92xkY25J+qfIhtf7jWTy56pp85ph3siuLJ6A+OLss
7w2JvwEUBN6LSKdkEvJCnWWnLyblaL8Yny671tDQqhaq2WH8MqvXAuTZkDKs
j5/tiK29Qjc+T4myS24pQAMhdLssohxHSLygB5eXEKKoe7bdZeFc74KBL6ce
FsEI9C9qW/Go9qrxLNLF/rIW21mXme+Fdu8hkJH87OhMj2O70V5lxvIcxxVH
sowbP4FC7s8Qccmg7P3XQ4NJ/vJgOvvg+chhxVTOp9llvyJlLLnEMnS/qIKI
vLvE35oReDFP1Q9YXf4RpeALcZOHmUzsuwNyUqyYOZDd4tZyky73znP4F1ZP
b1O+jI176CI6fZrPh9DHQgVPAizCGmncfFUtglccbtZO7xUgZlGGSH1YEvET
tsXoH3TZ0tKV68S9xjkm/+rgiHfyPg+7ECDh1AHX76y8XjBGTSTL7l1SoH8+
ZqDNu8mLxYGwu/wq+HdOF56NDMDvTcZgltNY4D2Pgs/fuGyKXFfD4Hx7Q44l
3mplcjpTZ3W6pl8Kty8clfYbk8weoR9OLVqjHA+KzX9+CrAcIVFFp2xrYKhJ
5vOSPBVbAjNBm2ansVNKBJ49AkcW9hYc9o8pgLVn/+EFbonk/pLh+EZoRQ7q
wMhJUZIAt1iBwznKSyF1XiGpooSYs4kTFUSZiFI1M6tvZs/00LwkyLb5az7o
7/iAAIAzHDjy1jAdPDcnVaIrO5/mN9R6vyvLFLE9p/u3tWKAem1HdVYo5PKq
Z3I8JlS4kkoS9Oz4cyRZq1ASvRaLsOKNrjztnuEy0vBOa77vUP50ImonVLLe
w/1pQRuqW1ohgHa93aUhveHcfjTxmYXE4UBsCoN8aQUd6YgaQV9Om4YtvD2H
rRZr0OzWW60nAToFaZcgD605xz8Riax7bZumva6oeLkpp20twjEp+GPUcfEa
gnLeZZ463G95XBP1gGq8Qp0ptTH9eAjsxoDG7Zm9691+nmVqrSl4i34TY7Px
h1GM3k3eHxTbeZKXne/XsxyiY5hpe1HDakjdZLyQ07usU0LTuv+0a76B2vni
O/FoNlZ1Z7n0L0FYqyaHDeH9TZcpy5w6FlRThs/U85eEAWt30k6oQKXXzlwR
pKGj801MYZy3zEod+56ugqfZhLbwze9Csbg9omcUQGDdQ+ew20e2F71d/Hum
/uddbvS+FOlianZ/gAjed2Zis1qJikwG3sMaS1mmfkUOTQgdNtJb9iKn70UG
P/xZn8dbs/EfmyaLeMsHQeAwM2BVNYYQb2BRFupD5eBXf35He/xh0d1UWcFD
11bwXBwqux9JvTL7SNmBVlDjUXPR5Cfg90lWm10Rvcy3q6z5mVfVAyLi0hJr
9//WAoE64pHi+mxDoxuiB8ZlLkdkcRc3C6edw3LBD2LX9Gcz75U0BiymQSwR
rWtPJrWLDkxLCRCppLuJjsWwr5nUEzRbLbnxczzOzbDcYBeKH9GPViSN3t0b
reiqNiGY/tDX+sr7vwrZschWItcNd0G/mMGHRgsBlTGsir6EhVfPqaHHwN3s
i3Pd3Bm0cpyIOdGqcQuCiLLrSQPNE/dt7tfaTCQWo3rf96KHlyqwpqgcuUaH
mcNYy/m1vfNIPSXYhiPMx5JQfE6iKHjy3v1D2uPZwtgH+017gsIWsY2r2l7r
HZp67bZ/UsEAptedsmtVHjrXrOCfHee8cdmOIBA03qX34kCGKXQbrALvMt8J
ZIrSx3KCts2eUoXAz4Tv1S5MqqvPRjfiB6hAUwrzQm9rVAXUo3Mx031d9lLv
ISzRGjS/u1xyFRMsWamyl0RTcclMvZTscQoHkHTqAVaOKUVkVlQguKZJNzys
I2YA0s0nHJx/yqNVXq1iYXoXhB8IMcFL5hkoQS+gXonSekDIqZ8d/TL8+CKs
2VehVsqvwA3I8ZXpopQUTsOAfLST1zMnJJi+2CQpbJXOBaBzyGCJopryrP+u
6heAwa7hSZFl54mw6bMLNcCkpv57PeTN0YnDE98SK/o1BXfRFt7QYcyrJWE9
WGraafn7m2GLT+YSlaCNH3dztv9CVFibVNb1UzeswqtGkx9URk0FFpqXvNWF
woh27v9TkFE+GdLiEgR31Z7qusL/bqHZgz18YhN/Ajtiz0TZG4GtoLC4FgA5
602m6SHPSagWJwtrx0FihQ0MrMv9PrEK61iHIBq+LWxP9rR6nwAOLno6TkYy
6Sx4oEHMkjgVaWrPdTXhpQQqSV9ECp0yJTPRAsQxXLRbn63xtDvpTR1IJM6M
Qcze3PYv1948XLsLm1hU971xqhc5/FlSnNnnDGHNgk2T7LjxWtUbsRO8cXfv
+EdvzPoj+PVm9Y5ZKcVz9hvfBoXE+fryZ16DV/1+Akz+wrg7saKu5U7qUxaY
AvoiDN/SlBuqhIMk0G3f78481Lawr657V4c6uBG7o80EW6U8xbCPpUe4foLJ
p6l20Fiss8GnaEc5iRK6s2HPBBPWf6BhshO1DLr3sBNOUPiXHyxBCvQnL19P
uFe8ga6nKXeG82HwYCD7c2MY2PArLI/gC4XEYmR04QMjkWYHXWkS9I3UtfNX
y81zS3ySvzB/mHiMgge3hzC77eX7UPSwnClHKZQnq875dcFf3KQnERJM51kL
TFUHFRBENwYrguaEmfOHPQqlHJQmxCaYKUU386i8VQbMVQ1OddFjfA/lj0L7
gG89VMoHGswF3Q+UUHWacGih27pn5RU6OvwJdK2cO0FeK9xMMrXghxJYLq8T
TfUMkj9ugH+r1n89HxRWu/Q1OCcsmEBO8ual0KKwAml5xUTgvwdDE3kcDveY
5tKw+ngnIqmPW+24DS5G2V9K4NDzQM3Ry2JhIJymaVFxzUgZBXnYcXO+3tnj
SXF7roMrk1/IchfEsDSpHQdKzFLH0w88/Jw7TullazEM7xAFYBKqZiPpPDOD
jqfAMAdJF1a7KZBhayXujsQ4tEmkgYg+AAtvs9ptfwIipm8VLUX/qO73cZo9
10bOQoS+PuXL5LaID0+f2gh0KbxYyR7ETkLHIywNnJKjPwLctSblC3H4LZ1x
XNwrPTt8QzTlFAd2UdqtuZJRTii08+jyHPUPzSdlXh1VxhjqXtQ2r4KY9gFN
xkMX35cp+qCdM2lTl66UnHvL9eefyoDLRkBBTq/knuDMhxo5+MUrbOMOTJI2
ETzOiDmNcKFY+7jY1CgTlDyOywyjUB46D72MhomDCwhS3UzNwJO3fJ++vMC5
jj47iXQrsceSzVvgUkukBNSSdEqhqNOwxfM19a/XAIz8hPYZiAVyvr8uC1fM
QWJijo4V0SjsGKbI0xJuZXDbvLn5BCWitvKwcHFlLn8QdR94WP3dKFiMi3nc
6yqNMHFpMQ3N56h/3jtPCyT66jd/C2/UlJh7d8kk3+5sNhrcx0hP1jkNvY/w
c343JV7hHESdtT7Yj9/+TZpRdH4q0IfkkkMd7xoUeE6n0DgVvhUT0N1hiU8E
+dyKDVgAl9RX0WfodTZHbqqBGlqLGdIfGWKvlFRTjHHcaQ9n4P6cFIwqRjEE
MY3nelrBOrc7e/qXnDA+DfQeotc/1JZd/cLCPSqIgDQ6KX2gXMZUm3yKKS6k
7ZX6tN3fvjIuANOogTndyIEF/F9V2augL96PmFh6S1mKbOSt7B5WZKR+NJtX
RPVBdtvfMHnrPlv4DBfRJXQpywuxsVQOYRMvAtXihwe85knV7FYhnBxhrQOe
KQU5E+yIKmLBhUqZWRLfPcJ6nh2cK06x5uKCl9Ddlq18rlSFRF3fRokmOS3/
kiYrRZA0nkleF+YdLKbYPRq9tPhMjZZpWeZrhmHD2WAMDMH9UdVcPAxDW7vR
+XCKIl/kVyz97zWBNeb9C0ndaP64tryFrNK/zhrV3CAXD7Y4HtUzDU9z2M50
mqdps71boPA6Bx9UazQ9FZ/+2iBEWMMDr28Vm0nE9DAB21SK8+FHv7b78nBM
AZe4s/BupAwmLAZWElRXs6nb3tfJzZu96BuS7luOOmGF9Vjy9O0yrmPumbKx
MEKfYIiExSYh+0dYxYvRLX7xMmO/ellPFFEl0o4Lt7DBvesnQYevbK8cwSZW
gW/ASHxVmfBMy5FF5z0v6cqGU1UCP71Wwr5sVHsrk0G7/KYkTCmW9cYZmse1
PsBbYwPQowFC6QfCRFo1mgpiMIKXDf58JbBZnzu9PDgoeeQKHcSkGadsBy4/
gszvpTXcrrh64c/p6ueZ/IoJ1MsU/zp7Vn55FPRiBDZnvaD2c82lX3mTEc/m
Pnci27/tlW+m/cv5PyPqvKB3st62X3Lu6UrR+r2FzBTNSOGiOulR1981wA/W
LeFyFwpZwC73R5Oeuqw3wL3YG+1DgULCl0r3/Qh4qh5MdVhjWIeAphc4vopR
Po0bdnPGA7/+vibyfKiOFI8wszaISJOzjkML8K9GKUYzQGRXjiHSJ7Hw1usd
w4urUjJvgK44GWTLLNJZJm6QJBA7Cmyf4K0ugdAri0E8Tyy7O2HMmcBCY8X0
5DAFX5b/XXfkVlKzWpCwlQXmHdsH2aoIhsAyXluN3PVs2SXiIdUwZxoh7UZt
ivQPMOTvZ/gwswbxeNDxhZ02WDDPZ/Oic8A6X5Rv6PPOR5hB+0SMVuuAlK21
OJ8+4cY7K4e2Uj26RMmgvEAU7wRTj6Kc4CcaOaCzvW1Av8sE8hCbd4DiISe1
YEU4COkMUO4NT+qCD4Gqr8CJnnT4Jygoz8825Xx9Au9OZU0zXWRX3RF6mZxb
IvMf9+ojFlQm7KI79MgW1wzXsNgDnBcEjmINmVdWMEOMx1NWrJ324bGMurqN
1EI1UTEYcBdbL1GYGpFrAH1DTI9eQ0GVwEoknXbVlOISkVAsrW4K2HZiMjcE
gyvQSJqzF7mHNV8/H77eOwMEWnVqIkxH9Z1rdAsFvEW+P+5UxQeUo0aXWbtf
l3Gi/XJ1dTVLhQDdZ6o7LTV5ISv+k993/WGqiW/eAc+l/89/jSm+VQumC3qP
xc7WR4RjGsV7D8obyT0P8gmBxr7CKbOIdf2q3febTdj6HhVnOSy9nA7dLA6+
mbYmWKgH973RVkKe8X4NEMNv85Y3JowB1a/m5p+fBIb36egGngSL8a6+tII4
ZCUTFw+q9A/1fyEV3cLWvsDLI4Nl7Fw4rmdnAuiYAPvVeNlrDH7oq59mCW1i
Eb2lvtCesdWkbraK/f76v722ZXDJSsFacK8mq5b334o3h8cEOegBxswC8ivW
H5BSO7N0kdLO5qPzDfZpk9hTdILc3+JCXRf4gtq/LzXTLz3JogVZTIHZNOfE
IfjWw+2+3LW4WR8YtyoR62WZBBId2MfPPSi0Y/m3jhh7n/RMALWqt/e9jzWa
2y0lqWpMIgqrdvmmwMiGTgd0vHraFrJ2uoqZfxuUb8/sn6BHWBg+UIWWBnXI
bKiPONtvuw4Lm4biIkcmrUv/MGHdRTVF8EGbQIg52CyF92kjA3qKx8a3CVvU
wILSMnUsvMY7o1eAIXVWuPHkCXUlviDiMX53DdbNvHiKeXh4N3bg6R+CRm5q
dvxcTZ05y9QqoJuPVXGmql2VDhR8nQ803BvTy+bej2wXDL7sSQJM90mD4x/0
dYOAx5pz0VGTY0z3LAijmYsTAIeGXGMrnWlZbjVV6lz+JBABl38mh7K5UfST
5c/z3gX31hGkemnnz77shkooSIeqn1tD7mfWqGrRn2m4J0VT9N4XpWJXxCpn
TiEjUIRBQ/3Tk3eErdCH5bvVSh3EgATh73IE+pUB4yDCiTiYcZxIAAohfiQg
j9TX1+LGBMUCtHQlqLUStViv/b2tYOxSwOeqqy1Sf1KtRYzux7dIuy6aRbky
OwFgJWndUZB8Ta6uY5iHXSm+fpH+XfwJGVJcTKJldR9cHvyZwR8FTlThmQl8
kyCDZd9JIebvGxXNwZwRrHL9633I7gfjLGZYhRnpzbhrdTcaE5Ypv7mlz195
7OFv00kR6aXwqDFHSC41h/AxC373Q23dOONi6yc6+sdsazp9byKbwdnyEerf
BVIl4fdHiCsF3iBfSP9zO52qL+N27Z7aEiZ01XY8ftSKMvV9rag6D/7Zqq8l
eoTTzkw0oc60SsEBlpTOgXDE0ndREzOIiD+9FRL6WyAp6tXnvcODrsMQCn65
oBk7hSVPQFOkvnSmR7F7Dda4MzWBEhjGiaDINVqiRVO9OPNIdetEqomVytQY
W0Ir3mo/dANMXGGK73Y2DZsgy0H5u2prwyW/6pi38gApqF2x4NPg+B1fln1f
25peBT59wE/ijZnbGQAxKOlpa8O/wzVF2qSTXJDmj9rlWqZTJ4/0/zFTSA8m
+H31CC6zAlClkzCe6KrR5wxH/sFsrvIJuS/998DsZp2RYlyQGxUGLQGl7AVH
7EyFHw1d0uquwwD4M0uKtC0EoPBSotvvrU/rQC89VzrPw/YbP8U5F5nhhqXE
fj5N9XwYBnKvWqAlWcBtyFZp19/z9rSiNskaaXp3gEetUDA6/TughrIg8VEZ
3MG6AwiECnwkdkJb/yygEy1EcO6MZ4GAiiEPXqSomoEkrxoDmU9b8NEJ8Lfb
3k9mtqlOJo4Id0r8+BbSoK0sXGdURoxEUlOI8SMN1MFLvKjMSir0Dd2V1Lmz
jc4aujExclysnGybbWQ2dUsotETFIpgVSqosSbffB3sB6O3Aqo47o9/5ctT3
7+OH4tmZ89xuQfYf1+0gujg5bVZg9rXimA3AgMXUBcIA+T84eoJCopy7hhSd
PiXyFqqm8zQJ4wSzX+NJVSy5SwSlTPod3q9kIGIRuO+MI7qJVl+Nw2quZB22
uouoSj8GFNruB8bizR2kZCvsZO65P2EnCOK3jXYHnjEgm4iInEeCHHO+MGa7
RmLUb6ytCcGOlhqANwiohuINqk3tWXortxWh8Fx8BmhCQnQxHq19sqzOYQhe
TmUB6dSeSPeBWeLMXmAlf8DF+xqeuims4D6VN0qHVFv/h6rrWdlb2z1r3+wr
KViPll/VOkdQ8S9XO0z9NTC5XBmeHyb5krwx5P3rnUPnkY3JuxEKyFOYHiEb
XZdYk7+a/WtADjviaowsefmwomFLBZ7Qprl4dBQm6HQHGBshQoX5s8+S15JF
Cc7nVH9IfXhhwjFk4UTiofjlFjBsS4RhiDc33KIND+FacckzRpYLFHU8yCi1
X8Usp95OIXAnbhNL36FpP90nw9tvsVyekJq9+DitdnaFN56sIThV8FNfVGLC
GanHtUTOEgXG3a4C6/6taOE6d3sUcSCXPbRBGKv2x04DkTPYmdr9BbxQ7wq8
CB0zACP8CiFe99ZPlsJ7qTAaBwhmQ197LfAd7NLFZZWFP59aV7yzSLeEUqqM
FXftKBDuKTSJ+haluZuv1Agf2ymA5AT7A/9IkmOjb3Pa/fTXdqnmy74rsjzt
oD1BY8N/SgO6RAbaY/vt3ZU1D1mVb2yyf0y4rGrvc0osmY8F3uo2qYgQL/81
loOum0YwQCfPqryFtkFkS2QAX8mPFI6Px1dzEtfgtCvRWQv07/KE0e/WoKJC
h644HXY7UUsa7EJsiB1Mr179zco7vdFA7FlOguMpL5UIPoqCzTM/WHIxPG/N
C1bAUBQu/oYArEttBDRNSoObQoS/iYHPLBt6tzq9e2J91Bi6j44ulvaNo4RJ
YmBEZW4L2d0QPBBR8qvDD4BfeKfFyRouQnfQvjVlNgX9Mks3BHwP1kyTOCIz
C/v0nvzJbz9ENgd1OXOVF0LoU3MKpd3trWG9+S0pRP8+JyvP6VoB+6ZC7oLx
/pBBT8fpJgyJMqvQNq7i+pUD4VRNCiBfQ39N8QsJzXzXtIm0BtDfIK1pi2eL
wGVzxlTJ88C7E1P16zmrosEZx48qjje4TOL19QnRFXqjboNVmv2EbwzjNNdH
0zxSdYo+FKO3MQWTk1ogNPYmDz1CwUOaWRNGh0Pk+64EV+4drPs7rfr5PyA/
tyUyTZq5EZLn5rBSRSjQrYSCq8Q3NEvEhOwJf9z7FL21GFJKy+ChY3/cbfGj
qUUqbHK2bHtQD2at/pSddlfB009uNOeMOdFHigCZGAISY+tUTOvPWOSQ5URu
nNxN2P21/lbU1pEJyST9Tp9cOz6NFLBjY9upc+qAi6UVHD4QLvW+y796/MBV
xtp28tKmGiBtMPKbQclZdlN3hge74WA9ODWWsroCvJ8Ta21sdX4sL76P44/N
h3w16V9KqVrCtQobJdkXX0GCXlkqFHpl59dFdpxmRgYaG67yR9Xkpb9G4leb
ke4hmDErPuGQL4HZoz0tV+KRlqcCEknPpX7xJVBBzgyA5bQsKLRM4AM0mVRd
SspoW+vww9sT2m6UMCGrO6ke9eJy0yYSUxJAQnJj6J9aKEBWBTTzMuMJotGm
MVFHr+OiDoW2nmuXwkRFdCZXeny3kvTsPfGpAzfobtwxiMKc5qbgC5MmWk1+
2ybe9/gJ/UTaibxECKkzlIeZjDNwEPBlG2psZ2IdMm2+GriC1zRVbxY0MkNm
xM7R3VGHfiQdFsFXAEdiVmOmR2vZx/jXSImK0ismN2XK1xBz3T7ObqL+9OBo
UETKzI1lB7d7o7yHc6VpI0GS3xSST6TknYbIvK8e7oRBs3gYWwrMjTLqgo6q
dDEbPgC2C62AJ6JGyhRmpFjyh3/iWILvAsmc/1G1HzIqgq/EUXt1quQREgh3
KHhBQq/Y7Ss9rx+IaCZ/d5bkjx9vSwM6sgv+tHYkcc4EE3BZZJJVtVlfFYAa
i8a3QGBMgJaWPJfoTxANf0QIfycBRW9rg4i4XUBLhiE8yNi4A4JMhm63vVBQ
f4zfuZwzpbUP3sP9dR9sOQrIzhwHrvqn+Qif65FlgDNbJpvtDFwno28GiDro
R91oEdha2YmEP0wSNG1ydjteZmMBbjugYhAdYFkM8HX1IdDNtGBPfdJN8YUM
PWntbJFryrBRBFfcpQH4H4FLCDF5D5BVtQKZK8UoV5FZ6Q2np52h49QJ7R6o
P3sndVRpi+kV4TmDSlCx6mJjxdHZ+8idej+WUIKkYFBmAqRDnrUyc/NqfEWP
pt1baYlSKDcFGAfJkQ8u+RcUyFRS8bHwXyNnwjr/XPtrEbIlP11pkoKlis3g
RyDKeYBPkkNHr/pQl+y9kbdamRCaskYtOWMam9m6ZPC6+rZdT4oQb/ZPV45k
HFff1BOth1igBnqN4nEBOZY8MbAstu5x8QxFNQzvW5S3L47OopG0nU6VGvV6
0zogVSgMtlzF1Y4+KuHszjSh7GfDzCipy/7ChuoVHGYuQrXXscrzsxX7C+7H
H1Epzi5AYMIKF2U+Rd8o7kn2NWJynffk0tBzxToaFzbsLj9QSA2KYtGg3EG8
7+W9U4CT8RZjurRKMzkz5mdIx94Hz5XtKABwJM52DyequTMBcqZa0YKOp/vW
QwiilMVEMtfVIkirjifZG6xhetbqXYXKEu1q56Gg/vLlvM30he9xgFxwLHNh
k51VU7gyWgq+WxHlDtVXH3rJlTdtgE2tv5aNn776s1nZqER21nJberLTLj+k
8Ol+9FR1dMWXn/ztFxOAkarLWavSgVBzJps2K9L9RnzKNSHnINIR5hV6ogLB
6KtFR/NNDlNv7x8GRvgHi63layjzTSgsJI0HS0Na1dyxBetccT53fYYuR9sc
cZwrFf/XWB5P8934bNl5lR6Nb24YJZbp1HMmytf5gyWuF3dHwrn4HqOtZQOB
4jQ5Elkik4jSQLhH5oEp9Oc8+umPHZHvOUKvBj3QXmaJx+SoPe53IRb/Fpku
m6tSJ0sKcPlP24gTXdLe5U4PLtqus0Iq6oINYkJ2fup1x0RYsqGwxcPRmMKS
4oMPBeM1B3OlHLV01prEcvJpt46/DKCQA4fTVKO9W90StVlfuKT68d6fRxRD
u1QdLAVFMI4Kh5mgshLSPdJw0XauRxxnmquc0Y7itmq5QH8NSou62uvId9tm
o1oSPOQn6SE4AqPmlBddAUmqSVwGz14L97zUmzCCFpg1B1huP1qvdAzI9C2/
769OS1MxTLplDMPc78C6Dap7V5UZrrlcheGKxQcZQlkqNJO+O8xrlGvOrL99
biFfyClA5kGp92xuf+fmP/jmJT9BNO52dpz46hHFHZpqpuNY6+NjsT8yGFZO
l3d53TIoQ4aQDHNnJ7zGeXec/0iaVOLl19MwPf6Eytd/aXepv+KkzukV/zs9
ycbAxYx48m3bVYHiib/Mczm44At2TtQWhOyu4Geg+JUrnNuHHSUpi1kYf78x
eEPYm4Azs0FxGj/7ToZWtG/TQppX6PM8E0/xvvZpXQg2JtfrhQJDgCV8J2IB
xHeMkUBKNa5Fee/1dBZJ7h5VqD8yXqp6ePrhf3RpMFoq+qzWl5VJzOYwSNrV
LIcFgUtxC/7w0cNjPCE0NOtrY1AVmpF/mkXHV0Fre2TOF6LJn5Mx1ps/nywC
YmvbwM0KYfMkd9j0yLY6Ero5nGKybxEWhAdRifR2FToeYarfmuk/g14PzhL+
kUtQkbIuk05rqLzmxCKqdBgzp1SHi+dImvDRNiK7uZ7ySYQ4M1rrgULVOgXH
U+POlzeA/ix+1947O+JAeQO0eBA1kpFnCwr0Z+lep6tcVRicYLbBpYp2BUhg
51IhgpiQjWgk0gEq3DZOAaK8PZdSdH2SAP4Xmp/QSs0RuLWNeGauutVERcr+
xs8sluaa9xqVyKojGcNnMkrLeZLtjMNbdmIfjwck2T9ntAWdRrNpWT/Rg9GU
f1JrdMwp2x9ka8wA2dqdbVpjnPctXlmdOhLhKysQvFLO5QHixLX/8tCyoKDE
YqoBrnMVX8l9e9g6gWfUidzZ0o972czU3n3h2JoL8LRYyHjoMQLe6LAf0sSF
EFNgWWLMOm2W6+LQnydzeSUD3mgWebzTiXMHeHBvEgfQ8RTLMH6oUmihrb7x
BrkjFyoT3KPpXTuJ4Y98TySXc0T0cDBjfo2OazQ6jnggkgxnksn6CPG9xfpW
yXTMS8ohZyPWeC917I10u2kwwg8uzo1RyLG0zajTCokhdj1f5LfvRwZIRzg6
3UF2K3e1FU5P19eFpuOPyxJ35TlI5TVc8oOKctVLxljhjxC3A22lspX/op82
+fQIR8AaBqES0ss3VrmDmI8r3jv0LS28IQiGrj5Otw0CxHHgrUkgCOhvoPK+
dZwCWQO+qntud2L683ZWfavKAmsHSOigGHdjauZML3y4Qw5jstYm5o1OWyoD
T91A+ckG38ItRRHxAzGDJ+Ax4JvEpoH2KBnj48SqpQ0PG3vI0oA88ebkYPfR
6Hn63bCbuhUo3t3TP7i+kMc2z/+FFTukxA6ZcbOlxl0PKh2vDQCmjYcUwY1a
AR/++Rt4GyfGt9CU14XRTtiXkM0ZiwmsnsZHCHTGVXYXdc/nlP8DW6noOydl
QycS+3xiMxXpDbJm2PcXAYnSKyJmRHQB4wPBZEW2ncyKl1nxEFrFmYWHJLpJ
TxXJX1PnFj2/OOlw4b69Lp5961hQEC1tvUk8liNOjJ6rFUY157KtDLGufkcS
ajgdW5iOXtfas/I9FWFPYHtNODlULXHt3jFzd1soBdQGTzkI85UIwrFneJXN
dpEAjh8bD3tE/pDiJv3PemRcKX4mnYGVa9snq7RMkSvvX52mJZ5kV0iE9ht3
P5A9Ti10mmaHLOTBeT5HLF07942nL2TFxOA0cZYtBtg7Env3YznVj32vwav7
6WC8L68RKuV78oxVo2bDDSos9YUL0B2BNuvUz3xlcyfXOAZeGLD2HRWXkYyI
uG57W8kYu7B6qUHc5kleey+OxfyAv5mrAT3hUOqknup92fPxp3DP1velBW2s
xcnPYstv5loBz2r9fD89Kt0appFkXIrbV75kfn0LAtNG6/GVpWyKpF16jJrS
R9F9y3NeYttYVwyqmRbOVEp74LynU/46/9raN2UaGECdthEZJIZflHGMVMlj
AW6kXvJIpnuuUhb96T9ZtJG5b6AvVmbfMLXOetvie1k/W2oQx4SODObMWUkn
kDiNJNX9MhR3y3BrmMlULOcr7mxCTuFDzGivMBOe7u/myaUIDMevyC0jbCXR
XuxuDuBrHZRhNEvS2GbBdCPjZ9BnFxhCCEXPdhjhvCyhvnEE4NfreGU1QyGs
uR3dSfn/LwAyts/SiXM84E43riif3v+7rbnkH2AwnmqgQeqYqsB1Q5xRjqL6
rupiDXL0Ar2kn2EoZ5kTierucKTXoROQyNWtU5pYi1Zhi1/dFQ5Vzs/BVFPi
Tk0Ne2S81MX5FD0W6wW4gOhZBlUK10eTXLGblF/MgUNoIpUHqatm/JKpHkrP
owAp63Qig3ipjBWyFOqMQjN/z84RIR/r53641NGEbE8wHW1DHKmflckuyZQ0
N7vStsNqRpzA+eSAbVGUgJe260Qu+Gzidr8z6qj0cAf6NAcWaaEPgRyNFmem
pfte+jc+FZ9hgWF4k59EdPcmMGDYYBuU3mlWgXO6ipLQc8YQN2rFQ7xVbLOE
8Ru168VEeDwhCxK3dw8c+JLZPxsYZLHcprUXJCEreXpQbmrHXVnvMR7Sn5jl
Q9Qd9ZNcFZT5Yo8sNxgaEdzp+16g/aZlEoDShmqu/dSLnWUDqaLGHQPwQKP7
4yU4r0E/Y7H/bt2/6OxN8W0R0oOkXoajUrk3xyitbZ7sRz/NE6JBxTo90gWx
grffQGVuiM8FJysUnR7ss+hbiTyIA8j53ETC+pYYlku7ULRi9O4EBBv4EPFX
e06mA/bvyLOuPdRmZjpwdeoCz/fNV0LtRfklMHMzsgCfpyv3KOyjOhBcHt2s
B6YiXS1H7kctM6HNrw7G+ZsSPKbpmA8DKZNJj3r1wWcj/GWyAvq2WJ2VcArI
pv30FJGu/OXVhkNtsTgFrPbBXN76dgPX9hzViLgUdq8gkUpT8kG/yIxcRnap
g5jrJQX4rzNmP+S2buEnxOJpp3S1sA/ricT26g41xrunMvAxZ6Ir8S0LnFdC
L3FgJX/6OgXs1GuSXbfYDoA1Nu4KrDk/uWssidLOzpGLKS2dhf6VvAhic1De
r7696OnGEFPJgvWyzSMTnawLh4NHi0j174XkANdqdoZtXYaHLnSx8qJPKyI1
psm8C2kSGFlXAIQCDPxygZGCHl464BDY2rC+EkXLe1RBTwVRHFMUHlAtzoP5
4MZIeJqAQyc8kpCHBwo/HPbAIZKwehF6Z0mn/ZAqI/9OKkamBM7yNUD4vZqs
vv2ED+hlloOY5+VpVOOAKw1TxdD57TeIOeAle/o5ki5wzXVeW77/PZvdkYGT
Rec1gZQCS6Sr7baKZGHZPsnLB59aSXcAvrfjUGZz1UwG1jRSXYucajEXor8H
2TwCP/L6qP15QHsoSN9b+AWi1U2HnTQSGmfTy+4tApCOBAV+JQGkWvHO5UG7
94XS4lXQwI5+PebqBCPjX/pAtZ+9fYxXrHWBGoo1cGIxcsFIVDatSvXkxA2M
dQskemuoAENKFXf1CPZyswbaHNfqmpKpwxBhzmK2OBSD512vnhZi0t1r4u5H
MxSHu6U+ThcxJsIFSXI0mdsSk5jrxoQiqpDTCzEg7Da73L4szOpLV4WK7wGP
gde44iDp0Nfw+9pszPVnHV9r+eK6hBq3QsB8j10YyCp0IZr3VrbLgOYFgChA
GsE/cz3SMWNW2AHgfLQx0oKe66llS060SHeO6qPnhBOjj4BEUuvT3SwHwn/I
UKQq70coA5Ui2EZGaaC98K+LLMTkcT/XMDOqLbK9nTKzSHm4qw2BNmAw51oC
PgfLmt/BgJdjCd73qg/xop8gUsdRh9invypI8w3wkbnalh4HFWK9Bq1RptOn
L5Gkc9w75haMZGq1NiVuD6+VsKRnKkKwsB+9awR1jWI7jqMLUqSIBqgEvvFp
xiqmlq1FI9sgdxkyl6VcA7Z2qoOjQXYahbyPedSr4J2T7H9lIxbq/wceTZLT
3vPuRYzh9B386VwZoq2JuasPJIrpCvLT1F0Jvffw/bKVEpM06ialqgwBnWbh
l5gKge0H7o46Hd9XOf0fecHJsQ78G8eSN+Sm6ttJUzBfqs50JXbsHVSEhkiJ
5KHWIda26RunYzMtMasjmr+1p425vNqCWues+eC+4Vd54Zyw63DKNdMvTlWY
8go35fchOOCvFBD0HPTZHS+K3r9TQsu6m3CSYjEjSpaMn5uJDOIT0dDE7pL0
/CTJgMXCoNHHkXpssuNtZI3bwOMBE8Uzd02EkYNQtfZJ7riCzguwO2PB9/pv
I2zl7bQlm5b1yCeTHMTG2o6M+FjyPFX/zNGgJW+XDTxP9Oiil8Z+KojWOyBg
G4/IdUUaADNp7dunsGxMZhEH5K62lKyZF0aMl+/UAhnzBA7Q3JRvF+H3eBi9
8hvGyc+kmbL0CbeUx5qv/BVo8JOKQ3GmcOQ0U8s1ueEXVRnv9yNCFxVtEQ5I
8+M+xSgzdXZ9qJHV/xykuLaYy8FtbHLfrg00ShVTlYutc6UGShILdM4i9dfY
xFQWaP+oPkCQbBKkDc9H393n4a8oiUXeD8VCPA6TJEs+ncAGQdTWwpi77EnM
8h1LSu6kJaTtvqx5hV2N+5KPdQA4yefM3IYi6o40ht80s1R4MEmQJhmhs0dE
Yci5ygSGa7iVUawkcJQZM3jtSgenYEoe9OvG6sHWFchDO5IZV2xhCjN7whxJ
PEyPr5gt9Ft0dA8Y8RtFQycvxwba9JegLtyoWTGM8WHcOzI2O+oXtAJ+jE95
bTBF143KRh1mfv0sRdalvIhIFM+iXjdlLgd3g5tTMrrMjD/wCtmRcobrMJ1h
qQVSU9nWLBNR0UC8A5nnQKB+9vmcshgpRPI+RVI9pmKL0Tbfbk+dTBklyvSm
OPRm/PDWo+Hn6kgIjjMVxB9OvBb1LB7GzjLcHjBSq1fYQpMiAoRVVdaaXwdr
NUTG8craZM72S7IVVEPPtvqDPb3Nc3CXDr4pduIYYOu6qvY9q31uAMWiZX8Y
UWZWmDV5eNFWE9FliAgUK9UsjKdvQ5EVvid1JJTXcGby9R/pzhLCwpn9kXdG
ChsamFpTfTj+a/xU86oMfm+rfiIKzrIubK0fAzQ97Qzalbj0SvzAnddCRvqf
b+fUduqGL2LGQpUjqLxz6n6biohY/KSoGOYAzSu54GXnhkbkUU3R9k8ghb9r
3JKlqO7GsbHDgbIMOSUjZ0K5dkiwkwdLAU9ZWAC7hrQJ38a7iMHJKC7I64ev
zLi1vSft/qvrNB9ADXc3kmlTAEYNxz8wItovbKFFDqg6i4qf+pvQr0BWLvWs
/IdQLRmrNAOd2JCNR01cHRc0jWFyo45/ld+SGhNvp1TE07rh6hmEIgnhq/Vt
9TylxcsJiv+f+uqEcEYgwwJff1RvTtkxWkqqc8LtDk8LqHWkQLMVuv5P2Qt9
lTRz+6eGKZSCndS2i3dbTKGq5Jc2fPFYS4dCqfxTHVREVJA4Goiel3z9nzLX
TbohE7fB9gelzzS3XG8vFvotY1ZnkArD4cspjUxqmyLzc/2+aNA6U194grqj
yMBA0NiYYEdHMgNVpNDLZibjdVxMQj4d7Gl2iDc9HfWQY6kkDC4vkzHrO2Hc
g2C+16CooZ8e9VZOx75D8NZvTykgS5fh6EUCdo9WBtFeOoe746ydby6+xlua
5raZpdf8FHKjQa5GbFnGV8+QwknS+1hd797q/PqBpi88GvkDNFl1Dr1oKjDa
WYSxKSp9k1UeBGnYd+InxBk0jyotKhJStRacqSM6VeIKUEnaEC3fA2TzJvJS
lLtaEuxKE2riibMKvANefn3MnlyB2x6i1Smar1+q04/N3h/WvU3P2QAl30FL
JcB4GzYb+8pB1BiA20h4JK5vUI4b4QRDgvGJOs/CSMS9T3WK+9vXQuDTvOpG
IXS1TGDCBiLH6B89J6XIx8w6n9jpVS0vqwp+dfBEbTnZE4Wsc+St2+ooHwr5
KHfXV33h+RnbJhZkkf7UDAiZVr5EB5uHIcJxNkiu9QvZkzYx8lo58Op77gOg
9zuUoMTXV+oMa7JEHzyPjwAWS+mbbWWQAqVwVKn3LTZmfAtcmflsTu02KAKg
Iy3IJipUlj1uXwWKNG1k54j+kDtxTW4A2wtwIoEi5TYhYgMdB/IeKAnP4eqJ
8o37kkx5USGgxxLWWC/s15v/6S5T46giNikeLGYjfNB15aRJKs0MR0A8A6yl
Fl5qOTwjzsTffyErReYDZASR6/c1dvQMsFHbS+PdDuwieQ8wqRfBuduqnZwo
Bez0UW/DfVowvdQvF7JF8rUl+TK9DAH+ElFA2iIFfUz9cQHL1IxNdLJym92N
bZ04tYFV0z34gObmznC92h1kYfKZ59d2FZd/HwSDmigiV0zViPXP9DHjExAw
MkLl17Iq3nPWeLB7+Rc+2+YAsQUUVCNBTjX3Su3hHgIU9OyltFFIlSQHe4hu
dhEIXI98MElOLctJhXcMKuaOcsPrOxDVcXvumvL33Daq04KBcdHPNL8rHw2s
A4cP8yDNYcMiIsA+BB/h+0uAgoAWNwXaJbRvktUk9i72J+AasTDKxORpuBLU
bdptiii1Qp9ZWUbaVC+Ys62qLEa7zHwIYGMRo0MDL+3mcCxnBFg1xYEkIxCy
N/0kg+dCwZKser3R1bqwJwpFTc54PItHqjjxjNv8u+zTY2vM2MP6uKEv6t/D
4wlcEd9dA5GfNfeg5guoU5PR2LbLuDTPQEksPokKM1jvBalXt1UA7dV2hDh0
zcvKnfweRbO6wFsiq+SIDwJrzfcMWAIGCPH9B5dV9T8iIP+KsZG7gNNRWk+E
R5jOHTI6I3SLFYWF9kgT1rnDrP/wJEfT8C1q+rBIhucd186NpBBXG6EzbwI9
DZ5cFYOhVZJP9cR5BCz7UbW5eldRqCd+o8r2vqkAgiaz6O8AVzAJY3x2MFbg
9J6AD4ZXVQYT/v6CI7e5xWr0k5pVliD7RWzozfsxPvG2evpSRpPG64kex/9/
gDTCANuZp+Cpf8811wIEX2wGcZeBbLQyL4Jqpo8QnbFl8G2Y+liSaWbJ62Y2
6tmKGmb3rW7oMM94GzDtwcRWKzxsWCCHeBJe4eiVlM5E2B8ldy9vNNAGpOQ6
Bc5u0qtiNm4dzYSreBWik2zP7eUs3iHJtsdQjjK0JcrEtb2bVapwUSlOCjns
SyieR3yMCk9MKniX3GiL2fUch07x8QX7m8qYD0IJ9n8290rIfDDCTalk0iEw
xJaKWh2R3E0rA3I0Mi+qADivhFrQKwpkDp2sMQK0gwk7pbz/xs+igTki7sxo
ApOH8JEVXGD5tKABhgOGAFdVOyOK6Pc5fWhq+1sSVHzwg5qNVqHVD8dm46di
oFZd8sdxNApuxy6AXbifk+EtbrA5wfhCYj3xqozsdjwrD+/pV5wbmU2Y53sl
p3pPxV6fr/q6/CuXJm/W5gClYSMuy5F3HtGTMKxYIS0Ian//syQcx24c7x2N
guFwwbkYLQkUL2gRquEw0vvblVkGkBmrpk7R5mx+7ckGw71fKeGttQHadVcr
ARLKr6lFTEJ3FEu8ycUDXfF8Unh5REIprR955eqlZ6zCw69VOw4Od72BQzf7
XLoJExzTD22OE/XfTDaycrBTsbuYLbmzUnZivWWIRWPjLh+GLlj3H9+iyP22
9aVLm0h8Lv6EOiOsqofJ/LhQD77T3z/4vZVPTfMMPhT4EbFBR+l6uIYZd1yq
OhjXbj9jfMopnQ7EPANTI8HXBEq5BBCQI/owtK0MFndRSzOditcZRBOK9Xz/
KDrzVaV60/mnu9fUNNFz3EgyVyvXrlaDPWlH/z447eY5XwK349NS0lByeNhu
nb4VSWzNS5dn32hoOpyLOUTu7jTHBzzpDnLXkffuQgfmgdpCtB61HMG3ECvI
/eanpuQpROjluHm6d+u/FwsakA4J9LcyUd+A70/GUSXc4TKoWoChVkume3Uj
kbwIZheZq5FuFT5so9nhWzLuUtJf8m9KGgERJLHq6U023w9oO+Cdmz/U+ff6
po6tYBTgFuOcani+ZOEV+UG/m9OB0itRC/H/F2iU8MJ0nkyf8p8Ujo4Uf8a2
gHq90QJrUFECTl97OBgxwECXoXIID4425Ye7zyY85GKb69zzTLqHI3b9AekK
g1S1wr/xtMSQFE4ff/1TiyVAeWDxwPb3EXTL+RJOLALEb9rL2MatSjGWeSUk
dlfTNVuOtlj/8QyJBfXrqlX074ZRU/4iSoMEVO8Cr5iY1gu8x09NSoht7OGj
HJq46BikKGQ0BlLWnaiOOUkJ5QT1GWWXGq7rSY/vSuQnNGp0r+s+Cj5lnlTs
5y0+fKyVk6Yh2EaAb9yA+oa29BHA4Gq2Lt5VxA8Bgor1HPrXXBY0bh4Zx7zy
41AuMxq3gsxU3CB1OaD6UNGqIO1qlarLNM7Qpfn0DOil+VBm4icVQwbkMxHV
rDJ9v+bmeBn1I0j6qkTrn3hZUsFjkH3FSgtVOSTooCBue5R3cR+YJyQBj0W+
8CkIRRkpISORIJLLNTfEAyNiqAL18Oq4sML7Yp7wT0ffo4a1DClYVqIS9k6O
H4xyaPzdy7Owb6fcc9py1U6kVaOA0FBOGf+EP62BDBEJGL8bWMUVt+oBHrkn
45kIPuW83GQch1FwgKfzbugTYXgqKjcm2ynU+Uy3Pd9u9DvecCi5EdOlwLXb
XxbbZ9q7q6p1Nvb4Pg0JM8e4dY0LTdeXynhcwa42soLDi+KPlo0o2NlRD6Wr
d000q9R8qgvz6G3DRKUzURG5kuRA5h8MfoSDJxRZrP9uWAgunMluOqRi37e2
c4GPeEjtgozew7uU9KgqDVYChoHvWn1YBGESVzVa2lnMVAfqUVta5HBplbHt
N4w/rsLtcPo0jY/TnCcrhkD2myLFSaUSube8O7pKo7mWOlbxt0syfryrwqCe
K+Ye7t+UOnOo5YSuHkerTuA2SgDc7GOjvnmPvIZ93G8kfvjUFpTy63T+cIif
s6qRYCw+uITmqZK1PxhIim5Ry/qRVF6tuPa/61kYxZttmJcGRBM42JyR96dI
iwCuNOM3j85z8E/QYT2PV8O/sisYLtkL7gwJptirv2Dj2gB7Eu5EyYo79VAl
zjAlJRcs+wkwiz9s3efQ6WeajU6a0Fzve+f5GSi00J7im/M0+ItSRaFle64W
vnmrw0Eep/YkkDVOe9treWcN92jPu0FSsLHiza9f5o683ZIIMVT0hj1qAtS0
x3vtyqR9MxAr6Srqyt5wdJAhgo2xElbtENft1/rI01qW64BEgTRbPxEgc+A7
FD/k9qWv0UW24p9f3C7ar5wlX3QssWQX0ulwvwP40LQMBqHxgbjrLumRx4Nv
k4h5+9SNL0cw3wH7Pn53X+X9X801mDVHTFl2xvQ4JQKXj9FnpSSfMs+bvK1o
oog8rcb5L2hQq2kEbWTz627cTec3Pt/PLMdd7KiD1egf46DgJcKgP3NrBwyR
S+YTRMmC720cG6j7688G037/uxXWFkCX4zchXm09Qhzz8mK3YyUL8u2sxrmG
5zWs41DMftTOHHc/E1Mhtyngwf159L4/SErBhRLlYglTh6ouxs8HPhOmGtYA
lneQPZW13vYKvpU38ljaKLMzjOF/r/C6B+bWXXzLS4YCKh0QNUHrW17+rSyJ
YGqNpFg1JEuWloEaA7x7TLuarn20s+5RUQzYdh49DLcAJqeQk8wK8sb88Kz1
VIrZ3YS5vaJPv43B4InNDfeiBCCIyzj3llJtXgoHCZtoA8BBoESZOAHBTPen
ngAr8C5Od4mrao3WT8Ab3KeDOReL8i/xedWfiT8qcpYJZcB2gyh9tObcO0en
/g2sB8nz2QJKAyg3Fo9rOsJ7h/qK7XqJ99Herh9+WiYcs+TxzzO5Hgxprob0
RyklJmnz6GhT0S0qvxRtiVNmBbg0b9oKDMBT51UQNRen5PB8P6jMjrNNVYWS
SFsNgnVrbyuAu6bOx0+osXp7llU+1Fy0Ba5QAMyV3udmmThWN1cZwJ6zhtn3
FAUj26mIpizTqKIRU3EcJhWXfGRrRVkAfjL6mL89D46x4Gq9RhHqfsOd3Dtr
FdyrLZD00Nh0USxyS+on2oGLVntLNsfuO/gft2MxbgCZhcCwi7qojtQtDYJr
HlWv6S00xmIyEo7V6Lfy238zwH6vUjuIChnoLmTLa8c9o9i5NOiGLysvwgWd
YERtEvkQZHY9BZIqhBIrCrG1qg/vJqO42MnbCxlytySpoO019l4urN7MlJOu
n/sCste3r/hs70oMxnmXNz3P/Jeh8KrGERfsnRHLNX+BduQnyhIjPkh1Ojud
EDVQc7uycDWY8fyyCYlLivpJ93NnRiGlfsDs0Fm21HABHUT396GNw9wGzb5N
a97TZr21m+lh3aLefCKNMw06yKnqK+6yeS0ZAdMJ+X5CzoQGn7a1HCP4QlZq
ecEUfNPJsofwW0WEXdF8I1QOQfabX3WWFBR3HkgqIpAacuC8awTuvcZrJjTu
WKbvqB04I02axHgfQBqqKgs8N/eZJZr9ShSJH8tYQt1ZpmxOvqu3qInmjXQh
zU/i4eoUo7rWIL4iOC4N9l5RiHfCg0YOfSEgx+mOK53JOd5K90U2tvSpwshU
koaEKh8HslIMvTKXrTZpY79m1NOuYWTfORclR0OFvtfSBJNIMmbrp0ZgrEcy
fvlM/fjcTfgvIeyCY76ezroMJbYXiQBMtG9xk9rMh+Xdcb2fvPjubbicv1Le
Y/kvrAwqby4YIFV+RTrOafhYfi6ROzeqqfyB1+2AOYD5QBh1ng1RDK3LlFnn
ovC/U9reNEcHdP7gDAp+9rf0GRoK84N8eVzr+ueZR9EmuiLzAdVUjnjPGe44
iUKaKL19+SdKjK5P8t83XcjSfceYeJII9CihdfIB03gbIV6E9XyrYx+WvsWv
fiuu/g70Jz5TsswJU1Gj0bfrvuDX2mkHRwM9LGD8OEneLUsxFZijJB1RrgA4
yE+ycGwt+D0EYChu1Y0StcBhOFMG/QBcCNGBDiBYCtYRO85m8/mcX/1iYrYe
HRMXr9ZauBCIayLmG2QHefMs2d+pdXl+TGgT9+bCYRM3PXkt2+SlZDX4pS/b
RDJfM+FKrBlE+I7k68WfpcKNpImllcXoKezum1IrpiIsid3szZtOBhrQ5RxV
H5MWZM8lUhmzUOdrWS+YLG/tfPEFqdTu20r/JbQ7ZwNWbG/PQgboLTitjm57
nS80TPa3icBOa2Y06P2gmtvaiyYOKw5Iaqqhlwj5+GYUtNM89JMC4Yu8kc1h
nLzp7tApnkvcQ/DKF/N5ROQQ0NrHC1tX03q4ZhT208dzM8z4oRHvXzK/2CPp
IMyRUkYTY93bUXegmYuTHRJei3V4ffWi+FoxjJ/+mZ2RS4Ge0poBFc/3wVXU
1W5Zw8IeMjhcO5Rq/Ia3rwBMa3mr1kiIs7gK33wiZ76X2uUDByWHcVbvJEuA
BGHumPOCBJdydKaxduboglU1CxItgCC0wujXihAwgORxVVQC9KN1SIMg3lrS
9EqwVWB/0FdyO+Bgr123IEHV5JUnRNbDnEGmG2w2K5cDBb2NcJGCCdEXlRVi
f2iY3CaZrtZ6IfnaYH2J4k4OTTs4gsaxYkHw5MfheK4fNOqQ8kiQULDgcErp
YRTX8c4FlD6oihdWFr5IQ9TkLEywrVhnbet/oFLIpuHVLQpSW3wj+2hkLo12
IH1HIFQe3fnv/JH9X99KRJe+kuilgeuCOkeGw19nWW95WM/8JR+655y+w7VR
gvxBXsMynTU2oHQzHH8YPUrNl7a8D7iNp8c2AnNCe6W+4yUOjHLhgozAeItu
QlbFcwX6mqnZBHaSnR6ewpS3HtF6mBHKqoB6UpFf5Me+05KQLTUtfqEIXmnd
L/Y5CTwixoXTnTDW9gNDU7nf7cSNXhfMrekX6ax1HvjMlE08E+I3l7il8J+s
hw3RBxA2cSn2DYBmAsosjolrU3TSrI7zX8x9vWVnBsWNI/TiuxH8CJdX28yI
WU2Kcd58bHd2uK7XKJEFB4G4DlAAzmK00EmSNJFFTCjvxDQI0lNzLYZujlij
QalEFqUPabZf7Olxx+nhnJvK22xr3GEOYEOmARmr1F16ga/i/5CYysbMXKdR
bmTpUxjyufmCeZwDB9G9nhaZchhfsdjF5hbsuav6mtRVvmMotAUyAZB4i8LU
JC7hC2exTGlKQrsJXiNqiFwZNhIZUhUamlKg39BT3zfkBEYpQi++Pp9QiRs/
yC6Br6ABBBzypJO4V07G+aT0UsvPMKGD7honulCnk6nldbOwfm8TEX2xZAWF
hKFPAyzMuTon/S87RoCqHWpYAqQkQOyWaQhLuBQ83Ygwpr/SSusRSgimhI6x
HFi9M0LTuI9ojoG562n8YAnY/zV2dPygd9lMIAj2RNcbgoPeWeXqqBAxcf66
Ev+DfIpGJx32P1NJa0Kjs4NeKuz9UcEIDnMae9T5Hzl7PWUslU7FIy+lrJ4y
Mk2vpH4QhDX0niro5wX3E4D0k4cFZmvEw/QS7+/l8d8ydPE32o11dZJPUeHF
vBOkn71AY0WChMC/dtbzPoQ9he+Nol1pj0V8yfpJdRyze43qkGq3P/lMBJct
sI4eqEXkRxBcuv495FqGdqeKQcUztb+kbt85WZmV4oolka2w/7v5WP9paU/+
7GUWbTqMFDrbtjzBLZ6e2u3N1zmkL2CzR4zr8yhjH77dlx5Db3TpsjEw/OZ/
EMgxhrU1psyIKkDZt6s5ABqG228I9+P5RQc/KI6MzDHBpF0f1veWclLehd2h
56jJ3VRLDfa4CvOk7qDC/OxlatCikSVJbll3JIbIBFsKiVR7v68ORoTMXRrw
FTalEd1G31gS+dozJpIAJCv2bKn1pdm2elkMmXr3lMjIsU3eVBs3xqJmyTOY
aiALCmGlz6RjIWp0QhETeQ6mT8Bbbsrh+D6koj2GHb+xw3J9ayzIfyx1aY99
X0Q/RhVZux3QANqMqvMlbEvOsJvPR55ow0xXZJr4R78nZ5O+hU2kC08iMGtm
oATEy59a1u8DHygDSUre3lwT05mZVvoqK0PfFeaU3gJa5e2usOE1LSgXRz3h
yu26wNx82YJBb91O+GQewJW9mdi5Uprk48Dh65UGMIPah88M75FWEnMTkriT
HmhJTQWC4ah6KWKGyhl52qgvzCITfPVyYEH3dmvVK7ITGGFVwMA+KnRM3SLZ
ViKhaVqizpvGnFbnrc+fqsHlEvU19tmAb45e3u2icGnxqoQBM0SRYR6FqCYH
Ghhkvla660KGM9OFYR39nWscbTaT8q2+aCltwSnBhmRXk/8Ou2wwq1ICZm9/
svTN8EfJuOYTZtNlaoKvan3cUgBdoqRQLz2M77T47imaF3gjjuNA/TwhF6Uj
tk3oVXuMH4AJ8ggk1FbXCt8QGwwsX5rg4XgkNgvjuGnhuF2PA+yUsT1N7J7L
vDlWNf4joy+0yx1VcioT+jIS1/EMGv416ZL8ClQlSkDDo/iqQoHUXMR//Sl1
LQbdt1LJUPOsHmJYgHxc2rUZtPR1OgT6MXUDdm2WgO6AM8ba4wV3fac0jEkr
o8UZxYElhrg/JKoDvzMBR/jnjpouirB9AHT10blF3vIp8KlgNMkV0NIP1vHi
dFLQHTIw4eRH/O344NcRNl6EwbBYNHKEprd6fsoyl9HvUVx4pmPfYIIjj/cQ
XJTgw6t182q1wWG5iS18DcjOUC6bvErmUFo43Obc11IwdpeDnAHF9iZfPPH2
+cH6is+P2qbbFb53Tx6MwttkVcjFkDKfwVljmZgg41whKjcGJV6IMQ2fbN4o
WODMqnSjL0ybn2GnitUdYhhIth+eAhTMt9KjEoPPyyPxRrZnJtIKeU6FSBuV
I+wpxWp8Bfwkpxy4LxeswpnBeRoiqoiNZGEMyCK/9q8Zzz+nnQueB2HcW4Oq
yTO5ZKfmfjzibAyChBCkueSNQFfqIlupMaLnae5F3tN+nntlsoh0JoeH5wYB
T4hPVIDo0nS5roJ9/Z9WgUhwlpPbQ8b414HOXBPOMJwR/7IoDsYRRft2S/Qp
LvTaKQj9Li6AgT92J9jIiXWOiJl/tMLcI+6ZlRppTEKRHT0kjR5SkS/CUObm
wBegShXdR5CMkEB06j2/9Q7ubv8F9Jtt8Iis1MFNS9rhXDefOFcINmVubJFt
sJ8SbxipHPac8doEFnZxL2+khTMPKuUp9E514ZeJs2k9yNKoLSSWtfYHToBC
q5O5kjqq1jYSTYIH2UiGrkFWeqvJdS2zYrK9n3QMPCWtgn6ys2unB1umDX9X
Zb6hKXFDDQU7a6ngPPlkQsTuVhFzttaxJ8PiKJ4HF2sSVUotCykDEPFDRZIa
nO0pr7NbBuHpQxbRp4gtHehrUJWVCfCCiCjbclDp8qvJniueooPx63IkNvz0
f1ZXrQfvIE3Y5GS6IJjXPI/sAFlR83uiogJoycXBq78waT9QXsIodTmyqjon
M+UbxNPQbyMJfUWq1pYjHnVV/pAIAzucFP2smfiXXwCnCykOPQXJGEzJv/BA
Yd5IPARVXvV88HsTeLlyPAOg3Y7iLFAggvS7A3BA8Bl3cMKw7LyFJfanwtFV
v14FvCpMeGHVPO+D3qWWQ+JeBTCP67B07SzEi68+ZNtwduuP1MqdPh8W1wrf
2Vq0OMYVovxfLHY68HcWQNPuc4tbXia1u9bJFOmJk4Aa/ftXEgjhtfRzrwZx
VIGHbV0PModPhn8Ze7zzzWnkTaBN9hBLqgVjLHJmXMcit7uNZPBe4rkRwhQO
8k9ESqumtrOEl0iaSTUmD7M7ZHPPBBVHrLQ3ULQDjJCqOMyvcEi0mMPPvjlU
YJGG7RMAzTptBcPmDIVxwlFBJmC+P24wUpnQJxXWTcYbUiUeq9PNaCV2NhZM
sfFOrDj7RWLuF6TC4GC/mGex/JODwEBaxXmHFrbcS4I2/MpXjwY6JUxuIzEs
FiCEMuY7mPxjsXYOe4P9PRXwqZklIhN8TYTM8F9bo/H8DmWUSdTfa8QvuPII
WGKPaJJAOKTzEwilBeCstsWUby2IwS+PaeHJeDuUQQuIcGDDP1lBv2CHei5M
0E+edMCGlA08BadWstY3+8S8Fx10pJRchjZbAjbFxpseorH9+3Idg2NF550r
fgemhOqMMEAM7vOoinzRv5gIj6Q4ChV5004MuX0WQf8RKsn1n+WMPm/JZL9m
u5sMg23J/N95W4BYa3VbAcb0uBDkvRo1R5awOKWUwPyUomKq62mI9kGsxphB
l5zVRW1r3IaUVXrK24NvuGDw1Jui2I6j6GIeNAb+vVBjjSKxctKOkcRxpcgi
kL6jRNRTaWLUGiqB345mDBeZjg2p3Dwy0ZkFPUffQwSSFSYmVnO5VYfyJVMv
Isf5m9/JsVoCipzmoa9j2tgDX8M7Iu/ypPX2zN17arzoy4cJI0tnFZPfQ1T3
KIIsN9fBkGkFnBAZvEMsNXxENkanw8OeEKmHVHxI3CqKyeAyaeOjYxhLfvb2
jNqyiJaUiSo1VVVPGsC9QYmk4Iesk229eOLIfM32tZQhxroWBx/jevHIBbXT
5LZN1gjU2QLTEVpKw3kZ0w5JAIBF3rnVc2kdgIyXF4GaxTcUL09VymHkMNRC
AHBQJ209196EjuxtkCT3bFIWtlpJy/nGf4ywpaxGCvQtdr3PS8GdYK526wf+
1eiVqBQZx0Jjyppwf6vgVRuodoWBRBxXP1mRVamB6MrTJBlLkfyyu6984+Lg
CzS8lRs5rMgF6411DCC5aI4Khn5wxvIeWLFj71boqJK6w1eLdzDb3XnAn1jF
R/ywKodSsM9k0Hn7Hu8Tyq7MTQJjHSOTLjhMaE10TNLoiSASI21UZc4TF4SO
x+0ELa5T5jtFPHHOtm3L8TaZlhU/Tj8U0fE1ardbJTQnL5g1ku7yZPMJRGOo
TYIPrMxrD/MHb8IymO5hmwrJnK/nmzIqHxJNHyQ5jCC4h3p+G+Om9Z+POjkC
Gx+y+0Z35dpDFyIXDbkyKGTbSrE686Hh3WviXEfwTxvZYaDwmpaowOT8qpJd
S2CZ11f3kmmpEA1oWoghHplsyhd5M0FDmKPC+sxQXnGw35etV9z5C0Dh/c1A
mKNU5ynJ0gFyDCwPfUyFyNCvhyLK2OiZMsCEFCGzFCfxinSGrMqAy1CBr/21
MPwEjixTypkuZHWIFB+nTrxyBEe9pVeIBuS2Da1kLMKraCaF6ut2iTqzgK44
z/sMd4ZRI8iz8r3gJ/RWx1tguKxXEC6K+RVcN5L02oaiMNWljxwIjHPdKkEn
/38FbEEJLHewejLOSGu43Z/M6R3ncPANi3j6P+Eu4D/LeYCFw9z2K5kifMfo
Rsl6G6EqPv+AMxTqxmCzTz9dndG5jhkl86MRu72n5Ia3ynf31zYGQPKPcIAK
NyO2aUm8cGmEeqKWfv5s2NCPGooxjdgNHI9g4z9arOC0Ph5VUzPcBHSfnO3F
PIbn6Y30Oem5/c/tqsdZ41/QCyb076gUD9xU26yAZsXZAIV5ixl15BKwrAkp
3SDCI83Nyn50Kd/lYRyGTU09szMZng8VjB5RcuIURpunF8DwxzQCj9qoWwlE
GX8nqUXoVt+7lA8ipS+C6ps4DA1UooKhA3UWtwR1TZbZofz2j2VaURBvqdnW
V/B10YwRFDmGZ4a0yOD7qCoRKKo13KRPCfub/VWSEKjXgngujTlsVKaAIm4G
knHdx57X7M2TpvER6INUPldNLTBW3XeJ8MKqKj8zxndcskYG3SfHomoGT7mH
utMT6pX7WPpDrXPoItHCA51uTVZGKiSXUJgK+m7hsw5VFricNibHeDpABTyo
NBV4IV9oIe7/vhaySS98erJpEVjlJbRt3lrnUTAcQ89acqeA2cWM8suU2Jzk
qOnsllyCEKz1l+rfQXOizqeAOIh5qZCCZ9c/ER4BcNWBa+yqJ9TCR/u2EI5Q
G/wJqnf2YLR96OvMsUMCcTR8GzlwLpBUImKZFhemgXhJsXQKpo35Daj17zv0
p1TS3odpxVe66OHt8af9NMMhAt5+KtKZV/fXL+US1SJiga1M8eGH4XqYvKgq
cTVYjvIKsMzLdJNge4Wzem1vzu36QPj1xubWLrZGxf5nTzqIYdEty7YER/xs
rUXxHAvo7l6UmC1AX/YyVIaunlnMuk9A4sZ6EU5QXB4+WJdyw8z0DiGZkGjE
g8q7NTeghFNUSFUzoJ/tw6epntJZZIGFEz9I3rluJwXWGn7CELIpJdm7chPa
TVijZh1kWDB9iB3ex6GM8zdc830ewOOmPj6hmBq2V3yLPwSjXXiJdI3QYguY
ad+vdrigusYKeIMj7bJZbsTiUkHAqVbMk/GmonP2nz9AI05hpp0l1UGCN49V
M/hGJwJcm/lmkvxLGbHRoLvJ2mgQNPLITwQojGwxH/ZArbh4rp2V0xIwM5ck
lEqdKRHuHbND3HPIK8PYFWYroPz4eXZRcqbP1TrVzkcXvF216ajhQ48tJV3F
00nO3GJVwd/XlfZj2O79i0bMZOfrbVLk51YDuI+awZzNoiZQ4bVPHZEti6Us
6lPkU3MnXoDkiK+MKBQPz6XFz9XcnROUM5iM6+i7FjQh5WO4TsNtYzQAb9a0
xBI98ZH16OvBlxTMJeJOBGt6Y6uRKwCTppM+DUk3iRn6R3uMNSGIobpLbNQB
rEUm7RZbd2TN2wvb+Nl7R+7jQ6T0flZeZ2TTmDB8kZLOxSAI47xxW4odVmIg
ldDOFGOJpuIK6avyER7AWmrXJ8QLIDRpMCbfWny3ovLiOuJ0kjIbaDGj+y7w
gYul2eiiKoJNTdwJedFmWnC8KY7gomG1PMuP+Rd5PQcYxnt6ovGAQQImkVbw
MtwOb+Ab8PzIaCXMb8OjOgcFa1x65iBqWRfz2nnxO0TF/R5NtskyGHi4maTc
g0M+F4R3bCQ7nEgH59obbZB+WrGNtgOBKtl05jM/7fKF1ry9899xlxdYmehp
8IwyGL3Iqn8lZsLAt19FkZILLHNcDWo/TwxVayUk7n7qbogn3Wa54s8uuvX8
y95RalEs+WTyBIQpN/RtBIPH65QL46wQBktk6vTcEb37aZMV5u6dQi0Eezh5
r7FFM/I8awkYwxtAVh0VXlUPd8IyHllXt0SYh6Ol+X2CArgGXArzB4oOcXXf
fh431Q9wWenZKfWHPi5xDMcmt8TXBm/HsQ31cMHERueFTA2ukjc1XZ6wCfyG
LpDHPe94LZ2CObg3Iwu0VVnYvz8HraPYnHRLNz0p4fsZQ7lMos1sLwLfpOXR
Avv9KACu1X4Ukcgk6rQRb0bj0E9P+4AT5BPC5xYZQdqhTvhlNfJexpmKP3QZ
FC1kJK1jrUmUoxit+b+H11umCdjiRQnrYsYpiQLf+uTswLCHEbOasZSFTEvJ
50LhFo7qZ72FCoGWNVgoil1A7tYpEjN5ik0posnRD8aB5Y32JaJd0bAjJy8U
sDjBqSL3eAcmQIz2m5JSWePnFB0Vj3jPXE1EkAbRXUM0Lj0n0xgT81PGTTqV
+HXgNmj/LcFbOm7THtDvKBfA+4DMmGzkTAJNyomuKyd9Z43K2D4BfQk7hU3p
VfyZoJ7TE8yZ1n1dGjyRdtzhVNAnveXhGscavHc5+zeyK9itFOgcopszijKf
dhVGTQ6qwaED16bTxBpYKFuyAH+U9nYu94VVcsEqMR6LQFrZFqIUhxgVziY4
GCY9tdEbcisOnsf1uVv7HP2jb2am7HwXJd1w9NcZToS82qi2Biczhwc94JsO
R7HxNO8Yo/MRt1pyVu9ckf3WGXMpa4ywUrbrWyNwAZbdX1uaZTlgEBnlR9Qf
Nul6c68Ak4ahAO/tJP1g4LCaq0vo8sLkjToQAZTtASgg+Jlwmn73z4OYNH86
kS8usK14lwNHk4gsgG/lW6tbDZtqhtixHH1cHB7S12IHmeRxC+qyKtb3V53G
79XMpkMkQbJvN2IvHkuHXhYYPkOoe6ghWSC2T+QRHhjzbT8K0ahjCaGiQIzo
SpnCGvul/3owdJ7v9lypbhIncRxpt4SQ82fCaXrpxgwMjeYUH0K7BoRk07G1
I5UM3qT6ibfldzFk2BFc+eg9Fre+IivA+ZWEk/UsV+EUFQkmOW05bXS8NCYE
mfDxL4RbAOnfBftAXWropiU6qxufmnmwGTyGv9buplgV1Po9cNCy/vLu+Geb
lugdLk+1hVUVG33Vc3n8fmXgxVP7zgMzGuWjpARN6F8VKiQjaS4/XG+Rb+dJ
86CTvU0eDQzfud8lJ8A1Hm4Mt9r8NOCdmBRu4s96oMMN7LF3Zp6G2tUVP6Iu
Yfmk7s6jDAATqVTC9zi6jd+9kYJcW5YEfiJs5s7d/Yscy7KCGg0wzCK4TSVv
fO4ttIEUUQdMkj3zHQ4gA3zF4BZsu0+gTCTT33VvBqVIq7bPOFsSVeDhKkKN
DLipRO47KIxmh3I3zbzaIdvFDoxrapytPWu5iteyiI58KrZbCu1l7Vp/rwrO
zyY/Wa2oKS65kkPYbEXjM0vHRwqzj38HPO03/sMOOXIsNrzHiBeNuFgSYgCK
MmcoU1b+RQX9FMFD4paZCmvOM8cW2R8Mgf2+FHccpW3cY1Ai5GemUp2sbuPz
XOXJCCF/ihdIZu1Oi9wK3TT9gHzbKl4WmFbss3aAuvkcTNDiRFVpqRqquz0g
IR3Ucno++o34KtoPprsIW/OnofvT0bMO150GRZdhfvm4aheOPHV8UF4KAGFe
W4/DSteApLi37OSUE2Ni27oFPzuzUpam0dm//Nxt4lAEo5ICaoi5NVj8LUn2
LDmEMGp629WmOcfqvYCsHbnMrchJST9bNMLqGdeAjPAHLCPpM099DqDgsr24
lIIGRPixnmQRMjOdwOiPwEJODnr9tEiNYDFo9rKIymcqVbF5mU7QPT5FvbrJ
fFksZ5c1MIfgQSenpjFFa+RK3EGNdyjcnolCS3lUlcoqwUazNnEbvGefOr0Z
7hMTKdFljqNCbtptJ4iaBw4xR+iE6oaR+LuQnhj3mycVy0PzwiKGSQiViF43
WXYJcmgrnOXWkbCzl8hWotlxDHhXWiH80vC/T3hVfvvHrJxuWVWbxCIGHr8b
AeHNvaAcF1NIQYwdAMB5KnQza+uv2FNIDVbT9LFxRdfccbT3JQ6yyV0pN4qx
+fz+SdXRzirBFjKbys0W6/SKWryShlD6t9nfwyAp94jpEnKXhmxW5AeXnVzU
e2oLl67x73l5A+3BB2BizW2E6hSrp9MSlMOAdjPCTw12p0GAPh997XtdL2VL
fbpJ1uCGD1eJD4ZuWKxFKwo/Ks44R+9sLLMhYp550iKBWiWVwP5kqePa5RCa
517QhANIHMKZ5luUIjR3GRdXzO9QA7ntoIK8D2oKxIZ/Ee4DA7f4DXZY3L5H
wDS5KzZ7pqlf71PbtiP2SInwtOT7TMEOikTx1fiMsjzZv3qALnhM0QM2k78u
bhI/1TS5J8tHca1gFaORDSlGphzSM8Ho2cRez1Wjta4YxjLINYujUY9Vfk4k
xO75ucRb8Vry3ep4MfDmxjhEjXHZCEcSlaNdP7IwZuryWpCGwnpgZ6ApJLcV
wFFSSIK7zGp+1pAbPXwhRg53bEKMSGcs+kUR5lRf3wVK3Hdy0g3qvX+DwJe5
sUIkZ+a68EG5er4YEZ0K0JN+g5w9TQr0U2iyByhoVZQjvL+3L09r3i0MMaaY
9Jb6zMipzObMb/3EZ3rAMtPOCe6u8tTC49tOJ8ih4Bn7v9JwYUaWyAmX6vJ7
7b0/bqBk4M1noBR8N1qmY4kbEB3EdkM6ZXC4cYWIv09bpAlfsBIr4nJAwXZn
7ichD6zQwreyz2hwRmbH1bgDrhihKrzxIhDIcH+TbVbx90p+p4FbM9ttjgNQ
UxbdXTPWET/5SdhEc4yMeYSDrMm7l+yaQ4/pWvbCJ3kPfetJQRhYuAHN4e0A
y2Pev8fbXkqxMrwbPfycVDQtj21/xB3Ix3G3A8o8EaUGj+pU38PbQL3ggz84
1ZzL9SWjvTLbMK5yPfp0SnyLcrfFBYLrj49PyFoKMpQC9c2Re5oHEgdB6uLO
9ky3l6yIOl8rd8nc6lU+6YA+5jLFEjNeN6esVbTEUonAewZvSbpNw6kXaUQj
EfOKP9CuQpQy9/W1Kf7sUUvDmzn39p+QQgAuBtUR/Luh8j4PbxuVIrWWfnwH
bNKy2otP1tEctpZk04Jde7pSjQkdLaqqoFqrBcawCol+W0stmzA8FXA5h6xH
YK8Wy5cQUC2qwBDlop5hMac4pBy6lzRi4HZEZTUCWeI7/foOZMs8RNzM8ptI
fgp3YQF4EPT0iSVe9kZWUT/tV5KEdLyTA6OyhHIMgG/aaU7EYKRYLhMqeGEz
ubv5KUW7ErOEdk2MlWBIbeWQPEjFfFmjbc6hO0yqESCraL2ir4NvnKhdeoUf
F/MCwCozfiQTY6LRoDHku1wrI0Yl/ovNsLMzqMIuoXoFnZbEF1i6SynnpS7C
KVGV3oyKZNsbcsc9wOmkAoBq5Pe3It+cEn7yQMFGH7qa1GpUv0kYmyLs+rRD
YVJS/yq5RCMsX6BfHwyvqeGWloC/khdOwB+Y5nTP8h9/U0NoSnuCyHltJox3
IsVWTvKnBNrEuHASqLq869BXIUxUDpYGiu0IFH8ydK8lJJuEF2daf/8K7LLs
m6qyHSGFmj4O6gLe0rLSv3KearHxCgvRVGdyGpADNYK1buZxhES95QMkWMC6
Tit1aAz/YVq9/2amkWBGaGsIFEyTTSKbks3at9977Jcb2Qde20HKZ3Klc79h
DzTU37Y2qlRmadFqCIrYnYu6Y01ieejxIHr2aZIxBIfT8McKxQkLlkQaKctB
t3smZZBuWjLBr/P88CAso8SS6CITvH/y/3HW9NJykaX8Ll0LYSvyALyRgwSt
FqCLjqC9JRw6s7p3KOd+/M0kHCkwdPlXRKwZbx1qKmlFbTr7qbBSfcvQB6OZ
Xhx7ag3S4iGjFwDXI05cnYjkP78vdYKB8JHeA2IjTEk1zPox/jRWSucvmLjq
y24B2i6BGkfDWJS65XSN2ATBv6HqrpWg8uMydhbgVDgS3FA7wO7m3pIsFCLa
ZAZlMO0lABlguxjYDlGRvOuCDDv4XfJ6BEwYrBsGfzl8ybVxMbkadq2rzaIs
lk2Wlr6d9WrftJu6Lit45sbm680OJOVqE6VPcDnkSUIfMu+EKvrXEHSDOnMi
mt3Fb0QA9bfJ2Wk+aF++I+iEK+SbnU9TF99/8R7i/0MrM00b4cs5CJWQlrlU
23QVJ9xkCq/oTQ/k9WaKLdRiMPTWVet8/nT7NrP1rwebrMBQ5+/1e3I5lyD1
7kBfa4SAvodrmqdqnHBCPjDuWNCSLV3OCTEUUTYwMUl9dXaxa97FzYZHvzCo
juCcNYoHD9LXMqU89+dVimVMymy+ajcyUbh0XlEZeYwMc4Ojse9DOo/87C8/
q9UVAjsPHtP09pSk2NUbvo1i0dJ26NJhqHY2kLzQUCnYMNR3EESMe7I3t0u1
dIiwqzpknee7OYeSE0LS8osteq1BQ0NToIbVFeWPjygxYvr4ocwUbapgi5if
ydRle0xq75HYOSR4yQAJo2kwIhp6VubncmtyD2lFZ463vjXXgwwsSqRjggP2
D6GtpUUr52Rju7J9/UCaF+kIJuqx6udImMNhEAbITKz7MbGdV2359CtCklHF
YJhhJ94N+vaAQh/4VuicPwVWHEh3W0OKWKvrfQkvSHBHsvmRyG4I2DOIFWsb
RWpVYQzTof0ZpZcmw+FqyGvsIV4zxy9PXq1Z4XKI5tlU1TQMiy77r4aBNA9J
TXr+Rs0UkZujtFgZJtL2wNqQdAHVlrZraXOgm+Qioo/HVkkrZiCgtJq9rn+B
W9hyRcKUl9fMCU9lXO1A6OwZWeLsvQjTwDREVjwB2y3VpStgYoCqvCIJfPh/
Zo0vADWdx1RGcHn/IRVsGe6Q8Fl2/YGO9OoLXaaLDYeXZNcrddZ8y6vRPTSR
U0yuVh/JsrMsJW/cYhi/03CrOdjah2qyUyJ/T8q2L2OwcgTd4ePRkMEoUIbQ
cIO3P7/G9edzZ+M/2pTHjfNigZeSoiPazel7UymTB9NbBvt3A+0E/otJ7V50
iJCKEofsLEhSTtsCfkDglieE0u/aCDtvjkp4ErztFefXoDPqLO560KrSTZg3
EHyYDqZSC1Z0M/pyMPzwr4jOzReu746OBDo8Pph0+n8RG9O1ODoAKRUPsC5B
qDVf/gbkHnvSIASxPrcnmhxYGBgy1FImccDmRFlSIL9+/IfRQXgzpy3ZaA/7
9gtcUBg+sm60QnPTDuRTg8rebozX45yS6f7c+cJRj7J53jdxKpWz43UbGEXU
xg71kWuR4ZZ5FqHUnHzI9BSdghpknvcVwWV6H6CHlBJ7qFqljQUceCmC9RNb
vVw7AmZmmgzKdjPKftz6SW5UTQngWeNS31W6TVt7D7YfxzmjeXHa0vyKtv/s
OWyF+lXyR9yz6E3mDD6tNMwKyVnXcIwX2EqBH3fZS1HFsABvAPyrPc6f6klT
tiowKlVI/siXPUuq7iF18UviZKO1X5X/eVqpYDVSwOXeHlDAm3eff093fCPS
DBkudKUALB6AKK/SBIjPWF9RWOBAWmV5VNQG4UA56MwKN/MyWoY4OVW4A37o
py5jKbOcFip5qfc25KLvLb4pdHcsjn/1As/pwKFiRlqjhYF1hWbrXjY4D3hw
yVhNkYu0WSl2/oBCb2Zq/EPVEUJypWHdqROS2zi1cFOCJRggG9ABW383/TKz
iZTpUjCjQz3YzmXiLYzjTYXKRBsHSloAbGmg+B3wwSOgQNewE/7JSenaujWo
MOlwEbYqaZqrIbX4gKnQFjC13od8F9CaE0A0G1mCIMPpZeubrPdKzJonPJZs
fIIoW+DVCNnwJ4olPT1jJWEqa/0AwuH4vJIP4p3dxhPoa43R2o6p1/2I3Ep9
UVYmJyFCJU5VD/vRjOLl+fj4C63PPNm3rtZ9RghpuYM/mLHmfty9/WLRya1c
oc2aRRu44w2kd8oK9b6FIDHeZwL9xWwDbz0dX9E67x5oDgc1sqgL4dm3guu7
EQ9jcrTcZvcQgSg6KnRB7hewgvuB6+CUNYjJ00GbR6mBRTK79o+l6Zu/nW3N
y2McUotw9rYv9tqc2JoxFUPWCGOceagrN8On4DwbDTmRFkzOEfMsTGbiqVv9
GIqIp3pU1N0aYTo1d9YbNHYMrI8ELoErPZqpj4nypsc170ewRYrkXw0fkeBc
cQ6bCJNlzi+6qoG4i0W976pq7EJ0IX3CysiMfDhZ7fi/jlCYRZVtS76styx1
gjZNWIp5GxI/2pjeborqNbxoPFNfcALxM53Ezom90mLXpe3aMnUgep07OlNM
OyNmogq6QZ37HVkMkCMnUy/7URBka3s/Bz40dPGtT+YGU8wH9rg25Pv6YmKs
Z+pj6a0QT0o9gEZuDLsWoUAeBGrvUCG1EbToTOyZCcBE8gYM4LrsHiDDokNv
NsPP5nqseo40M4Cc1QU7Elx9cYPCzgc8SdZDJsvKxHcfvLikywJ9w6YaXzUs
Sh40pPvwsPNL5viL0lGxveTdmYbUp30h/R1Pp+7AqL9nf5xnkhbh5uFgGGWa
KKBOzi7DBuzz4brccD2StCssu6huHVhIYRPM27++Swj5wsgMOh9X/Xs+b0pm
2/vJEifsPU8TKfuiCZUi5s23++WYEcll1jOnN+Lg+BgjvKfaJg583u/HprSp
wvWxWhMZ4m1acFSUU7PmOPZBImKOdIuRnx/W4bW62JY9QQMhimsy9lbqpkTS
2MzulzNW9PBiOsLIv9HbeVeyO+qOFcjpvjxeXrqkt8RLidlmRTGS4Ftfk3DB
8RXTrv9yW+jFekPwKT8ZpTTbSlrvbXm2tgUx0UAasmFFjO/7jVx7AyjGizp8
MdJCS89tupYurySpd+mWmta9NJ9yPFHzX5FZizxV9OHcRPKYU7JGwGFbpqec
VLTme/2wAtAHHCzgb8cXfcX/eW0k6cJW+bmmepI65htk9sfRF+YhkH9HY6j3
HpFdDXRTqegXxbmyH3iza6Y2bMm+CqLj0V7mOR0QLz2/0x+JbtEWVliFhqij
TbiG9juQhrsmuci/DQFUgmISe/89iKi2iY9XNDlZ5e8o7qt0pw2pF/XxUMTf
4UJlFSYJ7YKh8qTc6373U8fNaKPqsXEe9HkI5XwGfwSZ1nPYI2RvuGyl1dKw
b96zWJpzCoZLFBbtrsFTNhWYpXhPXxk0WFVq8SDcrgIPjFHkFlJd0TSo/ndP
TXkqjAXHdczqfgSBflw7ZA7/lGyGQn6OOpT2nUuOLgflx4jeqXTLnT3fO9BH
1eRsPPTyNdrIxT8ZZD/jemZNUcltVYPbezWWcsXB7G2BI35WJDiR7iI8PIau
cbzbXd4+P2lXa8qMXCaZCxkJ8UQa5Ks7AdV4cc3Fib4cemZnc6YYeUw9a0L0
E1h8WojjFC0e52b/QBh0C9TDFpTdWP1mWXeRwn6Cz7FeMAZC5ameycKSKvOb
RQ/1rFHFW++wWhxuuNd6gf3qGYny10FRnp/HP5BRzTd0RgsFqtABEKUljJCo
kGCd0L46cpsoqBRUIOTauXQ39jvMO1UHQw80rPbwPbOBK+srwUhq7Vhz1sZR
v2Qk7klOtIJDJOA0E4U3za/RP2MT7xWh835D+AWoDP7rT778F0S+j6pNkjsM
4MRk9wmWz5Q3AbAAebYPpR75ERIm/bBgjwD3xDx2f7G6v+4tJmxHkEDzql0Y
7k83GzGz57g3ebd9l+c4PCT+WfACvMF2DfADHC4xl9Qg8DQFAQAKYB0L5nuU
Yq9q3Csjzw5eLrhl0bI544ya1KeB+nGWay/84IoKQ91+zMnAq54m8Wv0maiR
DXvb3nigJB6X0M5153GTR2PNQP+WH6JpX4IEJdHg013Z8Iy9dAd/w+kqgRaK
O8Ct6ZsySxbBRqCRC7N8Ye/SfP2GMY4UyKs7ncynsKKXU2wmtK2tsiB13QzI
S2ZfMj+WidPev/oNJV6+SYMDzNySPwn2ArZf2kAHxEnU1TUGvzRhSMAW3YDC
9u9l0c0IAzepY1TgHylVfN+w8Ig4mdB6bpxPex+8f0iGpKg5e0JgsG1Nm8JB
zIyqrFD60dbNHvE7kAnDEsdfVjZk8AS2uTxWLbpDXYGOitZPuR8xpkxat78q
rHArRzoGw6KErADRbxuKpTUlmkMYbd1Z3XIHP+t7gMRf+sHgVJwdnR6ADskd
yIqTLRb02t4mbo4lGlfRsyJ7fxQkmRDS2xaSsNKyx85wg91adlcNZnGceh0p
ITkmvQUJxppURzazTsd4QXh0Z3A+RdiIf1XHm6s8zTguxOWwJhlHYGThyNfR
EmUAwW/e0Hv4LPNIRsV0vHtJGzZTBNua0ik5r2tMejnJqDd6B13IV3xb/mz9
J8DYOoLW5WQHlxFzoTAzT5/depBmyCDqHa0G+SmJCk3aufbrnVfCKbT4iLMD
NxQBAUgDHmkR22+DWQIBPhZrY09nS3H6WROD7iUs2+2hUYfxZqroes2iqUdu
WPkqVoXmvsTrSujakl7yXxFMc6S0oHQM7TGxwrPXMiPSZzIcViFU1PGwHrNc
gz30yz30Il8wwhYUYByw/w/ssPfR/1PZKDAqYI2gKklYTeJJy126aYN38pH/
/1QBoc+pv+KfQobay8nBKZaTaJh3R5NUtcx4KKJG9ZSN72cps32f/bjPEaPQ
Zmkht7Un0srutcY4AfBwSfSM9cm7m9De2yWXbsFVPplRdeqtMf45EHjYAZNo
xhxAMdtnjgt4DZGyiBfPlYR0zIwPl0rZWITXBkpW3pUehS3iMv3qrJflcDB2
CNre8Fv+613DkpDFQcs+QDioWubnge+04o1Sbt24CeSP4E92tEs3pVrVC3Vh
1hqsUvNjnq5aeAmksACIZvXLLcAHFHZfMVCmTeLxwICqUwYZfVIeh/JPkRNP
UI/hynzf/4oaYDqBZEl4fqTytWk28cq+LFpLk9TYmXLSHZW47UfJNeuyN8g3
dt5nPXNF3mMKWzbVLnwVrl8KvZVzkZfV5zz3zDMlv0fFoHSuPgYbx70ql89+
GnMJzEh/4zRbYA/RuPB88beiFMB17lTzMw1S3CRXNxppBgCjZXLfruldO9R2
bquQ47Can4G7YKdheGtmJbe4YdKJ3m15Z2jPSGlNE9upnn8RsnIOAB/rtjyp
4UW+VVehg82Xuwv0tHw7ZsHjZEe5kFjz0GQA0Ot5ctXfh5u7cBbg/cZgX3Us
6PpplFdYZchsQKMIYT3Ntu670ABe8oAKpa6Yhx+40qCTsOc3Irm5asqJ3a8P
igJRhIMRAQni36jEpzTieqarl66et4cFViHIxgcUAJjwCC+eAynp5/OXgSYu
rA08SmMpJdrbmsb0uAWs795sSGDfh+MhliU66IErigCtPwFP+0ds/7gXkZhG
bVm6eZOhV+BkFqCc0Ag0AyQGIJPK6kiGTut7jJx9Eckuwn/tWPRomfBx5Sju
h/RE7GjFn8cpEMKeEOvsir1n4ZS9AGBtHxSfQ5PCxnABtkMla+9gop5nYrXU
noalHenfUIlokJyc70I4fUgczk2E0e9K36Aak9s27FpnxTwiqsBHmWc0WESV
4t96iP2PCbAjufpYq+wViIhRsiCjBehkUaF3eejUyMJCrL7dljPEAw6eTswM
1YVS0jx5FO5vlvkUIIx6N+GFfxmUYIFyP4icWjx40PN3JB/6Jc0LuoMvvZKb
d5CqoJuHr0aDWJWT+1FkEbuu7LVxuaS68YyBLTSM1DEz1lGKZExE+VgFJGTS
3SZwQayo1WRYYjN3rLGVq9ug13Ul4ESxPn4Oy5JoXKDW3yVsMe7uwYFQycWt
FvPZrrdi75rCOk9vMe0EwAX4Y0Ba69xRRlMiJIieunRRa/1iuC7/ajNh5vKK
25zqgZlDojfbmeyoEa3rGq8N6fPMTtMW9TdNqY/Ogh5cQvI+XOKO3xUbyjkC
UZZ87q11EXn3J394YrDzHVEBfJ95yQZvBioIc1lwX6oNlIrcrich2kxJwY3X
+QIAJRUTPRyLMeye44weTczuiKoYqhQ/lKSf0ScElo/w6QlgYheSt3bAyPmj
fF//Kj4XY/vRNWAhevqKph1LotQFWKG2u4O3ImUYSKDddIO4IzMuKuVD4a1I
NL9iZWuYCQAPyFXhXFRjxnGDEPljM16UNXdoI8NaQgV8QmxntbIeCTIDcR7n
EBuw8CeiSaKd62dNRzimgbJmbYhA8NnPJVyhmNcJmKTUeboXSt3EKPRYt8pp
3CkB0VjdacnnIEpZPlReig6pMgfe2iFD0ldi4/Z0HgCr4h846swSVFdhSZGn
BJ3Hdlr45TczKHFnZhMaD0pZF27eokHpF+ON/BmdfLgHWl/GthFA1SopO/ny
31p6O5O6lt8ykDBjQYJ4jxA+dDKtiJ40LUxf9GIlO8F6UrtB0Zar2WwCvt8v
8XW9hf/JMnUkLwquUHpNz0PLlOog4IzU9oM4hpamhpPHU1AHcUhP/w3J5AnK
wax1MC64lXjL3GECysJyDRupWBtLqs3NWx5t4rEJqJCyFXEIyiJo8pN0tBL/
B7gpCx1JzI9u5tUtoFboDLZcf9ZW6ivpv3MUN4ZcKatgfByLKQSFMHrmN9en
75lEMkJEJdflRYMyH87Tj/834MjMkK1xg/tnYaNw5gsFbdvAzASn+If8Mtti
CO88lQiCzmFgeb8IZSe4eBLftwH/SnAP8jIlXD1DBdmXLXVflXmBuzMUdVYk
0gZHDYjhPdG5Q2GYRnK6mvyeUV/OaWUve+Qt+I6t+2pViYfDKNbq2Typ5eWT
8350wM1LGg472qphKmX3GLfz/hVwiZ2ry050CgfmNkGpctVlbPpqhC03o8Y8
mAmyud4KbblBPfQzQm7UYKGnduV3CmZ17aZPCITAC/qlZmDtTXdc7yTUNSA3
aToIvlNe5f7Nn3z5NXc/zsk+ziq8B9TApZYeFd3gs15r1htNusALaUf7KHkf
wFDe8jQ4ir5Hs2g7ibCGAbjVP1J5wCd/DwjpLPKtttye4vjj1MLHV494oLmB
NcDUClHl3YxYiSGkJI3ynMVJ/yeaguaJlRltHtjZ3TtPIHhNDGEmMSgyzFVK
0+Z4chUlZIkvMe8c710Po2nCF3pLu761pyH/efg82HZtEbgzwQn96boTC/Kv
r6V+OgMHVc1M4L3VjwmB+GTFKTLUXcinI67YRX4ytk8y9h/ZpUI/ULSEL89c
vl0EsfYk8pL3pYYpj/X1BCYpddyckgJBOULF0rO59tXpPsAURp3BuZBg/apV
kD8MQ9ho8/sEoGAIqGqluR0sGfMh+Cl8VzclM7Emhx4A80gqHniCy6lzCNuB
82yfKDdbzYe36aRyypJA6NrkH2qHu0nrryqRvkHUeMmavio4cQDDs1untLuP
Pi12VDW8sCI3ALLvTy2rpqSC+PNbN60ibeV0DC50+MRCMJCsQDjLkFC5LsZP
Hwv8wMjM55k8ukOiJyFePe/OOP/7kfVJ6pFkhrde8lWvon3AR51dBCOOx5uK
bRSSZ8db+IoUfynE4NiSK3EGZg+cogHeRbuxyyk/FA61h1eI9jL5KQnOOOoC
i/XvWQzzsit3jE0UiBisN3RqCkAv96mUMJ2+eTWKw20gdeX0ZRdhFC6oAy7t
NoqJRFl5qbKg+SR8T0I+ROc9mc76SrKm3y82jAjnYsR1HMqSeE+79/QTnZmg
kAzMlL5TrUqPRbk24YHV1WRstihuaaAmB8z+cW64BBtepMQp5ty+nm12iJKS
kw8/4DzSZOfasbwbfOZ4fIi+tJYLJM1Hb7DeAkNyTxhmejmR6YO1qShQLYGu
UzNIbwZBhK9N2p6E7dqlL95cH1QM8Lx4UzkUNBRMP8+UinpZ3HGoZuixNEMW
fnkAl4bDVyksbTPg4JfdnYrm4LQBJHPOCRHy1s8g8JI0EvrtiHoFvPUnq8Ve
xtBhsVLpCIGI5jvyaoFxJaJXdRlnoG7nhSEZoO936eQzKYmYng1PH/t6MEN0
Uk/SLZ1ouDH0Ock+z5CLEUCEQhlnIuEtPCEr4zD205ROT08ldHAzfVmwecqk
7xa1KEOvSzWRv6PgedUumXt5DMLH51Q8nZw0laXLz5ssbXuXlANIwIVTAVCr
rFmjNRIxEY42LTbBt4vxwbsSiCXBLsKQcNr2uxD5pMHRVtr/0J4oroGkBTDq
ly6VzQAwCfPnxyEhzhnJzYsf7a5QFCSNz2zo8Qma09zESkQK7M6Vd9hxyzwz
DmonAUYVuNeyBacjJG3msExpcYCpyKsGRuEvjh/e8Uap/Ra8mu11p/RSzKpH
pqSsgyYlAVQkCYmZiNLCBKzDFNkgkSocxIsNEEx+8Ox6sqlDR1QFZ2K6G68Z
LyscYcq6pOVrDhBICDwaVrQRFTBhTLypuuAD+mAL6qw9TUYdjrlY+g3afytw
i+mYKPLikSjnu0LX6BxNIff1Eb+2h+JgO1DdDbnJQJT0wlIqs3SHBEFLu2Zd
wJNmreOR/Yl5NoIJLMjCRQDIWuUzDjmcj8qdBL+8xMvncoPUFnT7XDcwodce
zYZt4Y1FTTld2AI1+MICrpQ0QWUZE0ClDZgxr6sdIlIqTHhirpDKpNawtB2M
E4rq4VfKqJNXoyxwYI1X5ZBWcLM3HdTh5hEkfA48t4TalhudWCLHxSEncOdn
fl5P1ucI4kEblyy5MTDQs9t9tPZERAh93lMaz1EZu5+UNiVkaouxh7WH2978
8eG1lgh2MsmsVx6ErJ5I/otB93Rg3MRc5ZbRBS8dhhwJjdiL+H2nppCx0VOD
Y507CijxVvAB/5iP6ya2U2sBcvzFGiZZgwfBy5zjosGRbj0ed8yFiXcfaunx
HGw8ZiWgaqWFAjH8+GwMTPbVV7FRFfxCcnGRq4aTnqoTshpTk3Pk08sV0rxs
gtj34kJ19n21wJoyhFV7DOI7a3yA8bK6l81yRBJxD9GClgBd3eHwmaabQ93s
T59y0oKutLJwCvYQVf92f6nuFfBTom60SWnSXBP1pf2VXmgVlgMM4jX5Jkym
ieapwxuNgXjgjI82PVTudPpExfBiKtcvUB29dhOuDW4pk+pMcQ+sKEZu2ahr
zhPSX/FBl8tF/wVhhvezMQhx9lG4mj3Ceh2vecx7NR70w9DE2cWLJnw/hz0Z
oExfgYMmlWb3fvVASkec0JuN9C/wxuv2LVdG9Dk4+oIIBDMWnpnoQpHQOgZj
5WmDkMEzZ+j1hQ7Q2QmzTc8jqWHkokFeK/3xf56L9SeQjBhISKyzimM7o6ti
aE2Ux7MrjBWnv0PLb/RAJqWzs+lmNgLVRuhEjjhNyWZpu9HHxC30OKZTKFtq
cIupbzkxaqrQyorSzq5gTxC14YsW1fzd/RPhWBjyTlKM0rgSVTADlzHGNgvS
Gf6OOcKntUgcZvP+xyoIgmGxRg+Sh19eD4vGzrDo/o9jz+k7H7v91Wdz74Yx
OU4lGSiGZMO813lqq0Dyve6i3Z3B9eyc6zcB0Y5pC9+fYKlmP5NlJTwn2by9
zMG/L6jUEr/nT0xrZqekGvmUfRMOlSgAXv5EKS9cdbE08WYaA/Nnc1/UvpSG
eRXEIjF7fCRL8gtWAyR9MLeCkAd4XyruhR3kFClYcaxWVeHbE6cmzaVILIj1
5JE1I8ZqQfXy/rDBwPW2NAjpCWXp4OjnZFyXxHVbyuWV7y3KawEc5Ovro0Z2
yUgRhmpHWYGfr8HLCJJ29FbfwP3+a/On+0DGAU+EdPgVmadY0q6Sz+hMqVWH
9pwCGxnIytiY28l5A+qugasGhdqMMBYxtZDmc8vWmKt8500lAXlmsNGjFgew
PdEBu54BsmyuUCpetFcKSqfATxNPFjK6q9k9Y9td9s75Q7g8YZmUSLqhNAXC
PaRAUjLm9hEnctjVpM1flutlIf4SWf15Ia1GIcoW5qVrhM2xsdZC0B8ZoTxl
AgEh7FaSwYnMZcnuBGupJzH07h/pud+RVggPJuuPa0ign9LOwym8l9Xhd/1W
wZDJPQsJ35OHHOfrUknSyeDSwRudXEBGUxC8/EhAjlLlGDvISiA6aDre4YY8
5jbk5gYEmTlkoWyB3yeguKOiiS/uRty6HVIfMSgOs+xuAcw89lRodE3HANQy
nsAa63aIww3bsNkHLYjM2SjSocxkyvJqrk4km7ZU6LgR+w3j9HLsSIkEpJHP
0yUvtNVeWhAK4qQyDWuuwRBwztgDHxVd6ColCzTNkTDoR64xTjeRXX4y2YRk
8zruQljA0WfzQU559lKnHxRBlKufemG9hMM56aawsIO3JdfOf7JvcP8DUjsQ
rxqtCRAqZQ0unbyfvhT3HNByUPbIRBWTfdTqjbmtC7G2BhZY6CinXWYWuoRd
aMJ6PgQk9ka4qgOzIGw1nylPoQjTXQLT8CQkI0a0qqF9/7d4oBmOY1oroeGq
ahFemkoGRDKrgRTjx3E+JUo3dLejcDNFLkIaBd7aUwi5dKAj1NiPnIuFbUWM
PrakNm23yr9qxia9/4tVZfm55j7Rk2DMfUIrlSCxwDm+csfHtNUoyd+f58IH
orSBqFHBg7sPKShFYMvfZSmB0ow9hF2yu1pKGjtUyqDFL0krjrqQNijjtCrU
rRzH93iYi74gMJARLWNr+YXh7tSk+qB2XpEGnPBKdJE5C87jQ85MlaW8i7rw
A1LDe5UbsRPy+v07zuSHhD2FPJOjUReBEjc0EMk6n0zzMe2fAORKxhQkHQNR
iCGhxyqhVaqJC6s5oNMVXamSbzj+VczQI7kPK8hC46vp1U6auDjSIKXjDoFx
TgbVomfbbjMIBNPPNRZT6qXtzDV8wEk9C85GfbzSvmzQz7TxkKJcDUSUKBr0
GO1Xw5tUyO7C73inlqFUi/RhFCyfHGx8VFKzHs7fWUPaIky8AnvFRzUaf6Ut
nR++6bpcE9ZAHHSHwMvwnnQgNOgK16zih202CBuxFAsFpDSxtMiBj9DiLcfC
0cyfwoj/wYa7oS98Y16Q4VwIjDjOz3YdrPwVtyaEV1wiHX0asXMxouBd7zu5
XJwir5TwA5HJeFqK0rnDtDh31A4YiDY47v/49IzDiZPp4xq6wCwv3abnW+tq
CQQzHLw3I0Nd9yxMscxbc4hQHklws4jCwaYBO9uRFMKBpi3t3Q2D9r4MUKNw
lCrC7aAF1YEl5xZPt+9CX9+CpkpgjwCqi8GUBR/agAdRYrsKDvcYkOpr1x/b
bSHpU4bAU1q4khToBHKAzuD5P5HIRaEKshlEJ05VQVKdS4/lcTk6D5j0BVeY
e2ukoMZgTmmA5dzO34jTX92iuwSpqWRKSyllk8/WYZYZcT24E3w8TqvasS5A
b8CixqJukjOCM56hErjIgVyg1IkbGIJ19vh+m6sosFPP0TeVA/u1X994ZbYx
KZpe5UVv+5EJcnrqav1EGxJpRcY0TgKhKS/Fn/4ZrcDyMRbjaWmImyOd3jrl
PzvFJ86K1IXK5xskIWYrHW0JoJVXcxCCmjIsJZx8++WEyV7KREa0dTQsP0ft
8qvMnrCBzwBzp+sPpGG9Xjuh35oTBrfSk914vSpjNqvqCttf1HYKTG1WcpJo
EjcfciYJt5vzo3ImCkrLSBYgQ/8miEzZVWCskU3/20KAVxiJ0ILBbugaSLmn
L/ziwvYoUdNAiDgPX0Rw/9N4n+uTwvjWMRANuQNjVIBCm1WnOh7frvxRw/ro
OX60QgxkbWdKUmqZHecsu98vso63qpJImdxVASHj8Uy9b+KmVaaLEBVmKgzZ
GapBfJm0H1X8ghZyxAxp66UsrNWGDNP/xW0/A9VP6zsNJG3B1wZLdsLrrcWk
MHKFakdh9+lWMpjfPq8FNkLQjBDYSYlH5oDjD5u+6nyATypE6VWloFU5a69a
RRGVnQ1Oj7HtB2laZeXq/+7T/vJJFLr4UNcm83jr9yI02zatD5irmG+JV2jt
l+dNmZnrQ4FeTKSdv+GLo9yhSXvYGHu/JqADYPBWPh2mWVejP+uToS0cVhta
JtTsTb+EtR8gvyU2SG+hAQDagZlceLTBsoY+HPsask7SG5iuSI3eEA/++AbW
wK/EwYi4EO/159gFpIxGNN5QapjLx7kN1Z9u6NTIEgKWY+HLqKW1aOLyg1u6
j9HNMMjMtc6xgiHWMxCqPpeXgwZeIT/yBPSuhU0nWuQZXP4b5ISvJAzYFQ/w
BxkOV8zRHPKB9zFcKiIH/zRXQxjt4ewLlRBN66XtHH0l/rX8N/NZAopUXIZC
sujTs3SJvLQlYx6UHfU3W78Wl7LCndH+vnptQIi86DVTKan3iCF1tezvb8Cc
4USkzpVAY6sTg0IRS8i7KVvf+EJvV9e3q3me4SVgEBh+GeepDYZA76lPNZxL
2xoqvzA0rITG8R5605eOJU587j7qIz2n697FDUrj3H5rt6MuHgp/weWcLrGf
0KWHoSTgkyGUqkG9cP1Lyy8vDU3UGkJ181VIBbmAQB7a1c91co5ks6YtydfD
MI/x0Mx84aUhQIL83O02oEcDKV50Bn8r3GkGtepdd1srz3VXb6/fyDu72B4d
krvm5Dm8N8NPBwuOOuR4+3Quc5e2Wx16OfLOkFKaw53a6pHJ2dc5KfrUEed7
cDyXbizyxyV4Bvbx4jAX4NQEk5/Wor8NYqTrxOxZMibhQZogY3ROgi7icIrg
qTDwnorZ2cW2m3BQFdR973OdNvovgf59vk+su/u3k9aMunCXXOE5xO9judUR
etqpJK7ZytITE4a79ljoak8lmMSOwunJYY0M5qeEtgyvK3/SpkDrRk6dLOPp
yNHX4RzZkN/Cs9mAhfk2q35kqSm9sZ3a0KuIcVpB/gSPx+WT51mca5QcZfqX
4edbys8oaBslPbh+pXJXK7/V++q2ZmIWeFYlj/DQjywXH3R9kXCz6UzTxKKR
8Mo2fGCPvrocywLSAQhbJO2LVErpv4J6tyWFF0LX1bxDvL0tKS34HRYvG4Dx
nkGVqNyXboshgVQaGIOac9bQ/RqCNOaRXICPhF1aBrIeQ4PfFfgr94oA4g1s
MHGDjuyed4Sgzy1FZaTE5bNIIejdNpN/vAzmNbS/Wnb64xdH3ZL4r76P/nha
imxdHGoa733TaLJiF6YscOL+uHi9n1jh/cCPQvNgd9Vrkd7RkE4U6RbWzc8X
6t7taGK1/AJ7REkEP1na2FBEomlatwW8BveIIDzIlUdmntMxroPMh1extqGK
UQCX7zJVID4jNCtbmqNAYA1i5ZjU9Og/oF9WiuSSCeI9kT2JZPYRrFlpjre1
KzwLRuE25aEwXgYsjkx3ypRj5RJHxX8cj8xvr8zGw5p7WlOtyXVBB2yBiuyc
B5XjlH22Fc2/VNUcvJmQ00ZrUwtFrIDWwsjW/l26ehWUhqvSyPPuvhviFcDO
txmZ94+CUwycQcbVXD0UYFGv6tQHNjzKpKqbCDgw+o+cNjaGNvH+u0bl6q6S
KyQze80pxH7swMJvpbAzxJ6LunM33zzqG67ZyZsyMlNIxS2qnGNc6KnjKmzC
EtpCHC/HCFaI8EaBxZWrgbsxPMD5cmQUAYJgApvxSdQfkB2UvOlgX1Fv6cLS
ibxQmSOVfVePpKn3Rc4IjP9TRq9oM1WorIq0pOR+DzKwdy6RqV26fJLXchMr
B3A8Mw2PKWjYWZcrzjvKgL8QDuboSA9+NG8HAZR98P8ape/hEgG7CIpQOtgI
EIeWO1Wyzk5BQmPexvOvmCGPj9B/62ugoxQIpGHutFr+rBFtAqYmohs3nZLG
zWQD3S2JNrHO4+vAsadfI1BQuPDHVUYM1y3fUAVXgeN5aUvVhIi9L6eg5ZfH
+3QcKAEYthLeu51ycvXkUTOIyj7MX3rQGgzMxD1W/z/P8/qTQZL1uI7joFjC
E2Hk8LaEqjFSCLSlT6lk1c+6j3z8q66t1gfLq57fgCEZozYuYPYEvexWzexy
tuttJrzDEDTG4W6WFQyco8RPpMznJ8MbkFlNmV1oU7EBej5SYhQO+9whPah3
Wp2kUyWZxdCYprZFutPXoNx7RTwsSHSbQ8Wk+xEjRHoUTb7tv6vwapsrO3Q6
khQ//HF81OnDkZP/inNxaG/+CQbvgJHxwK5BDjyfwhFPc1fp66f1i4RAdzAK
kqqPvlrvJlJMieRRR7x2KcuoBtUR8T8WtYwufvrMYB0Jlm00ZJAODv8Qwwub
n4AM0INwbIKzt7y4qOpxdN7aMVUXm8vp9AzDk327v/K/ZGywrJuwgrWVMmiI
seUajlEHZAyovsFnzvSA2oFnLLK1HBLIzX+H+6NHoz8SsUPBbsJqHh0NHBVY
K8Z/96yEibEhM5tFTzZH1j9m/vudJsuLa+X+h+Ne5x92RosoRXWXLNKvk01k
YFw1xJE5zK7EqyDHpOHCj6Z4XdOsPZ4Bay+fOfaG0AP7ZPDxfcEL/Au4Gn9Y
HeRXHivwBEtZFvnesU9SmvzFnnH0GzriU+X8InOYacFP1KPtLK+2jVJG0Wyq
L2bZhsmxGldIyCTwF5/4LnUnrO05nExMIheKSpUQoxNzASbSvOUhWv4h55vN
JodDRixe4/+fY7tjuXBEsErmUz1HMO2NJMO8EXx65Bjf2EtgpfSQXRH1Bwb4
GYd9x7wPlzWMD+zW/N9vNu697UPI6ai7dUUBIAmLLD9oC1jTRsDSn2yIziIi
tisgocM+XNPv6qg6x1nKXbp6w+7d3GVzpmIN9toz6XM7zS9grXtl3MnjPne0
ipAiAJSEuQFgHwLmCCQNGvZDXkkzux85NovJx+aSR3utws1omqMzMa+mCAiG
paM2GnC+A3JB3mo4uZEYLSW9hIcFRHFD+w/J0CltpjWouo62Ycmp18Swh/eb
sMiFPA0U5upjmsjlNyO4gSytsO4g0y5mYyx92Vdwu5qEspahhbCbJYqXRoot
NGnHVOpvJDLlur7cdlczKGN2VdnCPsvXkO98vV1Y5WBwdkjLeemeYDc/ZxC2
5W/PgiO0b8ofnNvbar5ZJDICOQZ70u6YOs3H9wuWpGal3CBgBAPLMVm0I7eR
7QNx3kcPajTkz88p3Bll04y3ZpB7frkOg2mRXAeUF1Z5lZ8nbxI2/nQ8kuOU
qZq7mb44HZYK8PD1ZOlHvxqpBHzK9BsBEgrBfRTyuMUF2hVgRVEw81Ptk5hm
V0tkb7oaleJEy7jVgJVRxz8KHh+WeqzZjJai3NpckgsXHojBSx0xetLanq8f
njEtMAYurzWFC3cDoJO4FaqlOc092BOommTLSXq6ufTrMrasOMfazkysq6qQ
fjEGMiSzJhtzNmN9cvYYlqtLG6X10DgbUWRxGlCq8UPJF9K/1PhEb8MiRVLw
M2lk1JD6o4wUOg9wAeae5A0yyCwYMd5UdDUacokOjsFheHZb7f0yFGZzwC6C
AJYGi5Gyr1iec4WOnbvNc9FBL8mYPcom9fBj8sy9NEvVe3i9I2lqX3F0227P
qNXIJtZEaoYZ3CApgI357rj4zSaFOiT7wMMdWIKmXksDXSzB7Q1sP9EmG1ij
DkhX7U9lwLuDu2R550lWJB5HJbej+9fbn+eHOJPMzpNN6Dsc5zWXR2xMMQIl
T0XaTRhABzMMTSClJyw3QQG9SI1ZhTJMuXd3JorgxV/PN0tUIQ40UzvJgJrw
ngfL8Nz4kK3mxaKDMvEoaW1DSPfS7shChhYaTxOSmEEhJVyGp/e1Fvbxmlrh
95EyQeBcntK1weLI3YgJktI4DI81WoU/QyFQKDpCWaiWYSIqqGAz/4mrgkoa
avOwwCpEWW5qobwJwKy6YMsBv1aNki8XLmjwSDy70K7HMqMh03PBj44Hf7iU
5ra4U71LbF0LIWlbKpoQjoQ1wA5wtjU2YhysP9OKfqFZ5Cd4+JJczT90pMqY
1Ugrdij/2H9KdDcP6HLqD8Nw1FSVyjpEn6epYsImV+28L4WR3DyMm9KpPtLE
uOgXPv2QtHeg2zQEE0bKIoXcMaRx9kFnhmtDY33oBqtgMv5BEnYofYLwUTOj
2UfN5wndpLNHrSFdBPSjv2+aGs4remJKdfEez72IPx3F7ETfJVr9mPoycYH8
0gh1OMJ3nrvNEbH8p1NxGClnq+lKUfl64bi+DRSNgxXEHNfLOBWm4kl6RoKh
xbsyx5n2xCq8wfE79Tek9ewwRX0H4UsaTATJ07yLW5sYRq/6/tFjlC8s5q3p
eTIxC0I3Pz4g62DJH2LaAVVqa5ROhXgI8Sd4/jDlVEATuFJxu2lJuZ4G8B29
fpEZ+wEbMlMHhw+AciQ5qP74aHXiM8aKxZxP5sIJqdUk0FyI0mG4OCiJ4DtK
QadJZCvu5zgfA3S4IPl8EqNNCw7M2CZwAnTnDKQlXuPopdNt9Zy7+QHD7yIx
RNFWFb8SA/oRW45EVX5AsfBSEIq3o0u0c0bBAmQCN6ZySp4cAdx4qaJx0bJP
OszJ6rVME6Sbuqr6eJkUv/hjQgxmjW27fi/iiicQUzPiw+V/OOEaH/ITjshW
AvaFdbST9tAfFdvV/y3ZvXVOZRjQ3i6aFchzpXzzfwuNiT8GQhYUmlmNTt6V
9ITut/hMXB/NKYkZJCFzEZMY1vO8WSwiI+yyhshYQ3cpCRc8QMAMkiw6e0U8
Atr+RXJ8H/5qs2Qhh7AkrfUyDBlO86An1PdFu+3GrCzOZqwCkVq/Rumf/9cX
KBV+W0B21cyJXCIm9WlvlHY4A6CRQjl1gUnlJj/Wn8plRrvdcckgmbjx2swo
GEtlGyncB/9QaHmASwVKP2kb+/2oxDXDcctT6/MlB8o7mx+1Sup93UXuN9ae
Oq31nMoMH11Y4ja6FhVNNvaS6mLlKKMLx5C11zNBxcVzpQY5nQ5qmeb3NNrF
BnpMMunHgcOtDfm7brfaV6AWERHwkrEQI8RTGHbDLcedhEnqjvhR4OHwmvY2
p4Zz7hwiAZPRkr/0yQrvvJcNvIsLUV4Ro5i0noRttCOHptq37K2V3OFBbWPF
pc5CIUdiFD4H1/LbFkfsXGfElnxMAHY/QF9acJ45Y9KqrKJVoI0oHpylBigN
IWPkYPVqhRLOtL5gxfMsrcyYEX3Ti848nGOgtd5rZPndtDvflsKV3bcgSK5G
sYUVmWOK2wsci+DafQscoZ30EeNVnS8CpBLhdtTbfEUkZhy2LXByZ8GRiXFq
YiIy211F6y+t3JNQbX2FZwf7Zzjw6qxqXRZjZGy/TsywGIib07eUqDSwVdFU
WHP/NtdBJ379lXUXhi8P35wyXv9ngkKeowffhccd0PpoYMhMZp+VzF/XlKdE
BywbvoCiCv2Dm7pHPe4BI59b+P5WK0BuOoalxX/Hpvs1lztQH9gSr20h21qz
220APkYCWM/IcltLP6U6GDJzyh7YTWIURlgAyddub1KWP5NfGoUjewD/lfCj
SMaEWPPzuXCY/GFtcOzwMG5jZ1Mwy199xmbk4CVq/1dOTiim82gj3Ptxvo0r
tvKIzmPX9o5oVqrvluWfg3nWvOTCm/11BQi2OKDS/O9XN1VFNen3KfyxBAbd
59mlHv9PcpBQDfHyqQWT4cmyH6Y4Tu61ZRzkUFXK3BPGmRpch0gX620Cj4/G
coAYyXrSVLCvGwwOQfeKZjNxxIXciNcD3YUfRFKXoquLGc8A1JoOG8gS7C5q
vAq+khJtjVuIGEcx20/bigQ5tI6HImuuxxOaqtx1EfxbrKJt9tursdgXcJgp
9wcKugkmGU5chDrVg8mQobpsTJsY8AmSJ37XG9XyHzpyOZFImfyCP/orAS4U
E22gx5BP66Q1QLlH1vHLJLmHbQf0IyRtY4aJY1GUkCHyvUV6BBmF8Vdamqs3
jZ/8kNerETyBcESbZXGf/JCNeXNoeYnGCjPcgoUgz3GYNXRUM1Lzfg0F/Ckl
/UZR660Jugf//0n+vWIq9pvErSfwR0Pi5kM51MfRBvTKksVfWayBF1nD2a39
/dY5pEBfIpoack/6hKZcohGekDKK9qCZeTzLAcNYY5FkNMYVRHMiu4N4vrxc
HV1dpr4vJrh/H1pEnQmHMvI1nd4XmwiEsHGxd7of7rIwvjlwuNx8UyYqgvdW
iSY9EdN+AH+IUuIMS0EuQzRRBsaXZew8NEJDMtQhwdL0Et+I7Ytywz77guD7
DKyCtuAJEbLkLa4PAD4U8LEBktr1Yml+eTmfIG2SOhwFMxGB5CCF+BsySqAP
+dupsPF7YsQVHZT6ml85vGQYEl2hm6pG0dKIrgO37FfC+c3MmkthF5YBAFQ6
iiJFsGhpCoCSZQPICB54ULLlFnldLlSOUkCU6nYjCqUoiSsNrG2YqrKWu1bA
Rbt48Ioy3fLZ1XWb8dimt8Nq2TWKRw7bUymyaH7Qhe6lTNOwv4Re63QRoluD
f7ZtxzWAkXdIlp1fRZeN9Raugjt8W2BNDzFGYdU3/N6pCl/hunhasI7r9BkL
pY5D+9WwQOAWNXi/ybC6Q+X66IQ/MgUWchQCicLTEuPVuX+4Fb9UbqnxUadR
Jv2oBkG7sG+ytefeXAL3RHIc4UDAhxwOLyaF11nlXarV86mNt76Iz3+DoUBU
HVWEb4PhjzR5Zh9NQKZIPgNxbOvIr/ciOZRqYcVXU1xXo5d6FzEPpaJjWDsF
UB1pUJdr9VUuOxqeoa3U2E8sQBOE/hyVZ//aQty1jK/mKHYp+zhTmq8gBxJw
yDIgvk0Xxv+Xqztlj0BQRAS24pLWUP4oYfJG1vzBgMwfm/jgFab2laKHJFhK
RdGwpCedAh6eV4X5RI+AUkoSHQoFRmztTB6eKe89k5nXicUqB9rsWhNatt01
jLWJdDPlxglV2pqL2AkAIIc1StPTR/FIxpkIeM1y2mjNNCEH0vIt549tDm97
b0kD72ETAdjy+Enr32R/J7XBgGEBqGwV13g2/EMnxE3wCTCJThYtc7BJfsts
3KtDe6eFSiBGH/qifoCDK8IlBHZiaXfRhPt6kUY2p4ZNVWTN3wdA/XHjAKtV
ChUFCnrHeOOh9CSJzTXNAoHmYj+DPZqUdJw/JeWv01hOKX2cAIGEmv6sB0Fn
9Dqk/ukVZcGiaR+j+6JjUl2vNtG/PgZwqpt58TEcOFbGCSdFJiUHGTOXPkCu
P75xXuqCdrpJvkE2T/w72Twv4exiD262R+KGMWyJzZu1ZrBcfl+Ng2PQgIXy
Sze19ZU8zF9+efo9v0ij/2fh67qXOvoxumrdpJRSaP/Tlm4Lm3Vj9o0SSfRS
yWIBakO/+rCsYM9EY2U7zdmY62kwVxWUMSyHR8T+vdpMPNvKwpYIcFK60qpN
bHtLd9WnnwIk3MkyLCv1mBcQJ7U4QTrMj2mBd8+TPPVqYmZbi9oOJ349O+Ac
T4g35QIFWuEwpeY2ioHPC3QxGRTDbFnlD/mirg4fRYhYYB8fGI1RH/1g6xDm
kMg78nJA0FG3A8k4RAQb2M4/+/DD3rY3YFAB1v/PThTIvMjAK4cZZPYOwZPG
JcxVFMZakGFG7LS+wgh/okPnaqQAPzhmcDxLR8ilOHEGrEj+0JJvDQG2WN2A
qy2+Tcrb9effu3nWQXM4GMeu1ug+s40vxtaREF1rk/PcdVCxuzHcIKz2nCLv
eW8Hiea6UGiNYSXkwXV3yOV7RfkviBkTayNPIJmrFSmflmQYjrahEKrNfcMG
pyvPdI5SuoqIto8ARaTZgWmdaHC+slyGeS+yG69jhBhzc8ZboK4uh+FgvsN5
Vbupkd6ZwPnbQufRwA1yf7YDIYIwhnxKCtbDzro1BkUbjQYqZnV/15dItk6q
Sf6x6LOh/Own4wpCGjBp7dC0rLqKXBnkvk/xeYVGSz5u8agTDj9KRucQ4nGb
CLvwr3lnZfIsErxTnvYSu7iFwLPUXAOIgoutpP/Soci3BJRUH7v+k/UYaUp0
6lJaEY/yR9rdYOA8pyIa71Byyjxb5SdDRS/KueMcCI6bz6mPCij8vpD3bov1
J2s6iO5tS9/0Yyktbz0N6eBWVFQsuTaRQsu9bKiW23vEsCp2DF6xQAeWvAsS
/SGjefVdQzJiDPqlwiq/AlQiE8FpjBGxTFX7IWMa3DPwGYVwJBsQa9egHxp1
88ZQmDvxtIA1bI4JR1SHahrqUStFWfwFPaYZpCtxK40UyslBIsKLWZ6m8I1Z
r6uDK6YGMwVlI2r7JF+pVHaQ/r7JKpdV89dcYN50PG7eF7JdDIdm3tbgEsQK
/RbvMqctGaSQF1s1mY/kVZxoSRwZwgPZHkJnu0Y1qpLC6JbMxSXjhzTqmY8n
2EaDH4Yn37eNXKleSNk//tmS1aNEXeifZ2vqA7pfA6Vmx2NVcJDsPyMJhbT8
Es7OvTJoHbXrJGhhQIOP+81vHBmlGmfQozK67zQDHhwZ6Y+/CjIivJqW57C7
h/Ql5ddZByKgu6WSEqQBZmI4Ra6UvsG7tMMSEgjlvpheTg8pWcf0wR3I7N9U
P30xtwGIUW9srWTM55BvG4r3HwvFlNLvnsR7mWrJBn/pXVLHIYllE9ZMK6lx
O4eM93vfIbTEebjfqZRc+Jbk8CJ7ZxWiL8r9ljFBMetYSN1LxEHaV9xQQdHd
fk3HsjHKs3/jkC9mfqvtN29tTRFFGLjh3NTp2KTL11958f4BXCu8VZLVj+Ad
JXBtUGl1DQE1sZv3lbRJkcyfwpeNcXVufirb9cEoaMiIASFvKPHQe5bKmN/2
cj/pCrza/AMqrfwVTZs6E4OvdSmPruXJ9PCGf6z31Na7l81z4wA7OlZV/Upk
Qf7rCjOlEcH1MfW/fFi1WCzoqKnl9Y1gwS9u0q5C/aF7JMoTCTXk0UQrh6aR
78QAuujISVHqC/8tfn0Fo1g4hrJhk9/wfG2zyOB2ligeKR0tx6LnBNkka1Pu
c6CrMZJk2+M0eJFZeDV3TOqMG+aO6FHh/+gRKZw7Dcvvw1sHczjw5kUqfCNz
EA2wdTRPY+fFzBoGjFwCLF4dKhpJZxvkpCnUqgW3AUEr6XmQZ3xhIBTn7Bvj
GyQoLu6aWDvThw7ifgET4k0Wv3bEu/1bp7eKMruBVj+ppm+E1I/4j+bp0HJe
JvuuQJ5iOlXrdD5jIXPxH1oDUDwhbJsLYiin0spGaU9uXT5Xl/83CF/vHE5W
Pay+V70k4C8LugPMlmbhLC2uC/zu0NqSiVN1q7RMBuQeIjrsfqWuJLwdPzcC
D9fwBU4QUm/2ErkkZ687i/hz5DxFY5MiGG5o+Tu2cG47Vu9iiRBAsJHnCtz2
fNLl/O59adAkMMtWeyPjp07mw7rtnnPcUhHDqrmUmfX+w2xNDs2u2JaWdTE9
QBHmKbpZU+FRtxnjv3Tssxmc1AatKv+906ev18iU/E/ksElNNLnt3doeqfoQ
ASITw7rtv0d80vaOmIE2mlQOhCGBxf4WES4qpP+M0NLCwQkMhO8mPxQfVKED
a6/NaJDvKJsp6Im5KSP7F2GHQ5JZR9lZUTcgqbK00PP3vvhGQlvPSeHW+lpo
buTJlBuDvFHwBICSYIw0yXLNpSuDd5VZHy8UTo0dfJpeP8jhGHKTW8DbQnW6
KYUYvUF06RdCxarpF3KLWvBMkaxMdejOVgrNRmVH7I6kSpnKNaAreEWD7tGC
HTDKXlTFw5niuRXqU5EuYqzCLU1DAeyZoQphuYxe/g8dkp5uj/72IJN7Vgqk
zlk4XQLMsU38PnGxYuwMAFOkDB/KztcjCNBVgU2mIWTAVkQwuy2v8xhTMiEG
7HxpAg/yD6F5D2kt9F7s1wc7QjBiHnkrCSRFPdmXBDEX42msl+NIpBs3F4U/
oNw7IwhvOrMYgWtmLa2dJIvlc/MQCgrjCLHJQyzmg5Qm+1YfySEQjvrxSig6
ZRJWPPEoCKvbA8Ibq0/aaTPAr+8HxaEJUd3fhAeHx5+waMLK+WPryo+YpeWn
dDRxiyqz8SLkcR4BDyUaj8bFptbVTAIG40ZurrkHQ9V2Qkdkifs4Y9q1jmGO
pGvXAaIl/IXjOW1VqkUrgA305vJQThBmemAIOyUjFQhMjmvoK/KVuP/+xWaz
hjIbPNSD13Em3LR4Y04G+xUm195NRReDziVrPvjwmaPxw+mBdhFdETRk5tiJ
B8oJ/J92RoSiKxqXYkR6LrZ7aqg/KKVtAAVmGRB2ovEn6sbiKW+pHGPj4MZ4
pfX9ZEiFEWb9kfvhrobA1m4qTIKez1UsMHKJoqOtHU3iT/N8uPgCbxzC4f9j
gDr9NsvUEjueFQ0TnK+Wc8f1ouNGCdCVpuBchODI/PMnmoL/1YWXblearRqp
ziNTG/f7U+VgUDbGOB1XEEz0CVFDNyWreXTKifbHxPaEQdTTpFmbPN45/p+B
Ae3UVT3pvd97NdLQQR1lYYHLqqKytPAQniy9euwxNWNAEX17xaUHPkf0khmU
DnzPuz3OPycVK8Xh2tYCFTXopV798vybeDmX+tk2uVT5hoJt4xIfXY5tWifK
Nsn8m69huQqwmQU3Cey20TYYmVQzY1F0qlyPjH8puIsWe2BWF1W2YiacFhFW
4BepakxIEQJQdczAAWTSaui54D0JFUn3Ky1cIjykzx0kveA+4VevpYSBusaM
pJEZAbBJMxBmKswgJrqxfdGpcwp+IBJNm8meVmDTJO1lw0NTuZWGfQFUfntV
PriTfDks4w5CZhKEh3YbWHVcS447E6U/4LTDQRvUqyYKkeYPIvNTzs/S7u4/
JXegFbvNFzd8btyaXFm2zMyh/7lrFa2n6MYJB32UMJ33HbmES6qOXdZC+05W
itwJ2YGF7q5Pouu1r3dht2Y/W7E8+m5Dr0HKfUQ5pZHUulynw/sX/qw8jNbn
9QzJrgGJK6Mj3bvUQ35eGQXZ5B18Gw2HrY3v7tY0quYO+ceO768zDvAS1LaS
6XYQ5sxcdMW0gBG+krbB+HUmy59McDMauyG7zYcHm/RF7HO27MBE8qHOi5TN
GE0rZk1q7bfYSxVEZsbudFq2MFcqO8DC5UeuMBnAS9FYzqqDQNRaAyyJsJnn
ufwr3lvwHXd+NqLMlBn47Y3Pj6mxYM7cyvxy6Bvvvz+CQpzhIzB5ub+JDq/+
9khWMKzaY+CCoAsB5+uMO6eJeNtVyryJfEYj9GGajQ0JuYYe+WS35R7erk6L
NqHVCi4D1DaT4KnkrARaSlNcZg3qe+umQHxBoTRBw70rmXNZPKP09y4jjYN/
aQcQGfSBUNYoamHqfq1tdLhsYD6aYiWkCm6UT6MPMBdwsO+ujJHX7JHwoOm3
u+visClk+ObhQs0c/tsvfuQL1K9V3V3Trd6D4yKYIV4HS5elUtk8ogLDFAwT
SrFKEg0WiWNvDeaTPl6u2cX8Jf1tJ7694v/ThGdxOx8b2B3wYXws9XJdxVwc
sQBr4vbu6J80SIsRhQzWyqlEuglDKgGdgJ3zP12aCh0aLtAKNyy6xOYYNMEp
REredkFWdbMZPoOYo5P31OBqD6DPKjtLlA2lJL0eoJcjr+A3JLZq0/0Prh1i
iZt2y3hDB4sR1HYNpurrFSX+LvmMwBduOl6UGDjihXcCVQ4/evMmjCg6srTt
rI9QDRGVDTDTBgHbhTfBBYc59Fbx9t2yv1smniwo3Y62T9sncmL0Njkh2M4v
SfLJb1eVe3btKVp6OFIDXTqgMr5N77pvN1dU8d8IWQYyvCzS6cJFYCTfJuyz
q3Lpfe+qKEaLrKaMl7vBkRMR5jLsonpNoxy4sJhK+Bf0GR0theK0r7Dqb02L
l/ool09B9FaRga+EfZEySkS2LzPqJgewXYLyST8ni0OBvWOkVmy6nqDfv4cW
sR16eFkdUSs2Fv8UJUCde5qljIwtypj7rwaeHtt6dNglit2Vfej0QwIQf0j3
jxpf33MfkrX9A9B2Cu8HCrrOLyh8jY+YxxVggV/CxI1VdfYwCLXZJJ8u4IXU
QkYDZsMoKgCXFNCpBUOXxgRX100taUjy8RiLRineuolE/EHie3O7BfSM7PB0
1xYeVgdhC76i4HdCiHyb6lOiY1MgvK8ziCVnzgJ8xvckcNcUM6PtWjqx5N3C
X/wuZil8QtQWGA9/kmI+15cQO3OG9Tmmi0xz5kBAx5oH7dPflrSPfvJaw0tX
0m68nqCO7X3Iuanje62GBnRys0wSlojk+4XrYOhnk+WlzxUBfHU9IX2/XdF4
BzI7CiJpkYU69LKLh+MX8D156vvVVUsibwa3eTNnmgkxLYfcThjGK/jsuNLU
XRS+YnfPA8v32LnwQrtRs/WNNbV9yXBC/r02czvLwcCx1wF4ObHtatd4QWs4
zRO8VcjNQODF6gKNZtIACn9pop1BlYMIm92zGpw0n/sFNxacVU+dxzqP/fzt
PAw1+Coo4U1i6oXq441KpA4MJAnRt4iBc2MTmMBEMxZ+Fyj5+Wl2Tvfw0153
H3Zt/nPi2VmmdUczuoJ8I68HDlRnSq8Ev7IYXpRSR1NVbZIw96yhQ1GOdQBr
2lX4YV/7vq+XenW3SRKGTlm/5Cqm2QATohcYJ/Etk3HmwFUqXQc7UPzWkLOy
5TdJhUgxwBbwKe3+KoOHlMNc9ctIz/dR0EzLc6JxCK+a2Y9XXY09zb0dD2oE
/WSOIOGn/o6lxRj2DwRc+sN9ksJ2aCpl/qC7WsxyFNK2NDGvK24DBZ7dZqqI
4raa47m0cpIdBemFdI4yqboTvzpi5R52LUVm/BC4QZIvi5QKIvQRpytBOf+d
qFYv8a2SjLLNYPEne5i4AHzoQU3TWrFU6JrRRBGyd9AbB55A+6Khz6W62UV6
2FJF7foCK6spG+oqdQGRv0AAsxWGFZjf0+z8BuWNn3hfXtu8ksfDffiOaUWI
tEsaSAKUayebb9Z9bmLqqJjyQ30VhuErSXAb+Ggw4TL53PdenTr5J9jVDep7
NJJV92UzC5IHugisWzjCeFhgGSk5kNKTI5PT18lfGXbTSrWvb+Wbtw2AO4p3
KCu5sdtTK0RFJya6TbqW7csN9W+OY1twXbKXXrzQzGRDctzYoEw6+iHfAUj0
bPO4l4qo7A45CRptJIZynPozxGYUE9Z+RqqqdQ+QuSYklgwEL8+rjgfJ8V8k
dBK/rpSb+7NlqnCnVSlAYJcvNs7NplIMAlN8qHYL3TQJHH+kksZcMHlhAfc5
HUdOk9BOhtzbbDXuWAItU2EHG8RzhUFRXxWXx8zcGd4foZ5sgyfF22uVxUOp
6e/n50B6gEEyZQj8ug+yPO5vH06tpnwdusmZVQbC4zT9sXpYU0vHSet55Vzx
KGMmvNif1+8QJ7bN/tfyHUB2GTaGpvLvpV1Y3I+rcyIWniFiJwbzsi4RwxMw
7FIPd13DdgAK3mAPbd05jjjFyyNEyknbMAUAXJ2RJqV9nthlIxIcCrMLAURG
/LBGS+40+dDkUmF+qXWbqj0ijMHEOGDTmglBlPZKtayI7pynU1PAdqKYQsgX
ZpPZlZqTeIRQ0bIMOxQc0VGBkn36zOnID4RY2XgPmiHj61aFBVf1IJXrL/ms
Cty7MoB/8FoTmCrSvwJaofhpTaak1ZMVC2fnnuebrfhy0ocubRO90JaJ/Mgf
jOvMhU2rgJpbOMeRDeuHDBMuJJ8w5m44+IeOE1jp3tTqv3m2dady+F5ha2uT
nYtvBaDLhfgrod/Cl0fQD0YCsf3TqZQL2HV0Fl6/ex19MGAIgZaomo6mB34p
ru3OgOsKquxs7CmuXPJzzo+kO8xI11by7qDc3AsOibPTzl+RM0zfmHVwW/gG
5QqBDNvvL+mVRAL0LFVMbhbaJCOHtOyWrG9mdr+s7dfI0DnsDjIuCOMmOLBv
oeWKkPXKgMUqlsTGSngpvZ0RnBhu78+A9imoc2rnkYrbpjTbneGjGb64MBuw
881cK1z4zM0Jpqo0XXV1uT4zYIxTCViJ2MBN7wD4weufuytWsCCv8EbPYfsE
oDz2e6snCUvyfbNgtP6i+o5dC4WQ8Vsu1Ogd+QJfNsSIA7hgelbtwhasEbOf
HcAgwzJnv0BQXnIAXEQU2rxeG477iPGCwxNoYnehSnO4dXWGsrOzQuOkeSdn
yyX4kl9ixxnVWj4yk2eNdxoxx2tByv52ffP/G6axXExLWNJxIZf/MoJJW73P
9vnp/0V1TFoESEy89Npw4dzR/cl/j7ssyyRazkmGB1k8XKlE0JN5UiOg2/85
v/40XZ8Xd/J9cX4r9iDSD7cePNidwyZnexemufdo+5M4O6t6RaXCvlORasPa
J8dKwo6/Vdfmfg4uTgctQllFhYfaAdFe4dOtqJ4qSgw1TTKQeyrtsUSdDGeJ
b4LYvrTFdZVjDkBZW2aELGDJX3hXB1f+P8E4kYELjN2f5YtkXXf+mp7zBqKT
Jz/ZooDI73+N0vwYjI8Y9HI+ctjc3XAleAerJQOImKcp8tbKltJoAzXeUr6j
5+ZFp/VIvtM4gL/z8XWzOV4Qpdujvzld4uhW8qhxh90K8qOK2YByZ1d/LfIN
o6tCQdZmTNNYSpMh+1NnWPyAoZyFqiaOsdrnoGX7jrgtfhCqgnDAYzGqD8Y8
xYTUKdW92zd8jVCVNmGNgcKHkBRx8mCu/WjFNPHLOam3gtADTX/CHkwPjkLN
AAHC9oo3tkErCWxPs/qSL4TPSwhT8S4kc5PC+Zh0sD7w8MPxeO4sAngLqTC6
PK4pLSIVthyitEevY7ut9OuFEpR2H8bDC5Vw+bPjyclkNtN1jADKLCUu+/Qw
CktWh1tbNz+kVeChlq5lGvx0RuK1hoQ/7OAlh/PrPvHay+DilZGJ4uNvSJL1
3K6zx5S8EP1eq8vtfgISqHlZ1ZIHh936+Lb2aMh4FNQ8n8Xiw94aOKJyI8oo
JvLAk1Rqwg03d9KlIUlfvhd86E3p0ewVTjlmna5L0aS7nM85NsrWJaHnL9V7
jSmZptgOGwZcH7e+nIF6Ho7q//cyjNTjOM+ILLCX2EI0P+mUUP//JvUclCMu
v/xZ3r5FlAdcCPH9Z0oWpit3gCmzdI57tONm+i9XFXoikJ4GBloM1mU0RrpO
XsfZ4tWGwgsUcVhxy96XEYLhTl43yjg5YIE6wABeyFPuELJJXpXgKIURdTMy
dWuYjJ7awRuuNrWlRoXCERNejvR0cW8vHBKaZRXkAvDQ+mI9jVp5c8p/KWMR
Z37l/KgYoy0nj46R3XHIcaYVvYNEHprmhQdrq+PL4QU2yAFtx8I65bk/Lb3V
7GKO699MBP2NHGbtVE3bleaDqCHcpLLdenmoHf1P4rsnmnBkPPnnEWiclKLd
3D0qN9PTzuk7oHjiOHZGjO8sYZ9JVqVqQNs4i/8ZLmcFDl553+oh5TS0tQ+W
dTafDh+YUOuplc78Qs9R3jSXlxTjTqDRSr5tLWU9MyQx0oh/fZb1IVPs8cz6
78qO7ayWZxydHBQSvXaSg30yaB/ezgjFEQy2qWUbgSEf1sBE5g33esGFMm3D
XSwae3Z5p2OKHES64AME40mnLzkkM2esvJ1+mY5Y6/iw8BtHPRO/8RIWEfBb
O3RUdEeT/z6WTsJOMcRq/Q4hyv6FzNIfG65QLh1Q/2+XqVYC4SXFEkmjzTAn
esHOceNpKmrsEY32KCwrIkQKFQ/nxaQdANIcmfjPFgO7/9MFls6/1Eewsjhi
dySOAccFYbRtYar4r/okbNiHjdDAN4yOqAzgWFQez86y1AR07iLdh1xu+m0U
UstEyyOAxcdXlH5qJVGyJtXvI9m9/RXxuu9eC2jbz/N4iukBFYq08JgBx5eN
Do0JVa51LE3W0iMI3ig/0FjDfXnL42neJxL2YDHhHEe1skbgpjZO5agQI4o3
SeEcujLGsCnFKXA+fjL6OVzMr+/mDqBZ+7iETpQKpZy/CmqfleqWoGnXuShG
Hxh3PwSomJM6agmLCWBMzEw+z7QDNg0sX69t1IDzkagD02bC/lMIAE7ye4Xc
MhCejmf1gSzkCVff0cge0hRAqiuUNI2i3HRDM2qzbVpCUjSxe0ydUvOTmRMh
mpYZTbIBl84Pcrhh2dgkGuZdqFbMbhHITYqxNfHXnHmpVCL2gZ7MMfQ/gQF/
+8QqGH0JNumrU+oK59u8dTzwzn2cNG5e7tqTXqGrSDNeNut6e5O5ugnD/HnU
9ROJKEShYsB4DtgecsJfG+0wNMMxkef0dGhlxprQSu+DCLWQY4YuHj8IhTwp
H/5OcqGOhBleB6HzgHcVzhjsmTQiZrZEO8vDF5NTzUWzLeQ/2RCRphM07ers
h9v8//kIm9alqJkUnyLFV1APGS/waya9gQGXB0RERu2+2ofxFq1zhFD/rhKz
MHFQrYmg4uAhr7/6n8ve7zkUIEjZ6O7jHhK5vVDPiTjOEEKSny7qgqQliAlY
RlGtcNB8KcGGA3qqX2F58bLUp0pLY+Ee14LRTVQjEdAid00mbbwZpvoeVpui
49kKOEnzbwn4BAEd5dHXpjO4f44k8MloAOsG43ilMZ/UBcVSGGSrrgZlXsyO
3ts9nrY5wHZPRAXdcKL/mKNJ4zbHL66CUfwspvtypi74y+HGHFODZPxpOHJt
VgrZMPNlz0ntwAQjiFSqZSnEIQIxlNZEZZNTfgHeKt1dVoE8L66JWZ+9bs4/
inm8AjSDvLaINcsxDIXs7EaheU/oI4fG6LmQfzIAIebmq+AzU0nJWri+VotG
wYCVOtXI1RCoqiBfOsQ+at63WIceercWqkH61vWAK4ky/Fz7Q9POcTrYXmnh
vXBmPr6c8PAV0P/1GKUM4TA45205wbOf5DGFydF3+rIcy/RdvI9imEF/8roi
Q1QxVWvQSpGJQOSXwYB+DTN/bfL5CQDCiEylSESu7dGJZSmNzsw49zuFug59
gJv4TQ9G2LYdMR7LwBlVuoAYmCjI7jre9XjTI2FwZgFpVIaPL8jSYGOZ3xu1
7Oxo1YW8KF1LLwcilsDAq7eUPcoTYSgOrTjZzi9LGRjB03gK9b69VDzgHH3d
OH8kztSxEQ3HvTumS3sis/gvDpBjICXwcWPhhQVkqQ0Hk11KoCc2x1P+wIJt
SEbVWO0vYFz5nrv+DqRRS2cIkHd/tXFecbs8xf9EJMFyekDJpeC1q46fV5te
Tbf1TYDPp6ZuYRMIkmyGqt02uMPCbWtAunGHDzpBu+Hr70eO6kMGAFozd/cd
PCdHu5rW3DRcPeHVSLTwoIfalaO1uM/Haqhj0gvgiC7iZ2JnqXJ6ldbHbkdm
hxku5v0G2VDufiJRAr0Vn5JWCceiH/5ms7GzHfmvdb3q+dCCkIrY+l6Gwbno
6uJy+iyAbh+sevW8RZ4whk2qeyQogjbNwSIiOPs0pnialAMoPifzwKHTbhbv
jXttaLwsHz1njtVpZe+zYnpGYALDq5HOprCHyq3qANT5Ne0vNChMihz0dInv
7Xq5YpXA6pV6MXO2LNdrnD+yVCH9umczbKEbNTfea1SYlkobMjRiwZd91nLa
Yt7D85TtgLrtzDBtzeYtB1wLmNPvf2rOS8PZOhTBEfwtPyIZbp+DZ40QQO/h
uP6h5duu9CdJjjH+VshWK2vc1MSFnsMEQrs+FO3o5bvIKTeB3ILupN6D3uWL
9Rm0nUFeiVLv+7wi7WE+9Wpx6gWgi1kcp2PG2+R3RrZmShbZYaWn7dd1luVo
H8EJitlYX48GonewB9dqbfeVbp8o4yJ4awGBAl1dkn0jTvgp9/QIQkU3kE5d
tZ2N9odSRQqh3EgK6Sa7MGbNH8fH3aRGwb0o9fcKJZos6YOj/LtwkdIn/IIR
RVT2xTsfD7O7Ghep0WpD0nyHvicNGsJJeWlojrdgDYvZ1F8Idi0lAAL/qI52
iaPTxxtS1HCvNZLP9EyMdKjyGORm0ytiOgJP+NYVIkNnwIeOI0HLpk2eoi1P
nfPRkpH4cR4dwa4UVU6NubJMbdt3DAVOZFns48UwhE0AsVrHI9/TKlTdvWli
o/Jql4CXb1Psiz87gifUV0vb5Q9sMkwtbwJ+LtkjZSUAdodE12Wn8+325aWI
ITgmoEkr+WtSUt5zbo0cC1QR+kgiYTOU/bF4xzrA4JXrHxU1D9sIgplMobcE
THKmkGT781MNc98TiKiUE+y7LNLy48cQu/28851p2FHfM6tCN2wFyroPH/ZG
L2nLC4Yn/6WHrhIC9fbQBQgfUXC+glWp2tGcpVNsitWI+AUuC/sbjJK8Bnh1
wOlR7/VmN00cLIHr3ziVr62VtXGmu3ziDqmQNpnYibJw1RvXwZ0OCUmbtcgw
R7QenreUF8xDQvAJkwyyc6imVDK2g2tRn6Wm0amQtffirI1Q2FqQ+7dLM9hD
LfhCgPh9f2d8L/1Q9i4vxOgCPbptdL/rTd9U5XF03L7Aa+gCnIuazCi8+44W
vG3sLLzZhJAVvOxwGOFh6KSySFMI48oY34khovJzmbqjVNJVLqF8pi3pSoiu
Vqefc9dy+KeS7gh3fATf8v2aXFcE90D861EdwNEYQ6u+Mc1sU0YYsZn7T61L
1tsL+O1Lx8683TDciq0uSz12eMDYHMZRydrzJJSYjeG2ym/JgaZYwF+mPg5Z
kiNv06WdyVrOL5skdkcG4F5+/qV4ukX3lWu2+zwIOVbKdLnzQZBOBCRLjx8g
S9V/eScFIxV56Rgw2Hvda48Shpu+vzWOG4cG7QyC3BjuTVrL+bco3ujBfNAS
jgGNSBgdZT3gKCITcnRrke8ZEXqCKE3MJQq+37k3kyeVse2akAGDDOXzdFDr
U9Ft9AaLBqitwAOgosFiOw+35xNxrt44QuMtpZjGH/y0GS1co1pdjYr6s8Bj
MH17xKrlejxvPnco+8pXGhzCxjL9XlQz1atGxu2RTrQKED6dQEu0zI3kVbde
J9UKpajb4rCKIXN3g8DKtgJiGySdUIW+0vMjtEfT0EFkqftiHP/4cSD30oBF
LaTcppBDtQm/9YiSDqpPiiZ2IXd0EW+hfqvI4kqWLWMjqBpq6wxLUdAHASSf
qsfbuST43UXPIK5CEKcqQNIL4WKsv/c/hfHCqzG+SWVXLJdyQROzKpdcoMPl
Il8otnPWDxm7mRnYmFN8hx3g/A/GVDy+Y6GDWuhPYLm76ieHKUG76FYW4fhr
zIq7iu6CyAOLWFIc8Kw2AjF2rMbH7nkI57SLh1r46IlTwX6F3DL25BIL2XA9
WGEdVGJhzUZp3yxiFgQHnM/wz7kvmwg036i+SdQjsxa/NSRfa6kBpe5dVUuJ
YtWP0WCgSQ0UMRyHotwtGMSv+w3EXHvolvJPAuhCj/J4Ao0CFyRj+SgPf5t8
wTCkmQtFAS/0FBjZbEqVh3DACS9kDAyl8rWewroZSFVyK6LNRMCv1rqW0bBj
wmep8pBiwXVZIVOgWi+6rqo+B0oeMk4yJbs1Vv5o60VlgCWlrtVMCTTLcocv
AHMp0QvYRNAY7TNa1PG7i4dZEfldUn5nONDaRUhCaXXYjzB0qNl3MtK8AqN2
eUxAdUiYInGfG6frhlybXbUijGNEYgH82ePVCRIPV0NKWHCj4XCLzq/IGNqA
SAGH8MDPqtBWJ1twaWPxsxAPu1NPK/r6FBVmoiFynRO/3+Qmla6XJWM7ztQZ
C75Yy9+H4QR0j3UVEwzYMambZPBbyBm7/j48/sVx7IqywCnt1i4KFwuxSPC8
eka9IGyX/JN0C7K1DEZy2miAT4JudBZdko5c27Vl3WulfHuNm66KV/4vmayW
M8aQeiwYiG04LQbFfLufHteqraKgVbqZEnbUGsz8LdRKniH4Qlr29W9qWlKU
5DQUP9RyMZpKrvg3B66aCeIWXiuoI9vIt+NUmbVerjiSfzNxhZ3EyOsOw6aA
TCvIgAb0iPXH5Nk42JMurJKiBvACGTTOCaPrWV3Kc7MdbLo86fMsYIzXdHyI
KSOaHp1xDXNWJnOFvE51gK3ceJ40+2qjDz4JLeVGId5p9/EqqI9Y6xHdtsNE
1hjH9NtJwb+jLQL+/sps70/VXYwe4KgfcYbl7o1OHbEKZq6Z5HMu4typbWKs
GTdyJA2dMX1ah9vqwzQfUnELiSxL34NdptrawTg6UBX0fNeIIoIhAbBp2R+M
T9LXaSovWueaM2c15PO0kK9Ja643cVWBLxrit3m8UEKRwJlm1gMMsvJuiZGA
BkDSfrd4Swc7tXxZ/GG6Io30Dv9/Oxtsb++DL9AzwnL6cHQzJs7Gm2drejNZ
pTmKxI6BkNTIPayw3csbfwQJ5QO15h2W3zMzc8oc9ftOPFiK6ZaBGt9WvEbR
hW0doyd/rdV7nt104Tn5PqZI7S/4sViVUv0nQwbeNyGnOVkqGXTRk9esZB27
cr+JY+eDf4cN/2JhHPUDwceufYq5y4G5BACeL7xLhH/T5xCUp5N4MIziXwDG
lgFv1+rbHwUx97uelkpJVQweGAvGrfsz7xZsmcxAqbinkC8BZrRnybYLKzdH
GB1ZGqw0a11cNDgLiZwdxeapcYuhSLy7qwYCfE6wVQ1RfyPyKlWLHVV3/FsE
kmB7pTy/xG5RLhiy9t1Uf9U9RPig2GHZX0mhR07HbYfcdiOCI+EMcjSJOyWB
41DPC9kmZ8SGDGp8xjCPnD2AVqTj6qpr80cx8vGjbQbbRToB13IhD++QNe1B
9MgkpyxvjBHs7eZHX8hf4eYHbby3S+K4bDBiWhs3e7Fhbpl/O1MRMvQZ8Q6K
jBf0hcwJQC5QHq+cVoR/3HhzSe954Z/SJ9x8P+I/g0il6oyK31SsLsNL1MNb
4zUBN8zDI4WAsgnGWJnP2fkVoJLOyYoMKaOUhDvwanASuyeQiM5G0q0k0H1p
PhgH3KvQuGSOIsqjM+f308Ri7l25NqtbOMIb+K9COhKu3L/rl6EBNG1Wk3EK
s68qqKOEtQD60elfyghibdx1V98Zs1A4vAvRBwC2KqnXT/1MfV3nmhRUHy0N
34yPvCuKhesDTJyzOQUwUyhusmsLneI9Py/XcuQ436jt66MJmXyXXtIxCKUh
WLpBem8a/RQhoj+jyrQ6uMGbNHxBYEXdAAQ9309+CFfUm+4NziS+NvNUt0Kt
fFlf/LihHrsSffdmrmJ+1wBhlRkeSDvRWZ9aNFjROmSxbxoAILz+vdoAS9/t
5zpHi72Lf06vXQ+43Qqpjw5cG8XB5taowmuAEClVth0s2I9zs7WW7VjPgh/u
VCykyIdFN0/+zACSTwLzGHOkkvSs/ZM1tN/+Zhy9rkF28RCO6slUB72vxV5i
t7YuN0yupCnAzPjb5JmS/N8jAJJlzf/2EqiJF/XgifeorhUml07V8Jsn1VJ6
GYCtWVSDDTTncBcFU3cMzWMnaL5bcmQ7pu9vZInhNHWuNRQlrYODKJi2/YWI
gtAHnaxVb+STyrnbz/pXPfDFHx+BWWP7LZAS3aBiyPg5W7+mpT6uC5tGhzI2
pkSmNH/CxuwPKP4g2gxGiZUHVToPCeaXTDVHkjieW6cXGBBNRNfN5E90cm+b
Zmi3I27r7PrO+aO4rRmSFpQVZP/hzBcbhatreRKAwOMr0Ry+cizU/aBsD5CT
TbDLHYtA9h6hgFco4bnlFpornkmoFL4+Sl98T8vkleMLq9eJX5TBbD5LutVW
LvO6y0KT49rBOBWyvW25r/jDoLbhY4Niocp4bZYHUIaCV1R+tK2IEfjT0cBF
oEX0go6mrRNECyL2r5Jl5qu0PzOw0IQDb8DBMZ3fDW81KXujYd+ZoNsnG2Xj
1FNSCXSSULmSutFYTp6m2fKWccg7lsMid/V1TmIXjPtUrgRBlp3Yeib5tbsR
a89Yj2AjWA05yKYbeoIdc6RCFqEbR8ejoQSwIEgButS/JGEmLdHltdON2h8i
KkIVjvnsjnvtQpfUOxVbI4iR03Pfnd4h/CrxG2l7z63+SP46V0II6CRAV+Yi
G0/VMc1dJCtqgpx/K4RhzZZFi0Kz5qkFis8eKMAFG3XFRmYd0brnJPL/5Y9x
6Dd9+CgDG15Ncx06PoAyISFFbR9mR6nokj5zqvvGkSn8bMhpW8PDBTMOHkhu
ie6rNdCW6sz22Aocvp9+IjcRfB5KVA/c3+1Q5ueqZdqnF9X4Eb8QYnN+5W1O
LREP350THMLWqJTxK7GKoug0QPzZlT7Vk5vP+e/3XrPJVmtc6x9Hnw+Paaok
5H4iBFbSQz+RbivjT0QaKYfKHXbYI5awnHfexofn4XpACrGTp3JT1VXGwpG4
tmD3+cLdY3wik6cSWzLcme+WjDksShqnGjBlsfFrNeFDGa7fVn3yTCtbN6mM
ObkzsBhKAR6dBZCJ5A6n6sZuMSIjxoATCLrJfr1q5pTSNMB/bGiQHSpOKpH1
bION7W8BeALz1bhPZMKBOosfIIlRu6vf8NLVBATY3d/IGn81dvSIxtdvpnnJ
ueu+iT9dXTe5OsZStqyMLebVQT4bk2//P9/lRRm3Pvb7mIg4w28FxnY+FGqp
x9+5VT+z8YeTZxsb4hNtSx44faja3JE5RroFwh7IKTZ/9u7F5k+XjINpEONO
lhkVrRf/AnOkIeyaeCPBe2qvfccF1fI+d+yhItwLTWOARUAMH3z98tO2Tocf
Jl2PQJ/sOGYwyRw/BVqPjSWq4zCTgw0/oZVTYPnt3F23bK/y0OsNivyAxh9e
6tL2QOQtTzxORCH9PBiODFemreFEJ/3x5YOcCmtChlpeu6CYcNvEOkbe9wmB
cdDyQAP/s+QI0xaM9+PWf3bDySdy54BrJJ94eHb90+gAKT4KZmvyJpcYq9qS
ctDYmwg+lGjC1UV0xWTN+J11OF1DuCRfrj0MktSDwFTAKAYpYaBTHPM7wff2
sa53uzooGHmgg1ePsRptHcMx5c0svUqhHFY84TAlW3QRqhyy6ad8lfsyhcXK
l5wMZmGLwTNNTKKAWn+b3IwaYuu11tQXtCSo3vJX3Ix7BAjqVAFmNd634/ZF
e6j/05xngVIcO+1pW3UkUrblHvFo4roG367F1HqYZ+/p044x48dteGs1+kfj
8EKKly266Me9vefImp2Z2GNGoTVvdgztTj9jvfaFYVh6ZD2PstnL+2lGA8Xm
iAVEos/QiyAKQYSYSaITBA7lnqtlUzRPoBEdE3kpvxzgkLHfMC3T4SYsS5Pw
OLrFmX72ZLt7HHOgu/f51fMqeONNiVE8WvLxCwQYgBEEzh0UweEfsPtC/DF7
uEHt8erxF5XvYssRp9M2FoxHVOd2rarTpbGXu/Umcpgmrz14pFvt1/+JsVhX
8ntIuN853I6SXW38bkYTV5HTXie85Y09/Sdummp2CI7aGb2uz2GliKn/FKFd
T8S0VJo4ED66i2m/KqtdAnRFDNWgZ374BGhvg9bILZ1JiMx6ohv55YuXhnof
dId1F5qASQqj+12Zm0ALMbIq4tnjMpKQ3EyKqemdP1Is7lNtq1kHhuuC0ff9
0SWumJYS6WqMAzpBPcK85pE067U6wp4rpUyJHa6xHwhRJG375MJZBCcL6yUm
F/sy5HipmsdYzlsXKTxMGvy2dCGDADjNkZUjV3YNIx63kRom/4H7rjOsbcOk
Hjbvq1bRP99GvR9rJuQDyQ06hLCJhyIMdsIk3wdALJoluz9dDcRfcmYuRoQP
eTYEMcdRm7w4qdbWeuflvkiqOo0XqbOB27nAeEm6ChxsIHRI2W4ci/at8Y01
uGPlatHvhBYY0YHzayuGRZC6JeesEW+Uf3c9e2FxZNvPhcetXERjEoBPe2JN
YewHagKS2szWzaF95YR4wXBdHXbTmxNJIW6Onis37bkFqRNCVEE7jNyNNkLK
IsAG7GNjh0FnKbAjQ7Ymot0aFNws/Vka/BD5X+Trq7cNf5DfGG6S7tt5PkV8
Uzi9qP/FuXycOCRY4KVsb/CMb03m8xk4c0kwdbn9TfaqiFfmx6MeY+E/ZBY0
ZUSCvX4XkLLocmOQOtONPSzV4aq8W/7N5PzM15vSJ4Hund9A4nRa+UFmzEdm
LqiCbD1OLTx4D8naAAoyR7gOcI+ryfyMYy9gqzRwBiegjvlm3SUTamf702Lg
ffPMNeH0AGDDfuh6dOr6OBT+ehCnC4tT0vPFctipCYJ1MV8fOf0iksR8OlLw
7ma3ACTOqvPOAApydEgVpELzwjStELtrK5Fx8jsSb9pK5Dqvl5BFYHvufcwF
MhgpbwDqzNzo3dL0wDdZiGmlbqczICRAoI5e3uIaOVT66lw94i7/k+iWyASA
j9YkfQIkmo2SM05NdYU8cjO0xnWQGmflgwdoA7eW8BwKmfWXjrtZPG90uiLQ
s1I0IMooUE6sHwZpsJrnRxVi8pSrjlx7976cMlzNzt69NLQdWVrUu+fRHQUS
+ZUItYPCFGOJRLU3bvUV7nkhTKz8OdJNCpKaL4umhXW3uYqlugHzbozP0VMI
ow4E0v05WpBlSpW6w2gOxZeKM9x1lVHDreIVr61saf9XHNvrpKuP7JpmsSR7
SCuQQMvLwFjNE9EwWgGwAsET6wbsa+aenU3+o9sXw3ChVlTle36kdT/9Nogo
h4GEXdhu3rNsNRKnuZzXQaSaHfePTPyWZmruOuoNCSUWnpRFNmdLLOUT0rPf
1eJL9+bw6tpZF2oaA9c/E20pUGHBgIFcXmBKyli2mq/H43HlGfd2LN5sMauA
48YLkMtjZlJjXvF4uNt7MI3frGSVHGrjAAJVq4wxywUmw06r5GeBfu24qHZh
6vRbqQVS9DSUORBbRAKsJ+/9YKIZTZDFKHiUWZwR1m5RAayGFRSdSCkQKS6+
n7QHi7SDTUp4DZsNLkZmY8vQ7n96jQzSr0mB4D0ypr3D2oPAOMD7Id+umQpJ
BgYRITmVzmbnYMdlXGA4G8CNLmBo+egzMd1sM5z9Pg8u2Zdl+FA1SPH3S0uF
cKEYgdemcLICZKY+Urn1CNSc1N8KapWsbpks8Wikw6pzXD60/EcYsaG58zqB
ULB6GlFKAxuMDZXplDAnLvkhZ8bv6RxEsEy1Y4yQpX0s0Q4U7/cu3zx3bLq1
sREoTKr8/FyMIWyh9nKD9i6UUcr60awQv8ewxUVs+/xT4/rzuO3Y1rkyYdAM
Ue3CkT+ydVJgvLJRg4gGKIlNQbv/M/bTn7Zu8/kx9dvALf92hnTg/+IadaYc
z4YbogEvSdxNXrkFMslkkZloQeAvpNLLVbnmPT9wQYKXNjkYjphdmwAwrB5A
47jaDsGHsQlZCmaKcoBr+45LtXppz8ym2XR3XMg6POWAo8N92ADnr1htVm6X
3SS6vPbWx9yocuj1sZNOcSBoWhUI9bW6qYthg2h4wWm17g2DxngzdA4XvuPN
Fh9ZCE4Tyu7RekceYlo6mZ/ujGZjEnhm8cyMRyg7CeX2x12Rxoulcj9nhBiI
ywC/vVH2HTuq/tJyjOD2q8XR0ePcp7xr72WtIleKn4RR6Hu8R9WEcmtf1eFL
ptNsEYFYaSh/P66pi4+b5XrHVTme/8Hz9kqPtSBhhbHNBjIqEythVAi11Arm
jIOM3zz0/YkXszboNFToppdmhbJHOEJg2YYm/3oZkvej6LDhkeqVHH5JpphK
gHniXX+irqO7Iuhv4cH3UYoI3/DV5EvOqDYyAf9dWPOjZ3mbNjtlEiWhuNft
cJXM1aIoMd2MXeGc6jB+WBu6fkg5LD6/VhPuGtjxQAwk4xOHg7R1YiO1C27z
5zCgRcnBYFZyN13vXgGA5/u7z9ASOoXM9/jSWwhI1oW5vU846zulaq0Y0DSO
vBP2B5zhqPRuFuKDqnCP6//ASif6Hqle0wL+tl+lrG5Su5hwE/f4v+wHI1nk
ZOgErR/wIvIkFG1ehyU4O1yg9A97sm/8JdeBceX4NbGUnrWJ5N6msWqTsYYX
1VeKqhpjx9/0ADstuUFgWhs46Y9eFbOxbiahSr1XtwRAdj1XGmJd08GW6Pjr
ofG9H7lAKnUTe2sqHJBBe/9MNgF0reZrDsCn2nE3KiLdkDzMT1xoRli9ReBZ
8/eWhXLdkNzSmboPp4YNldE5VLo/y617uyKWtLj/boxAnmg5CD9PNgDnGUwZ
zIoHk9/z4WFrKjeDKW+EXXDB4auaglh+wodkOl7bQ5EBcKY8iiR4JU2tOwLZ
dK20u91jZbvcu6j/70iG6ydGbjc/cW0i7Y7k4trrLVp5YLKnxQImKebIHPSi
Popu3dIIm4cTY98FLZmov6JnwLd9nZz2Zvh5Z6e7jxZB3bM3zQ/YW1oO4weL
qRFMHzsAsnS+4P/qnuvFiVlZ2N7PV6lPOu2qPTZ5M22kte79GgC8vBNhED5S
VuTymtmhUDyZbLaYJuoWVjoq0sIAkJvCftJ8DSyHzuQnHEa0vzt9ZJXW4cco
XJS0n55Nge2HbFX745kWieeLpacfAENgM407/tECZIX1LSRaMSBWPkTdDwGv
Q3dpBOn9C4lr+YjeGXl/QS8VjlaKf8LrL6FIge/stR85xUd6tcv7dT+wnZw7
yZulXny1iXHzwJsKAILr3uccEfEA+N111MqjpXEvRVwaSJlwPSTUTx44qmFU
NnfnqZuFjLNmGMyFQzIBXdob7vnJ5O/jSsVB+vH3igt0PIg898r/0rE5+MqC
Y+TgXVS3KR88qKHdqXK3cF1C99X2SNaetVrbpMbt+Z0PCYXA957SXes9RVRF
63AoBUoGcZWYlSyW/+HWHtYcxfKqOV5AjrDElUP0tlS/KzI52upUUKGzB9sC
O9O/kA2pIULIL/bO1pL3iLpc9YHNkGlrXNtWzM5H5w4wEMA/8WlpPxH9omVV
uUnfyIP4yhjEJbY8o2Y8Ey45PMEsIvDWv/QtwD2KqEKZXwtt86GzdMgWCMuz
RgRUwu3xNVGqHl9HVLDFTvufFtp3K+1ZVRKha3o+ps5rHUPrEtjSxpm65Xbc
N03YgaeccyBvz1SPvr5VmgEFk3mtcdSNOGpvGcbeEyDkHAyZC++jWpRpLLSg
2Cz3z//ue0HsMT6EVdsA/wZyX9vzOQtxX7b4gZ5gDsJibm9IMFiDdFk8BQbf
wPg2L2j80IgDaAEjFM1ahkPgq4NsuInHR2u6OWMtYtJrLRqW01zmP7oAb4FA
Fr5kFOKapc70yrYjsmlbIZn/dEP4b8elTqP1Ux9NCbHpm8k6AYPixfMJFFpX
pFDFsYInFymbtRxh1Oq3ZYNgl8g0zQbEF8tJGmmpatMs/ophaxAdok3U4Dei
w3mSwtubbQk/5Hz7I/8xv2hMff76j1RfJA9dJFTtK6opG7fjNQAJcoPRs1xy
lJXFTzX6UU2Q7rQC8UPuR9R85RJgzpavaCBlV1keYcCPjtl6rSVbZzwlg5fj
ZiL13xtX4gRud+aXYJK1CpP6I4E2IxclAmh3UINUXzTPqhuOr925EOY+2PKD
iywpM5z80eeUYB8EIJPf1rj0VlI71H+oWfdoWypDD9p5snaHmyCgw08yLAQP
UVVF9uwR7U0KXpibyC1Bz5KMhu/YPB6gWcodQQ7IOhr1i1fu7L2o22tAVwyy
AunR087C8OjDuSxsFShaTSYYeA3wkAcviFKAgL4B46r+giYjoijwIxoBqL0J
Og5ZZ8XL5k2y+pWGouxMc5ooAIcHMwxjwQipan6VaEkcW5P4TBtLvxBxjkMI
RfaUKp2jGLnWBFYnMLp9w3IDBonUpTJS6hcVNnTH8gb32LindEq/ngP3AWMS
GmOLlMsC4r8n3AWyQMRdvS/RO14Hn53zjRsihUU4JhfFS41F00sRzQxQDfPS
uTn3qEzbxFrknyT5xoIjtJY+ix0dbDRIHNAvlBj12upvJre2AVareM5LJxOh
z0KTrgVJdW+U84t7v6QgHA1higTNLhr93p24/1HBZUUNackQEgklEmezuArd
0rVvH7oCcs2GzjYOXd0/PlKtbEuJpp93C9s6wlUCiV+mNyp/S1Qtkxv3yG86
WMmdzINbCAUWmNGsO49vfKfSVF/2nLWyBCmsII/sv3xQZvIvCFKrQuaSKkkh
xEIDTLkIJdtGXi0HneQz0QpPgn0KMh/J9LLeMoZH6xZomvRIindALHYswwqO
Frp8nYjJ/OA1t6iTgXxaNheitSm30FmMkVvNZEtB8Dh0/4OibvVX0DXf47H0
kuNbMkEg1m4XdbORXXSDFRvXCyI6+NhvCOcK2Y47qAg7Qie9/c6+tGD2wP0u
7gnOkwmxkap3vkYjCX8MOk13rttQQATc844B9QB8AgGvMvUw0f8AwMio0G59
VmusOKFXVI6MRWHRSUV0kPyWuaOHRoQ7AGCu5OiQgTX1Ef17Ps40tpJOU9uD
2P8Qg6esxp1/UzkRVJEKfFV9kpZmqgcZw2gvuGGv+SZtxYftfwVSvA4G9Nje
Wbh6515ZOIA0A5jODsmRH1tBVaKtG8ecQE14dXta6zVGzQvBqllANQ4Apcmn
c0SkoOxa+vYNnuPfRuFL7Ceoj9b1VWNR/ybrko6Z3vpAL0jMQyCSM8pUnBwY
5vFoVCRg2CqJbGxB1D3129w11nJGyaXo1ARKHFYY2y5wi8xNQLqzMy+lC493
ckP/psCHmeQIdmMYGa2nmpkCPkusoxaYxaBcM/pGRh87+s1ryNhAUxOxmOaI
VbcaSVM0v3rVfT1Ccc7IQXNmLIs3I2YBCBZXnrIJKxWghZJD5LCobrn4xQR7
ZeZ/FLKXlNxK6kAO65vZVFbODlrbf4aAUAP679N/pzRqnIGYLiaFOKIIkHkM
Uvu9IVG+zf2qsonq07OX6g7lgnoWqyEkCYiIlKm00Txbk+krYobuXfIv1FFB
Yg01wQ1xO8GPs8vEifYhbW7eUrxY0JiqZqY/NSUZ8wvAdhMVvYMUASs6aYh+
xwHpQM1G5zwL51IzR8DmElmJy5cpHhWqSCoVIMe3J8B2QE3Oh654fMlA/dnM
3e46if3AKmaLslBRMcmljW0VQ1SuDY1xruEK9/lgedVsRSIstWQao7iDYJ70
jEHEw6VGfclUN7I62HumJ49aXeJh6h8D37EzVdwosjJTR3BVYwxVi19ZH2Zi
q4SNS+riA6xBdXo1NlZB26BFuIivBxvwdbHcbdlJlEXFnc4qozNwRDKQaQ5p
gLLw0r34KQke52EP8KEMSl/u2TavNYDyca5hWwaVxblmiNhiD7ChICHgGE78
heYpznZqigD2RxeSFZxhGhSsHcAc1OP/DeT/tgyLKjO+6+TFO9L1CDswOdFq
Ifau5Gj2EHYiMm5QWoXaL3SOnXrQVWrZt2aXM6c0XoV1xbzmYDL+XmHnErln
kMvUVvR/ItOMcaB5zBgPs24jlGSsvw76IF50aMXodOMtLFZPJW5bOfS0j5nc
l2eLLsjSXZzaLVMzJMqrjlB6atcYQdoq6JPnI5c/pFPyeCmPUoKj5Z4z+o5X
Pc+iR5k91BiHrUuzsQVxlkZTLTp75+ZYSGt0GNW9adRAU8U3P9/t37PdVubA
HMRZ+58KpRJB58f6I8kv/Do6bzvRzvSdJMGAXvn9XmEyip9nHurzcsjZaPaH
7isV1r2NdkYdtw7QW79149UzSzOYPiVXiXu4UgcLvlhUGPrH7jWCYV27WOt9
tdecIImh8ZaWgmZ88unKeM6Toq1A1N2fJSQrSylpDeyqtZ3VmcmHb6hebpzO
yTYhsYGQ03RePMtlVdyURq731x0HGUqBr6ecSVEwRJJqyl8Dhu3TXLvPxCQ5
eAvWxLOy4zjQ2GsxNeYYEIpF9w0IceKpv1NowDhX9LdZNyeN5Oet67FojaVW
ltj8C/TjeWA2/9UdWO4wyEbplLuu5YjVPS4dvKGMqmcnXCqx87elZ7WUlica
DKquc3tAl5cf3lMGzNp3KDIT/FiCR3lAAWuzPtZVf9/4RWRfziV4gBKagq9r
+CI1fxp/zN4GjWm89jgkuspV6m6PQ0e4UOSYbw+XTL1lLn4Xvpd3JKMBLDJZ
zrDsIAC2Ap0Ro7KhGzZhVTNQiHUa0R43hgwsym4zwkvSH8w1h9PJd/nimwJT
sWmKSRP6WHxUbPax9GD42a8DTHH1IGKnkaMSiRRViY5ScxGEyAOayH5P1Y7O
Pj889KKuTW+OmAb83jxr4nBjeOITf853HkyvlwxCDi0w2dROj0SpnGdbo0+X
65Rbt3Vjuh33T0v4LQ3D5QJW0+kEhglmY1PDYUFxvBUOW++StZhmUBhnu0/p
GcmzOM1mgPBxD9vXFggIURE/MukheFIVRMp5/k5D7eJA5PR4vS+DlgN8RxK6
lHCXMkYFGlyoy8HnNzxNXmhE1b6b7Vj9tGqmlVI9oz+rxTXeypuGRHjIf7cS
4RH+IS/ltfdt2oZ6acQ7iXO45aeuQPTemMJuzZTsD2rVcHUJxgPCBthEKmW5
H6gQtYn5PryF3yp6uIL4en7vfzobHmKI+uPR3WFoNbWQISzElLh1cOkhCnml
wXc8N12LCsqn2tJyD0y8USZrxA5tv99wruhPVEAkM+k8l38mn/bWQzB45rBc
/zJ55803VYK/MNo1tgDFSalmlhP46oDkWsFqRl9lzc3aSbwB0Ibp5z8PI6AZ
wq63w6Es1xR7v0zd8JHfQpUt0yzm+VaAJIsVruZ8NTCnVggHlDze8qtda0tx
AilFCUSn6cBVELpJR6poJqPJK5jjjseKsxWWdtx6ucTjsKeVGq0x4Csh5Sqc
q/fHnkc/emY9pCMOC8wb0M1ImYPCBqrPq5YMzbcEYIpPonkZW7SgMR6NE8iO
at7U4l95ZrHjN8EdDsWsbZDXyK0mqqyrXJH3w1rszrE8csRfQsnQEDkOiV83
NAgEIeT99tE0kj12JoBMEre4MiKVuqL1Iawhf9Uy9iCJx472lvFZaq6C04zj
y/eUE2KrWQ8+Pl5wR5WDFWHkI8+MeVaM3aVMepCzHTgWrH/TlYtO22m9o1Zu
+siM3KGLAxPYnZONywJNhJo6k91F0qVHl5/p8fFzI1uwcZoZHycipBi3SCdJ
Va7VChZdeRnIp8bMeJraqoj7MgJ7MHMH3WBiZ2AoNEm4On39FE/2SbYK98qW
H16hioyJPFUDdEbsMGAYVZ0Vpi87e/l4TMYmS9zK8Z75ghyAfXZblNmuPssW
OZaVDmkkOefVZrqz1y0ufMNlyLOen/+6uyBaUH6i1X5bEpk7VRrftQW7AjM3
NyKsb1qyZQS1N5o9pXbl4Q4HdTHpw4N7Z/FvqPBVTDUgQ6DA0Hzwt/i6EMDI
G2hmDz//qZUU/OuLPJJMlXVfsRBfqBF5HSAfaM7loJOS58i7zt48PpcQ/FQr
sdqvCWupswPwIDIAX6iwEo/DC45mwQLvy7vMKNrSKb1XQ9pYnCWk0ScuyU30
lNQONBFLimouLJXbVpIsXGl2eL8/cXpQVyZKZNnpQAUsmH60cZIbkGgzCe6h
fYILZGshB5rkQyi0sx3lpGSYO4LuBj8h0J2+xUbxdbCCkd2nTH81D5n42bgT
truxUjoPscV1kmNnakoaxEpnHCzdn7NJkUWlTmkjNFdVXjq6AfGZHz6hrIOr
YscA+rNS75BkmIAYxQ8PENraoNp6F1bcuYr3t+aV82rj7HO9fovoQzYfeNKj
oii98WZsfTLAJkN1e9YRf2SAkqSkrDspFLOMNIkOYpDozjVfPTeBVPq5WMYT
YHFXqjtTR5oUrTLPE5QjgVwB+fbxc6AEzYVnJXaaNiRkMzhaFC5FCZckzsVK
AWWzGlVqJ4QbhdOf7MJD8jzrU+AHcS8Iq8gh7TfLOdX1sizFEAOqtlE+h0Vn
XSy/pmMRWsAQvyxq1LtxEn7yuurS8oLOZCUjp2nalIAiamX7qtwWUfrVEr5L
Itn0eE63kMXraBcfqxTEW/Hd37Cj/eqW+WtLDYgHG7gF4LVVB7B4uB5o5qMy
aP3JnD8klf7CJBVZB3EOO11QBTMcz+KY3lHRlj+01ZnG0I4cuKmb3Z1LOyjy
su/VHE/4GpIaX8B8fgInIv8TtUBvSEQbc9eOjZpOKD/YAXbrSs9iJKldUrIt
y9oFuGokAfQnpDPFEtSBsUJ708iaUQZekNog12q0Abvz3JuxVAnO0MLtJCTA
D7bXIbfja9E6UQLadXuBLZyoKQUM7moUxBdGAe6/hif6N18tbeNHBYeu666u
1hwkCQyOZSubmFdzSGS1LdHtZIMIzL2pd1Jhew+r02Y5HoDPexIBKcH686Td
6NvP+ItMXCcGGFtaJI813qFgYJ9GaSJMO5rJWlBxwXa1C6m0m7E57cZu2UyP
UC2fxqQSnV0W5NSOniNO8EkAw9DusVEOj8/KnNT10/Y55hi2K6Fl0jLUbQ/Y
vKlQqgx1Wl47JxnTGITvwTQw4KQfaUgWot7Soz7vQ+HxK2/UliaIG3HJkgp+
gSDxzaP58iaUa3UNXqBzLDLCrF1eChKitUHjUCKVr5yR6/fcW+JxrSse0Doh
4SJYGvxDjWkJtO6D2tPzi/bhN6zQNEKNaobaVg0OG/BtPyimlvzt4TNBnzvs
HVQoGpP73nMaYPWk2pY0f8jzc0IExIOveyTeBjWxq0pflRxOxtjOR6JuHShg
cWcTddERfQPbFH8SYqEHfKCFUKi42vcqpdxz+bE8hNosAfGRgYo0pW/ngKMc
9ov76FUdR81O48ND+IyKMXyrSvwjgonB95K9Bq06ae+z8c6+nrxoPhttLfN6
sxrD+WxnXQFgKlUlgV4cx4EhiEaiTmRTK1LoEzT9QDff83iFLLIWh14ySS/o
yAsRV3fMf0w0Exq2ZSaqCLVOkqwz4DfgfpMiTKH0kK07aZ1n5JHet/hfavYl
kidihyT448ppizJ0eE9GM0KhHBYRvxWRO+M87PVaYI54Y5v/4QVtemfy7U+G
wQwT68fqCO67H/0kN3EK/gd5aFlD2qgb8g4ZaPqfB7cR6A0Fa2JYd53upJ1A
CKjAbkyy8DbB6rC+1ANAjzLEIUq7C2FOyhGd+hkYfoHdPsnWnlPdCsHpE2Zk
ZqwlC1wI1NTufVqNT42bILqmGjIHFaOPovULD9lIj0xuWZ4Lmg9mnvgl4Qh8
a0jObjxPQGFSUO7rS1UV28N3Cga4Mh0Fx0Rc2SCGyhI8A8tJYAvRe2EMRtP7
6P6X3cPgKWMfWOWnQKbKqUcPIVnIfSHyIsMSJjdcOr3psjCXMpxgeIlrG2mR
7ZxDHCzRxGA7RcdLpWrQlwyvzOqznxaQfPhXxEJ0YUKXVZWyFGHixyVfm4P0
8Kdwxn79Xp7DZ7Qm8Q/yZdJlQUNw0eA/xiyOjmFcVj/UxI5a6/6akLY5sbmx
rl8PKtyOKZawS3gHdqpCN3SoiHFKkBWun9IuLrpAHQTRy+vPesNwaHauaCNY
xYmsqacWrPA5oAd+Lb4a0NmaEAVNSP6mZ+PfPTgF/yNF5FInixI88oZx2Jbb
bdihWPgAh4yUF1Hz44HUsilPAEH0F4FP7ffPqNX5Bf8OIJ9RN4cH6spUT+5Y
njVVXV0+ZKiIq72fe+CXfuSdEFq/yrmeFlsqobdZ93LeHtb2vHKth28gty2R
NTOr7+TtaxFcrQBAGJw3F4J1Cudh1LCdKOyG7+L77qJXYzOoQeHW/dSQnFJE
cSteWFsJllJ4oEGeKUzfvpzkfIAos6JUQGgVxkEw9jnIDN3BJMxfZ3pefb0V
8iis5f2DxuCs0ibRwOXRa8dOKwcgKqImcvcMZqUoa2FvBh2jeGWe/2W94O0b
zFGN//MaWH71Oxd2Jqnjl4V/u0BnKStT2dg2hhq9wEFQ7XWOSchDHhfq9P7n
gv+sjU/XnqouY1lvHoEK8hyWKb/TlZWSJBwaafwTH3sboi+6Rfg2bEggh9ED
T6D+1Oi0Mp0ySWZNEbeJWvgWs+vdRK6gCTOJZRqsiaO7NNYbDNIfk2wCTEl6
HuvjaVnKIfb+o9pM9DtLRMvRQNxU0Ww6lF9jv1aY7tjzhvcY/mKObB+soGTW
eJSAAsTq9RzsF+U9fXT0COA9mgLdBhXve6ht5Z9LvxkONRGRx71s1o8HnxB3
T6rFtF5zxSqBqwWbeVofYdpqCBtYIudCU1OK6UajX83Xl63k8SSKFm8SafSF
pNXoHwsKL3AVHybkqXQ3qCzUhKUk0so52eL9a99RFKTIUrzCovrbu1GyvwQs
4XHH6w6yO7bwI9nAAm9QnDglqUTWHZF8EK9zYUrwCAhEQFQ/w3BXWPk90Lmg
nZY1PzubGsYZ/PbJ+8BvC42hQiRfpoc4Ljl3q8Sidnp8uUEcVGp68grg6Eo1
AVyYCpphVHkojBtKHwgVMH3WoSj9ja3cQoiSTUZ93u/JnJSpBWzSPo9hsLts
64ihmtSCeuaFQPsJf5S86BxJmP5adXgjfviXwdaF+q3Jhr0ryAqpF0RxWWbW
tbHA+StuYxizsBYOAGiAbJ6qWJkqfBSLFab3OpnstgMQeVtx3LRyh9kdZf54
7ub8Xmz1XMtupHggGpMywMis7TNNrqxwmY74mVtIxdvLBRTr4rNjdCxqLWxY
/PMrLlStdXtZimju8jm3M9qLECZzmmoIsafqsjm/ItzjDYwjhCzFkFXNSNmK
X0ywJYnymJOY0lXX9BD8qeSYw9JTZNe7HX/dYBmJ3z4fEtbt4XyK5bDQ2nWi
THWH8KbQX3YQXiuE/gvLfYGbsQUcAIWaVvVEAXR1SoGo5/2SbngveK5rUF1O
3Ir2O2iA46zyLWqeEXQFaPj/h8dC5PhSnCR6NfxcBieGLirtOUlBbsGvH8vX
htktS+gqq+qUxrWUe8QURsXQWQoolYSVGpb14BedxSbxCV1gAXHpDUHUASWO
q6SzNcg+SkijQtiqmRXdwtTyQXrZHm33KTvSd1g7wjLF6cs5YzRs4wVDyp+L
SF1Z4gB7u7T/Ldx3QBTZu3GcwCZgIYbqr1gcexvoOtK6pVnbzmy6D4AM4zva
l5j3RsK5XTNsr9Ce7oc9+P+Z7LEBVZ2HdatcHhA3JB6KTaoINar4brBXKFCV
BLg8DI8fYdiuOkH3knLn4tY1IH3nhCEhlHUT3n8Tne2c5ocbqsyPPfxtVKFV
1fhbbS29s2IzYFnjMFIR6dUmVhbXwqKYtfQvf8vzFte3ZNsmDjEyKbiI+/aK
ETpDXewIB5Dm+fh51xEak6DeFq+F3wobwBCD1pLFYzsiAn9DngbsD76aXnHs
po7pe+gekMifKYw8BLypezpi5ysPS8/9nM8YGqp/J6MfVgdjfgi8wdG45SFK
bHZTzP7nYOqTIpNFRnIp0kQWbdSKhCVj7HYKW1huaXeRfVqU7qWrWzkT6Qc1
szwKc8ygGC56mXWHudmD+Y0CkyhgNi1p+cizbOAcCdr5zh4wNouuhbSKr6MB
YvN9DhuU0q+WFQk+crdSTwHEjLe/jauBdJRWMHnAwE9nPPDdmFhBA8qhFmFp
rgOscvVLyDNe6+mhi5ylLwYoal0torszrTgU6HUMa5C68fjWD56GhYzwM3SR
KKF9dtTICw+eDVMaMimK+oK9/kj6TO0CsI4gxrDZkCr8Q6jF8ZrgyL4TjNjN
9G8RDoW8L6eO+L5gOdRn6hKMlvEEV0TfopCcktbxg/DHTty7I5+z7a13S0Ce
srgfXWmrzRT9TxDatrvUPdCdZ4o4OB8esZqJHhrtTdp0p3IdN4dPvKN8syxP
BlWFbcYikQZ5wxm102yQagU6iBm3uJAWPRB57BFFhdjryFeRvQXj0ghxeVlj
pVxxIftJaeze+GUUKc0ZRin7OSdGX4vfAS0u1DxXw4MtS9PiHZMJKuaORzDj
iClcxCobVkrcS0p4F9Hj4zlHc4XEPpXVO8XWhSY91+rg2VjTkrl0NY2eZncl
ZN4sDjX8Zg1OaJHpXRKnEOi8i6bkncBdOXI5JKXnuIDihcZqlRSIIfm/rJn6
3DcWORCWoEJ6oa1DN2MNMOB4jwI/qT7RuvKAVegynyPFeJvrc1bib9K8s+ao
lIAhiiXahTPoxQNMf3jzNVk5x2U0HYVNn2lugwuurvXc37hyTNSvn3frbcQD
RtdnRoX3+Gk8qwfaBErceF9nI58xse4YZCvXGa041Vpvlo6KIKLd8cbaw7yw
Z3ApHKmKkoFg5XJCLhqZLNK8sZmNB3/uJWKzJdPu29P0VX8MGZ7sx7jIlviP
b8qoYqWiM40T9qlPHPlwhSjSNBUNlMNlIFHFv7ksZvul1dhpX+Rai7xUOlzc
WmOO+/dXqwtMBuY5ckJ2jd1sSKZ7sY3WxnOeI4O8+lv6OkjH+N45wUkeugny
7OaQzbQNfX4kb+01QAmKQJdWNY+HRmK55Uk5yN5TUUAUJguBQ4FuH3lxCAU5
AInMZZe1GTwW+eM1ieznRNhGCqsHVRQmhxJoDCpRKskgiz5G4XQtt+kU53Ak
w17bwpeY4rfx77MVXYPb1PXFsIrXNyTwDvVqufiyxu5HUBG409yTbNwCK77R
ao/MhhFF9ylrZDWxvGNO+kKPEiHK32FDWNQgKrJ7IOxQQUoHcEfEpbVrz6JZ
XKQowiJKJBeM5jD3Qao5T3eZjYUfsTWihGM973Zku5u68inO/14CheuwYttA
35HNHRsxXs6YrJvzWLymeWXjV7r1bXF7+SsmuTShQYO+/VQJiplSCogH/EQu
FaisSqo+t4gLn3tJpIGmDa0+jO8ZOqBOFh0aRUs0h5BaXzNLI2mB0ij3S6zG
TS44YWoiJoNe+gpCjGGS5VRaamNKpi2M/A08Yn+40iXankMWx5fMLXrSMXG2
vxa+5w3/e0Tr/Z1G4w5gIzXy++PWxQhcKwiZb86V/0UydNZL9XWaKqcj4TjW
ArM8TeSk6Kv5sBuxkWqxYC4Hqiq9oRMtK16OgDOsn0n/HA3e+XUFElX9zhEu
MouL4OxHUMMVJT4SI1z7+X1ZVSFzdrUxiP5a/ciyu8pjck6mYRo8rlMENmeF
SrvNCEukzHfqGHs8GyjqoR02ewgyTf7dsdEyB1reRUzKA3Q2ZkYBVnUOauQc
z4fNhIaQEP9uSolTK2kBTefyg0Y+BdYkcL6zhW36suWCf0IfmN2URMgeT02c
TQitW2DHeSVb5OXDOhEKJtBndZAgVMCDXskCkoG4DyorqEmlh5tPPMub91eE
qVt0lftWtcrS+26egeS0ZI0+2kuoTETZ8dEElB1DapYCQwJwd9x6BQ15yeZ7
fvKLt4vHSYQ3oisegQJsV4lmJK4Ztuwym4UYv63asvw8De9DUC31Ulg5qZka
M2CcDCcm9qhxFFVtiBoiQcRP+9JNXyPZO16rnmapZd7dArqeBtqISCAFKz91
BZL2b14vbJafsR8VbVOPTjvr+ioOpDO6xf+SnghzGamDZR4UHHn5oOBqOrxs
kblOe7n9NDywzK7mNUPFBu3W8G0zyH3mKDmfK6Yw3FxiKuXMrM6nHaQMXVAG
z9YGgzlbYwZb6nGoFrDgbG49ejo1OXjZP7+fzfS/3SuuRrQ4cIC0H0r6lLaF
i1ivr8Muiff+6poNuwdX5m+6bfBRI7F6Kmz9Wu7uUsXEEPYCYGWZdm217PZA
8na+6QnICMZ6hguM/8sw2fzBF8OVJSB8bp/wQJvWqfQldZ2G45Yy6e3W6NRN
4ZYRAENpJG9Bn47sp90Rsp0SjZYVkvH2exgBhwLqMlZhYzS/Yg7NB2oeiFCO
O3AIoiedpsbjamdKuzfcN0/GH3zcTSpIebSjo95C4EGt9SgJ+/qvCzYm2bmq
02Mr+Csgy3uRBBVZ+MtaLpO228qQLg4LCxw/DbgYreq5T9DUQi4YYMJAMyT4
11WU100SvisajIfJ6gD0qLuw57i0bLD7XjoSVFzR/kLAaLoVQ73ByxtX16Z4
Nfjg+fTot49r0oZOop0fj0Kq5c6BgCVOdYMWxJIdQLCKT0np0DM8eXQAt9AV
nWwdF21HEo/XAT0cT1eqf5Exf8tHeX9lKLUzQAM1S3fT9GUPJ3B3kD3ltsIN
TVGi9VL3omVu2j9OnG6Y3EsRyT89PXoTgBXNJAUw3vYT6EhIYKFmlaYA1/MQ
pLEg6dxK1CDN+yT4iRXHaDT41ZrBUZVqdS+6OKgu2QfJKXifeL+u8BW4fHIG
oemkfRnDOPCG2WPi5gyjWwnnpv01mJMkRT5nC+DAPMW85TrqZZ5JAkTfC+0k
y0tX+2Ikzgrwy/xRLjfZMGPjNBb0Xbqfm+05L3YMUjQh1OG9neJfC0KrdP75
cEik+tyJjy9z3IyNUAQVh/KMxGDWk6CMmbAwNSyvOFd/3ow6I12J4FVc0M31
WiZZeprDY/B/U3Ab33RNi87B0Yo/FBeXzBtkl7jpPhAl4N5Dxh6iNdmGFdw7
JXKe+IL6H3bbqhzL5Te3rDASdP69nJqU7ktNKP/TYU11PnB3Iq3em/KZB0Zp
bItW64dossErOUxen1Xxk8gkpTD01y49in5fGcoLZufCBySvkTkdjgMFcz2i
h2WGrqmAfF30pICYIPOTL3aoD7EBpbjGTbMLaYCSDxlfx4nmSDve8t8HsGre
Imh/7wpLjZdsZBGKaVG5H04sYeSah752cn+Cb8gmXsMqcCJiyu0TLLkS9j73
YrhPlJmVE2j9mfSP6A7yiNVVAORFi+Ashxs+ozx+U05IAMVkinGTxbphx4zA
Fsziu28Y4qAZusVj7omWGzzeTLsysJ2dIklZzEEa77gvRkOnESgACmuG0gn6
QmuLEJmLRBjXyHoMHFuTqyvTbgEZ0Rsdrt8XVBQn/9Po/YbdlKkm62cogGn9
ZVgzGaiBoZxYIpaVg3EGGeYAowL41hLaw6qru+W7wUcwsB4f/P19JzMNDT1T
eJaL4hXAQSHqZKxU2pO6ylZBuM+4ghmBZUglBk2tEHC0ZKKN0AP23juf2aOt
1CVL6MbE2MBKW1TZfwZyyaYSIEEoFqqA4dXxmcRTlfCckgehmbSSqgoE0dGn
dLDmHquYvSOCU88aFgL1+daELqyBpPHDFkacVTGIhZcdnyO8FmLRBcyDGjQd
mo6kQt/g9sa5PuNl+1qWJze816Eagh0Z4ZO0yt/qUw5ORr2C55jTVO62CttI
zGuR8IEkZVUjVmsxZX9x2jaRI0RcjZB/Hu4wFi7Oy9y774V6vJRG4xRLqKZF
7jQs98o68jCW8mRBsEr75v5MPSkI1V9xib4oF9lUMbGiTBbHicrE7adV4UN5
V/fy552MwbWhHeTmL+/RNfIXaKUzkyXldPwO/6R9ZJeCSD9T9l9OjB5eq8/U
x2/xZKjc+12y9aOUt9TuNJYyVJsBsp/2UyFX8bylnCw7k43PuHMhD+naZAEn
vxya+N1dkdAQEJ3PZapip4MeJRxFld6IBXLobSwKSSQ+ZIDbgMIBlVWsCejw
vFySiHCwGZLeiKz5Z9nEBw92MQ6lseqT3kkskpHSKZsHIBSjldJ0nMTqj17y
UNaj1LSbP0I694giJJzdinwWsl8TDpp665vTIeaH0fArbJjNooEpw9ZcHoDk
ZAMN8sU+zVmjBKKm/oZdNKLqvQ8YQ42vS87a1MMDP4bumzwsxT1Qm/kkxr2Z
hbrzNG/s36opGmAlHC8De3Lv1eTcIBMUq2YRCsJNHwCLA7vhvrXZDm7gB7lZ
HkaYpQ5Cj10Ztqwqj63H9KqFrSibqBlVjTUJXWv9MFNqJ8Rr+beZMNKzpgPX
mUkm2m8u028xQCoNPa8skXOwG3dFGykB0flKEpwSCFTK/DUZC9TatFc9pMMK
UaQ6JisZcr4wUMouY3Z8QnZKJYvlQ0eS6fvIu5KBSFQlnv7Of5I5prrMNL2R
h3JAybsTykUQ9cElqHxjKoW5i7cFvzhIafFW6LmTicoSNmHGMPMTOQghzGsR
JfXHHhYj17yj79NMXYrODBDKd7WCxbG60fqDjfUBteHbhoSzeb991p0vMmZs
eH6WLOFtvg6wG9whpjbZ17WFfZ2NmXAraHpx3gEs2Kbb322sW5iQvHV5peiC
L3rrHUHKbpF+R7kMRtbzl0aZxUL1U9Y5eJYeNbeh3cKatF6VKwU8PeBEPGL1
2KjjGPmWEL/YWcsL4WFh8jNbbumOzbNQeMoyvSQpdhPh+oTMiFJam7TjFmPI
nHFwb2eVM0JLuJIQmtZuRZenXgEocRsVIm9dJ5L164IygEbQoShFUT87w9NR
xBIBZhQfGZz0EXnTw+VibrnkVI+/L7Dt6sMhdtcGL/GEipGKGAQaNjfwPvS1
hTStisGpA2oWKHGmAFWWFhiCWW94IntxOcfkD8fjoMfgfb2H2PudQi2imD9Z
FUiXrUIYkHeO0yByRjuYV/fAG33IC4Kwr7pREHcKihYUOg373zQ9OI9z0Ibr
j/jFktf8E6+th44D5B45wA0OFU31IVVMxb/ZU6M0ttgGYNeET3tcvViOFnoD
yccZg7d/Ken47ZjZytZzRbGaoUVCib5J70Hh4r9Y8qwxxJFbVwCFpkewc99l
zmqTLWMDRiy47yO7mgXU/RC9Qh8vCpJGX+X4t6O/Cr1Rh9Jm7E6GEfJolHQd
8LxiUVhrwv4gAbQ4Rajl632hSEFbE9pNQr2sLa6OFKQeWNMsTAF8BLqHeXjV
fKwUyRjsKrX6VbL7KIzf8UI+A7KF+Cs1xin7eWMGdVhMmHyhtwqpE0FO0rkx
D4GeTTFqiIO3JktQ18UFI760bvo2BpqxPSuEmC5pyXiRHyHEeODBFoojpcXi
h8+vQiNQzTGN1vLOhsTUHLrWQ1aDoPl/+8g+WwU3LVO9nCq6bTy9zEA0oKMr
HeW0uEpA63e+YbeL89vS26PSFoqrw9YHeCX2xl9C3XSUMoicHVEQ3ops0QJP
mCA7QWKO6ehsksWuXVwEaKz+Db0EbIrzM+mUEAyow9iyOCfiLLNZ5H6BWFFG
VAkoC9VY8SQBV2ibzt0n2WzL3O3hTPWRHmyghnS3c+EodJSow6CQd8d7aEul
7JqDgHFM8w6JOtao+eZae+FKlas6vcG1uJbcENkFT/gSz3/38RH/XvrJb91H
nqE0r/alcxfix024K3jmaM1dOobIxgqczU/r1mYVdW1t6chS5rBix/bTajWB
23b8GTV1adaVTlRCtgJoMcPmJUqfeskJNv1QEWUmj4Neno+j22UqF6w8txT9
WYjdSkmtU5mqxM9clwxulxbXxs/eFMXIq2jaNfTE+Re8QYh9YfIU+w8vcDtp
gxP8vS6LM+GA2euJekmXoBbNJcNfXu4EEQHYLC8Qn3Xy1wZjl8Ht5GNyloPE
tMKGeqdmsJjGIUU+iEg3EvhJGIifyW2pRFMW/sxHt9kBnYz5lNhKI3LW0Xyb
guravGUSaGiSbn+6yHmyF4MJo0G6vjkX3nivSIcgJ1wXGjKO4Qy/JSwymSSm
+G/w+9PfeFf/ssHOq+ZfzsKQ1VrvmNKqPHE0gkBgsWWUH2NBB61faESZH6FK
JeQPK7a/YGqAwhtaON/HsZuEcOow//isbLj0313RlYtjCc2bd6axmKLv2A3i
sNKUeupmDVlemnzlGueXyzrW/XMloh6Ge8sLFl+MZ4Fb6DlOszxbvGy2IHv1
aQkth2HRSkK3WcmreXQGGr/h6aXX3NTurwnGdcaXoIP46XYH3BPcpbxzXIWw
SIAWkPBbBEcMF0ahKjWYoXhuugPqcm84VDzj5//E4dw/HpSUn2bQivRGAfs8
V1W6WiuRN0/+E16jOUSC2n9IFHbMRDiN+WkVURpiNu/enVC3iyURsGexCyJ7
Vs8l3Xw6xQMhTAzSuUM3e476GrMAit3FrDt0yF031KIZz3FJoCousx4GG7Zf
WEB3HwPyqMyJzkL5dg7btMvl3MIzNz8QCiC1fMd97pDG/I8rh+4PAvWO2ZXP
CEl71jbWy10KSjLzuep97FSnYcsExoTZymLKh5WlynJ9uVKiqLlcylzJXtvi
hFJy1JFj9LRnpFIfbl+1gUqmpJeF0HfEScHUiAVZapnPbPdTTHZM/qZ7pyhi
aRVsK+OaH3RcbajdEDTrb4QRw3pjrTB4d4OOyyqHq8i1xXw09xaDHjbIghYc
AO3uBYZL0Geb4MoDvz1N+RdySBvAcsJP59toco2rBrjLm3C5qmjrOqLG8pRc
o/Jd+QaO94mt0EutdPodq0gvj/RNbvca/jSsrD7IlQgvyjLpIAG/7JunNqMO
zBTijyfK3W+1h/k3fvCxoax5Gv0PVvTyxJ0Kjqlm1fmzfXzuR6QMDLNxyHOA
NokhM11/8fwZBa5aciDIutIJrzjyKnoyCiS51QWU+DKy4T2Ta5i+aIaXcDks
Taqhl68jGsbQFLYC2n9SIx+kmNa8+QOKLmPMAJSZmmPcVlWXy9nIKiq5EfqS
EpLR7f0TMFUe68T58jR/4jij2j7Xbo2v7EI/VlGIPZU0DpoBFbnMYLgyZ+HM
g/JPQjMoJ0ApVsWaEfCNB+8cNezBbXxHuDoOzinj2qZFOOPRgdOP49qAY1XY
STYGIHrMOw4hZTfoYVeKuDIYsIQ8U8xgwFG68hK84Dv9rxGHxGG563xlfFsq
BjRt57cYQfy8qRhpo8qhnjIytrp3JcNNwSIQI1+BOG/P2EOcDs7szWcgoX+3
bn2RZrU2qRzFHpY9VbBWCLrWfkkvWWn+QCl85k1JnjORl3HqTQ9a+ZKqdLGx
hILqLkInDJyUUw0g85CQhufhrPyP3feKeZRFxanSsm9ZXgcQgSffdqHMhhgk
SyQRkcvK0IO4LQolXur/t/f7Fu19VBjwrUU2bI8ADUUNRQb9eJlJK7sEIfZL
hLBwz8Yy06TNLAx4vcfdDEnXJO/Q3tAMUG4vhEzB5OeGA6QiPpVTvQ4Eqr9v
1d0H+QvewdabMilXATyPoDqvG0VDTosLJT8+jP7wzwm7MW4ToIYV04iQVgvE
vcrnPFTFhauMGBF9DfVW+xrAS7nImrP9z1kVbHpzc/we7Txe67W+Ck1PGRxY
rfkDl5o4+mD7ITFSSiNyKzZTTvY1cL8GF+Xwnh1UsBo7bn45orARveWcbKra
OIX/lK0/uHYyO0PqaOjxlxenjvuGumDOKaTE2hvWccvwvzJq80j2QIj0NqY8
YOy03O+0TMIUre1q13eQTF54RMuHXX2Fsj0emfOzGLuHXuzZeEFAo1bPyrG3
gvB81KPXqIfz1pvrvO7RQw+iyrTRpmtyMK1oqsXdeVTO4xrUdaJw1lwFKNSM
wxipiZTWHXaku2lt4hEgYmas8wib+TNdTvXCiD5Mtj/PI5cZwFIgjEYwv/aM
WXpIX7b5C+Ijb4aFzYeIE4uwP0+s7oRTN/hsEgRBvc7MFQdcXvHP+HANcbsN
bJS5B1OMjuVoxaSh3WUaJIemqeinmBIEi8wVl7oKwWoXf7fZCWOgjEUuQpXk
5j9RQWXwA6cbRExAJyIVYWh+Wb6inUr+3wSpzrXdfhVHi3gDguLr1UKty+Sx
o9uUK6B3nXaWbC6PLD+toRfWTWmCMWkqkUJYjn2jYwAMlDhcWqrkNEHGHNb/
MbFLmRJWLXZikoc8VxNPdR6bapG2WAjhXbKKZte4VZWQcswBFf897ifyhq9i
FAWPqYGl+5fsIV7EhkCkOE1lz5mqHaweDC4nH3jwCey7lxJW6SjItTNHtsJt
dNJCz4p4sbkc43HpqN5m+6PJ1bhC4TvayamQRl0zW9DCbbBG/eGaxg/yJonj
/zUpspdI8+ruCuAo3WTiDBqkYo+vhR0VIg6uNwrayWMpfMhzPH+/upL0Xv68
9fe6Iub93fnVvGQDYnP1MAjTgECo5g6HaUGMN2XNoSnfxhYo2pVH/8Q7drZK
Bbd1ed35sODAXUVJrIoxCrm1RdFpYwEoIP+YUvTqy96z7JSwjrVYu3bNLMxI
VAtVIJlrBUmtzjplk1lYYTx6yzjJcPIjiLqD2S+Y0SPvjcxAJ+9fmN8RLVZA
7I5nuFphBQYMy5W6vqJpcW1IQAsXvwp/CfRqpb11hsFhRpBBMkehHWEcY2Q3
+DO7D6wx2h6b6h/Gexwg1HH1jCtRY1dEpSgpXFuYNEqP9x3AlJPku50hzbNC
4SzBJX1UfGZ18VqsLBEPEcClt0mZdrIxopCtBrxndq8TJ94+uzU+bSaVm7GI
F1FWM0fAzWzrL/HyBmETVu7NXte5Ivz+MzNa3fxLwpBnSk9P23r3+mBKyly3
XgOKP278dGnl1WK247kgGGaRbqFT/8HBSN3a47dtsdArTt6WMF7oj9/bTnPB
OpaQu2VyuLIrn9fT+Zs2Gwn7xikmml/oBi91UVLMzaNTaoJww/QQQ34/xFl9
CK+A40RibDwprytoyH++/F0eU0sS30+bKHWOQaz2R7AAPLzR7zQ1CiymQiRT
gWxvXccqdeOc/s/zVPeGG2ETpYrz9lLoRKVaeMPArdOxaNEdcNtT52w1ablN
DRy3A2VKqm7VXMs6c5mciiCRXfOHvD9Yx3PjuGdq/s2uvn5MjW5urOVgtI0W
CokDZiwQ6N0XY0KS1Q/ra1bQ3Zgy+8fSTw1Jcfzcp1mlW0zCHFkzk5XbpEtP
/7aclXCBszEmhxK69NenTDdhNTO0L4JBYt3+wdSjr4nDq4HNxXMfe1pJkukq
8jD2dWwQD1hGxNFXqVIWeLizkCR66sqBXkrQowx9TpgHzSwV6tDO8islMk4B
rjLtpleiDudJ9czlVz/TpFRpuh0hibZy6w+W0rcQivt6X+xcxVdNn2D2G44E
jMWKLP+uagTPcGTgF3x2FhoJ/Fby5Wj/iFsPA9eGLT9uFACGIhw90nO/XcdB
QCAvFlRhdNLj+AKdWezCXJYkBTNwkUe1eKLmltqKx72DyrIvkJz9yFzQO2X+
UyixClVxkBt3jAXyAqKmc3aiXAxqPVo9Lsl4B7c89u/gz3imBh46s/u8yoeW
DpoBr8w0yrB+BKX7SVcXje5FmWR8tkNZt9ouqQb7h8mpyExdLELxCbhVWfU2
DkIM+M3TfE33quWctrk++p96VvckInpatJF9DAODZ7qOWrsx3PG8v5w7AuDL
zIlOEJz39vkm3wORg7bUkGc+6jEMU0T9+W6D8wUQajwH5qjINg/aS0ZpCS4X
W//AU3LiAal+l2Xh0Y4Jrome0hXiqcXMQBfqzEgROwPG09GhPPUSiIczj5MB
1F8+zkIKirzAb3MWtqctTMqomA62uldKRhEIMJ3J53mMvSYp+Vi58ySDmR+F
w9hjfZ9GET2kh50TPtx27zLdS5uP9gvrjTkO0thVVOLyn5aGU4CdE2iKoyVP
Vjasad4UeVNhm3YgHTgS7eUp2QEnoxg9F8XBy17pTGZYUyhZVHM/v6hu3lLZ
ATvpb///kEYTIZ29ZXxBOAYx26ZesXRn+oD0qGhiw1Tpo1iPUe+jup+XJcLQ
NnyFTGpTtWh68VL/vbLMNs5bYHj32XhG8eRy4ndyCVSGBqvMV+8qovLZ6wBf
loyp7RYIEyyO9TM8vTnLVZ3ATiZgula1Kg1VRqtZdl91hg7lQdbQp0GQqikw
x6w4p2P0zozfOBozue9S4GOpMpITYfhinxfAROEx6fr5cCg4EEc9IeLrZDEj
YuJsAMVPXNExvdLe05fqju1F+Bsp1iRw6iy1sQCEX5XnpG/LmFrOSmDtWeaf
Be/+D3T59M4I4jp3+XS1wwcystclKelPKhv6tDhUIIz748YvhGNBkuep/qCl
wskSi1dG2up/f1CSguiaWfT7w3gnXN/w3Q0as7J8kbegSSTeKvjFKNVXZlwc
lzHd9oYQJMbbGh5QhfZXa/x0J0pD5jpagf8Im6eBU+dlUEoJdq4chVqOIBAF
Z6Ad2jICOLEDsN3eel9f52yOmBJ2DygY28btkBv3oNIeTMG9SiMBQhKPqmCF
qmE55hqWEN4soGFSe/3MrAtjtg32ZCG3qcvW2X3ooIdh1NetQkJ0f7FJ9iX9
Fu+mu2adV+9oxtkRfJGpAAfhwTvQY3haM65kb6uIVW2MF9r/6MAU3MVftlJV
VKNZ0XJ/k4e40imbiITDMFTBRGK3aZxeUa2/5/y5diS3rBfIsV2jQ3K2M1z4
alX78+w83+FgvinRYFfPaZtMWZNjJRbyGCDchWQ737Rz/gLGfAtmr4pe7DQW
eX6s2ZXVOAi/6CUXOq8dQre8PuuriwmrMrkEH2lB/skvSx2Eyzm8fx5xnZHS
918tCIP86A+BwlpZjb0OI6R2WUYiRgAKaO5GTkCxwG9W+Slxdax1iqdm3Vm5
wUXxQ60V9Rx2Ciwcf4p4lNS19YwPmsOKD05bIBWkPUHQvxhjOHNnnbQut6/m
OCJdQqBZqBCh6BVTyY6f8tCh0rl4Rbw4oNOMZlqR4H2PvVeJYW0VoiDh1WBG
G+KJE8ykROseeaLrxgRbG3R/7w2jJG6J/dt48DiAokIOM9h0GucwVcNR1yvn
mRCqunLozX1QYPTepT8qb11V7YLQYVRQzfKQVWhUINKF8sDGaxTl3cyeaqtw
TWqABi+6VsAfJrIsPaK3FcmEILGxTgW4pAhQzDInuxsuJ7DZH36ck7yjM73K
IsBuHMaIZvu6/S61pPolXII4SAbSz3dZfzWD7zg6TtFIcoqgnga7MEbKIYFJ
ygNlDhthG1VKQXdigv8xyb1fkR8TH4BI6vMYeboaoGUWz9OTFDkoko7dhWoI
30V03Yxy52TtykU4J0pnusFcdIP1tuLg5XsR7iPf5xEce116neY8zl5y2S1H
QREbcZSANd45tWeaA1lIggSkpNNVYjmBLRBeAPk1AQLrVvInQMCuvcIg/miN
eas9rWaV4He5lGhnLWxtyER1EI/eIRxdTeUxA03mgrikDobkAibSg4YcNbM1
g48n4qmPK+RAFWuGWwxWWqHGABMBwf7324jxW64ogUU6gANRMN8H+Qor1Y6M
W+JwDHwREvKrFUrREYQyXPAwh2OP2moRTn5iH/PTuyvr3uEVOKbdxLlJt2F3
lBTLnd6pFe69OuQvakk/UpGnW7iydtHxNTpLWMuCr+w4NmkTGG//IJoc+Bpx
HHxyJEKAa8dBEmlBBc/YGAMArzzwboWHD0ObKkfkZ0TttIq4mjQj2Bblqy7q
vwaipP+MWP/6iQWqeRn0LjoWByhe1mkTCfWcOmok57lrwI3fYGE+ZYF+VsK0
L4pqGjVsh3wdYZSOzHlBlTdiIUistdW1DyCttTMKYm1T1lqt44iMXm7EzwyH
a2oV3DgiBKq/XtvRH0uYsf31M9GseAtCF4/OIVmdhI2a4LJgkRMS7ntHe+g9
AjLFwNH48tvlQTj0xpimHXausoeRIj7Oo8G84IddwdGPaC5p9DxEsa5OVrar
kQGK4yRe5VN95YD/7tqxpFmqWJTHDNL02uPdcR0QRAXKQKFTvENQMhsUm0uw
i8CtuJHefCTEvI9WkaasT1cjl5jzVJOZqslwW4TH7AcISLteQi1FwiPntru3
DmnreqmovmhyHDeBxmxZ4e7HeR/mJV5thGkMtfYGV//TmqdQ8EvDColfYJjx
Q9sWYuf4vDojC0TPe7lESJbdGxB0dCelagZnJw3/A5W3T//PtCC9bTvaHmrm
HNAG991dn6SuPTSLDWQpcCGZ2zZFyDIB6ddaTSQejG5u/31qYRvAos/HGyji
UzxCAQ2Pp4DU8Epj3p3YeITs/5snb0yf2lLegz8MIuFl6ck5Fhsy6M9oTPmY
E2QhgwjSpRC1wZgVtmhyvTrR110nzwxEhv+lDudih+Unx5x69bvrC77A4ooD
4KJzul9oYSM0H1d96c0I/ZptWNsPiWngqkAc30aF+MIUJfK0kEaZiUzWJ8cP
sEvwf85cxChS+dhhlomV3619UHtqVlNUtt67T6G2p7F8Go426jmfSwujEjx/
FcP6+t4IgHtVuON32RUk3AvPttfRhxg3ufPjhLim7tJsAK2AabPd41x0/2ha
K1ZjKqkwY+yM5MQfdUIIJ0zjmgKGF+ZJ6xJ5Wii5H1OQ2p/0SnJq7S73pH2k
ndL1SosWxrSRVJZs28rBvDKe5GMTgx4IpBbztBqOn2oTHheD/blXhGPIj1ua
yMCY3PEp83QL7YkV0tA16q7xRdfsqT/X5Wk235kyykZ5CJm/Xnt42TBd4x2/
ovun0dM0/N75LTlaeJsG6Og8InYwAxuEatrpXxn3YcDMJeQ7KNpe3i/cO4sh
LzOAm0H+gAw/QnCYbhTr6QdmK85SiJ7+7VbJnkEAthLpTg6H8fAmnNwqTt5n
F3L5+pJwGZb1RXLUp5K7LtyMroDZ2qqmx16ks1v5u28wdimDbtBicEZSEUt9
nO3WVWiudhWNVsb7TvdVpjPNra7jcxuVdo1lhoT2TTP6OZgf4V4Fpx1IguN4
s/FSsb1gVDkgatJms1dgQRet8sY/aT/DcS80qr2d3MvpWvn4Ut9Vp4UYdCeE
IQgq0ZdxFEILLpSf/kx2SPK3fKB5ldNWE009Ibvnx0MF7Jo/Pmoew7Wi5fwX
z3hNgU/2UaoZdWSvho6VqYfxzVO2O660FmyAvYR5eeTpfJu5DGgIgHaE+OQJ
OwFWLqIpJUvZ2BywJXIM3dHcYzbq+QJuL02TGwVRBo8EgwVE1u58A8PuHmdN
yiaaCK3WPraC0tKhrCfGCpGSzkD5PKANBwez9Tg+2sH/J73+jyYaCR1uA1Ov
b3TrN+wc1PnhI7ElLrZ3QgSnVLSg2u7Lnf8yja7UhO/zlwfQVEOgXzaEAk9d
gLZK8fwKPB5e9A9P5T++jDN+mDXUjW6dU7KRO8mYqbmtNiKOHi1YZRvBENcj
d04Ws1Chntbb3dtVu7xhbvVr0uqA8+sWKEekAENzkcnBtpiMbi64xnfybxct
q0XRcMezLyV+H1Cf412y2V62hZPlIf0rLJlKhJqD224bgAy01GyCKuf1Aaxb
b0WdGL1cEVR69dV0+jeevg7b1eF0yg/o4mdxlTJS+dBBXNFU8gIugBbZr5Wg
EfWrmUeudskG/tcaB1FOdFj8KDX7dXybWs17Azz8rxCv6DF1D1s/d28WTE+Y
WyQUiUmbfmMunn+8FphoPwTmnyDQZYZZ51GKjxHKlvYYhSNiM/70KcMp+wL2
YEnJkQKsqsEGuqEd5125sdDv+d4yB9V6jtX5LFJZe2fCazRIrTCj/W1O23nV
M+KP4iLT4wRxip0A9Mz1s01+oxrnoiQtaj+tXjYXVfqJ78Lyt2pr8+ffpNSD
IJWptbXAoSMgHetJRLadOE7Z/QdwfC4dfMtuD7Yitm8doihk9+9XO0UlcCFa
gazv9do1/QIUpym0xWu91ZaKZjBoFe1rI5AOC3sFo4vZ9t4B64HhZtSv8vHp
K6esBEIOQyVJ9+4qBO0dYYnQaI3kHC1j6QNrFO1pmYV+a1P5symxxhpTBS0J
leCzVReoyUbqC1IrUJ/XciU/CmmA4+ZwdFdTvZMc2SWuPoV9t9sWBwxZzR2R
IXSrJbjiXkTFFXCf/nmzZNVNipzcdG739mHjlvpJVAW4mpPcQyDqpGuvldQf
IPzOptf6E5buBBfbnK1QGSNV3pdInEYkDUR7OVjqN17/+EPBR2EAl9d3n6O/
APkLlU1QLkjPBmxX9PIeOSRO0Ms+5hvgdIfJ6CxDb/H9urWrh/27hcUrpjsN
Q+VFEh2kTFvhJ0dRzOebJ96nsevA1EniOOQ/z0QiYnf6K5aYsb4gbxA8Q8Y9
3lA7+ZnmbbgJWlpWo2w0bl1OX07puTx4jfmbWoPmrY5ZnG6wrVhVzKni+80t
XpaYqlpZo0u+3FElGceDDJaLLYGRjFgb8vrkiOMgqMPmZ8Tg2qPGCGIA87G4
y+ENlc7oLY1VhLWAuSy/Gk5SWKDZka4dAqJP/sCjiny4fMsyzC2sLCqQJ2gy
P4GEs4UiXEpbD4F+mN3c1kuv4wWoV1JNYEqYzO2QU1chLKxcfWF8ACes3rBy
hhFmaw9oAWTcAI/F0zrpy0oX7u4PHv2onmKJSc4j0Oz9ZjQPTNsrqdA3mujT
hcyZ6WHfHDNh0l2AAgMRTKlzyKbEUIkRMbIf6a4VQZd1iRDsyNLMLgFGlI4S
TnQ2dE3xNyXaKHDMIYJDgTPCHu4SO5pDCjYWp/+695tTtwO4seR4vSEGmpSz
rjbHF9M1Yv/f753tS7scRrBMOuiGKDVdFrGNe3Y4N6EoyBbuEXZN3ucnBnvW
AHw71lbpDHksU5yV3Lw/1Aah+eo/l/OJpUjF/K9djoVxgQ+vZDia4ITpVwVV
1/TPxhUo3U7/zXNdaizKEpsO7+5Gz0chVugIkMNpn9IvYiM3vutI/1Y2LvS6
mz7m57yyddlkP8yRiGP86b/POaLR35hbFBBHlxgXAfyu7IqqDq2aPIL0TRXO
jD7YKO8JnOI34E0tmMhP2WPU+ZbuUsFYq5UzqUgUqNWP/NxxdHMWrtKsYxf5
Vqa3yo53GBSrb0LDY0l29PIg7bJcdGFVa8vKNcd+TliR9Bp6laUAMoBxScDb
4RPaeTjtDj6NqFTLm1raeZgPRQ2BPRWvsMKUgEeCkxo6nOIzTGBiZ+0ENfNs
zqWmIbax4kwkjJHPUhUePPZASzLhxqVlLAeQ0AtyaTbVJte5V7fMreeQpG76
N1BiF3O6pqZaluZfeEoRVTNscv+McK6riWGnmuJd7hecy8+RCmssOhPi7nPa
XQU2/H3YvlCddqbbhaGVx2aOSG3RJjq8CLg8JiAf9fqCqN6gLA9YSykXxnEH
GgZdcSXVuM38IohAqnSHVh52RmELCkiNsiD9BTbn74+16thyep3zLrHDkFmp
Z9V1mysn2s9HdwQQhU2Z6x2TxzKN6cBWqnEfok6IWWkzRamurOr3bkzLF8r1
gyEcbPiPeo/uSupu/feD+FJXSsFer/05ciCREZAjWPFlGeumHoyeQToVc4Xm
AiNrzEdd1uO/Yd37hlxSdL4FF5yBMUI8V679lNoEIulKi6zsSEAN0tBOgo4a
pDdjgynTTge1+gBBRZaxZqULKWg8mTBvXDyP/ubHq8M3XkDKxvwzt9gv/8tC
jazU9KiLR/knG8LPxehARv7KxqBxOtH1WP2WtvNxie+te4szH6xzdPVx+jY0
xsFmscItBlROUn78GzXeftTp15v8nXR6lfgSiop/BCJ0++U5SOSwoXK3p6E1
sHWa/7W2QrBy9am4fKjnztmOL2b2FMQkwp3sH8lscDhPsSZ3BL3EpB246+98
Oti2F/UGJlFch3sUT6505Oay6x3pLKIzwyvL+qOwDN2KBmLAVMnOQuP65jOD
ZPub3Vzag4sPRqCj3kTNx5bfDib4b19xShmt8ww15NKoaciKVkEd5EcQWExD
2hPisalH+monybckRSPZeeHAkY5Ixt44WniTSoYdQgzG18i9OQlJP0HOYF+F
xterDD73iJ2Ptik3Y8kUC56O5rOopgwXHTr4yBm3AX4WWaL6TSZxfNaLj+W0
BdV58TyXLqzxtiuiSZNY7D21QMYPdCbbqHQNDRYS9JJul2qzApC88vB7RoI7
QkLI2C9hZVqLvwcMd0DbZodY62jSv4cmngGQMehTVmnL7aVkgTwzRDQQoPft
R2tt85l2T6qjRgYQvBgik5pHH5m6g255RyoPrl9nf7C6l+30piVVVJUqg0RR
jLACQsS31ZW2eRrD/B4SytpdpV9U+kQgDAeI2b2BAdfXvygn69MsbY1YNq/N
joFhGEGeiJQdfzFG2pLChmWj/E52Mucs0YdGSLCmARZc/Ee4mMvnLnwuBEm3
8IfeR3G376/e+I2NhtC0nNKEzmBrfYt5Cq5pLbaIeJCYrUeg5zqi7cqLyENq
GDEcC8c4RCMv6/yTX0TkEw1aIhbZzh1beXnQeZ5p/wrdkJfyEOSIZMkBnnkG
8yGZzCUBLtcnfIb/X1eIHibmAmBr1VbV0PD46jgQ/spE//vMcnoz5eMHC7pY
iYM7kXZFGpYRVHvONVHwXGEVtG6zsj5W6AATsYcfZNZnYYDPNHVM8OQCj+LV
0n7HGomE8nDC/O6V7IJP9xaTPlBdrY3KT7nbPzKkXfDAJhv12BSAC+DV+QO0
gDUC/lXKoORX5KTU9UjYJXZ9rlGik+zpyyn0QbHCtDLBw7evANj0WcFth5rm
ZdK30zZpfdIlyhIt8JXfXPj3hgGcqUhwUzIn2vjEoxSS+sWIjxukPAZ4CRrY
TQ5k72UWEmWcYzEWdg3NbgcJlcdY/kpk8Nbs6C9j0nQ5gZ5d+aCR6Vi5fdY9
6cAMz3gjeYFBxj5cZ8VZhDeeTahmAwICrTQIBNfhjD4+rwgDJ6IaosvLXWRr
fTBJ+3r6zLHpY1CKbxwnKJOUOyf7C9B/yab1hromG6r1rvt8r0GjaG9hRrS+
8KkQ+qJ6OrrRSUguFaxiArEZrLvb68zJaZU/UH7ll/n8QCoh7wE/WX5nvIef
t+XbcJtJqMR/oag+zxiCYbsjh7rwymMIuJmzUPnaY1dw7TuWH1f+kesIhmmw
4/tIbUr4kIY17VGOkknH7cnmLlGVgcV63MVzGyl5We5qDRKNoplcMXDhcYAS
cx5+o/WpzLq7zdmoejQDo6JIY+5SXVMMC4YuKyRgbj+4uotJfmVphQpFl7KL
6rGgiuiaQiAPbyDkUoMUZWgfdgZN8q/eoDd/W96tKl48GLBdeXFSYzQa1kf3
7fr6P9MbIZfADQm2XIWKh6uc3mlCd3twy8YPuvE0EcVP3gWGJM1+b+enlKha
kPyRQSXKsX6FecvCxcUT/92r6x33GWMrWQWNyPqGgbi5yJCfXmmD3BFG7q9w
rqy8BCc/svD95IFax2w0LPVmbIKYdko3W5K7iEpJmTn1zd+Z20Q2T8xyJ0QO
SrxHQMZbl7DGBCHeV27022dZr/ZhEDgycUM3ju7lIRAW8aiMUrNsxvwrrt2B
eyC5JsReYdyWQf5tbqPq57GiwMeaOzHdi1UnI5ytVuRjgdiApUfsuJ/SUOtY
Zkdt8IBxCab0AwyWIe8rqwLNf3emaIskfdk9lA9A4M5y14WfsmIUkozFCNwR
Cv4fz+GspDV1PWwzj7Mc2BCtpyi7F3JYUmuuik1vg2qCfXoA5yOXPD1ByGAD
565o9ZW/2wLnt5Mi5eTkxKz/cdPdseCVLH0ZtAOcKEXDHgcuDQYzCN9wOuko
8tt9rWqio12Ci+OdXH6uc9fDK4jq0hmZn0k6m555vC2b7UcCT3GMsGoTScUy
8viDNB1k1/7Gy54Z8eiJHyXlllnlHoEDaufa8J40KD+wXXJ5F0QEksXmWPTI
61laxxN+ybOziLcrCsodUo2t13Vj2vvt2g1o6G4DOinTNJ424gL3sIK4kQyP
a7MJSBE7J+TJfqngOtGkTmwQSL4T/Dps6jBt4kPKCqZESIPuy+REFMsC+mFm
N/jDYYFfqzq1wh1nCF6goI8+im4EE5j1K0uo42TqDlSRzXRkF0HNn+3a15Ob
xghmBJoK4Ltxaw+6ZhZX8N26X94i6Wyw9e/zMKlG9bprmCZXijUpl7512UCb
y7rNFLLceyk2Ye9zJDXBdU85vUGN544zgVSJR/lf9bghdBbC42uciygoKrFP
eIm0lkD82yLFrQlYQZ9BKagMNoiX1b+Qal2v0NBhp8rQptvISh4fNWNqMf1O
kv5x/6gKiC1pV4sjxENZ8KrycLIGTE0Bwn5XeR0EeCxQWvtAxIei0Kp3eg08
rSLAyKFpkyU5OnFFlTrTkcsBXmfMke9xVsOuWrbokjFJt2tQqY7LJ3kJyG1t
/sTWw5ainIFDSy1RHt++bEu4KCEhfWbxZ9nBvbxtK6dQsmoODkVOMA04kq/C
MWFeCrSKdtJ7J3LqcnJP5Ya/aE1nJ8V4Bf1s8GVfwBqs6/kucVCklala7HSQ
STnp1xpFrgHpoKePDqKJNH4Ji8grumdmHeOqUZ5l1GNK211iOLiYLy2WB8dU
ImyhEtQpy63hVuwWUHdVIQPGxTATO6LG98S2oQSYDakyP/D0RUkfvfcsZrs6
OX61BXVW4os67B11Upa0aAD2sCGdAzpDOkKyfo8iRuXJgpG3PUR9rqEsrNip
18LUxhUVjeN+GnpVHDk9x+nNCG3ZZvFLXQh1FGR8JvMpqbneqKlnEckBg3Kw
nptXi02HODoDolMCP3c6eHqoipv1eonUK15q3urE5otj22PXxRnVaiKDRKSz
Xwk0Y7vMUr3r1vFs9WDxiSVquYcO+2C4lI+jJcWkWExwiGPFOYlgDMTJma+K
5bXLiTqE8Eizrp5QXobnHGGYZFpTsN+b+oPJUL/0AzK7JFxTNUxh9duvBwUj
jbllmXvbeismf5v89i26XyqDr0EeFzNRagZRzd3JfDNj+TJ0tqXTtsgirgE5
WzDdKUUXCGKR1lPcRkw9jZNxjTukyHljids46ZxPIdToA/xLrf7LkPNrPDHB
6pUsTT4A+30++hcDcuw4Ppw2SVbtLn5t6ak/UUG8YeRXdoPpEC9FlFS/PnjP
p1cj88nkExXz9sjDdz5Fqc9WQM/GzMc6x06qpwmyUgsKcmxxiEFR4Am2fS92
s4vAQsu5D35BEhOVQuaGTv24TLHVRnt4uons1B5MCm35xtCTleQxzWL2NGSY
AkZwxjG/Tfm4T23OBM87YX5cOCA4RB61zYpdIpPBl1y1A8MgGPf0ilQ3qCHW
SqncVkuB8rsM91DXPXcaAbcuufUMXzn4rAVjUn5laeeDGRxmPpyLRTr5Lx1q
btWQXlGxKwvKrltVeYT8/2km7EqJKjKr/FA6vzL0cYrDuDu8AmcIAFKJh6yM
4rXQ4+CW3l7+p0LO/8oQ+mqsYTRXmVv1+lQ7s9nOWFX+oGICFkmz1lnA/YZA
JLRPckAMbHShvv7tGsVThmjMuUcDldhnXR+r+GfrY8coUdXkIU+7QmwonK3l
jXpBUitDvdwNOYMBXf2CUaolJDMPD7gEh2j60uMwbpzmETOyZi2NstZlCyxs
Mycv4fpPmkVFTQWx0DuCLuUu/Px7ddt7/NGZ1n8bET4qA+XHXPvCCtI386uY
1/Qvvl8tC/U+tqqCq5nGHLc/pJP4xJtjVd9LjrJagsEBUrAkn8MlWmq3CXWm
9IJzR2XjyXjfpDVvP7PYDTN4uwNtFkGDb9gBpIBSJkgAtz5y/W4MscqjM3zG
1V5HWkMGydVMA8vWXDZEDJdCXqHtlZt9OUOVfBLp3hkMah06StDICK14emvu
MGR6/71LuBMvCe9kzN7xkWduuXVUQPlAJH3Sa8Tzfy5wt/AGh5xbBSE1aM0Y
u035lnhe8ZcIHg3DCV7/1jTMILOOFf5aPyS7YCxWsZlpZlmM37rTcl4y6SR/
VZriZaJ8i0BEtqYr2rjJCVu4yQZcZiVewjtx6wTaz2pbp0tTXyQGAPplBaTz
KlY2E2Obb1ql6Etyb5vVgV+omgIrYUfPjMq1qa8+HJ36a4tinPNJQoTT2K1h
c/KVDgtrRMhJjyc6vMbcp6xsSU07hlet4d31H7D9z1BMpzCd7EEP3VkozuLD
TCopagseLDBwDcPSPpoSqOa9o6FBzKw/FXcaC8ZMbRP6MxU4bXPJ9ctTZw+8
tEwxI7yjYgVZPufT+jPKVCHWW/2Qb5erILiX5Iz1VmdXgP4AZBsd7TTaguFS
WPU87wWsSNlP44zkQug+WamaziVL9H5hVZfMVFVsOSqoiEuebhMu/PtVltDH
t2DMt4Co6e7CJpUAwn0uxkAkJaL3iQpLPGNVUKIrhzseL3cFALnPZ9YZJCYT
H3bE5NjWZ17w8lyazIYvZ6U3QRsXwP1nR2nbwxV8PgDNjlUME4B1FCXOR50e
g81UXdKC7l0F0BtZRYmpUGCTiYmpyJ5S/eBqPBd2+ywyJx04za6+j4eBu+ez
s1IdmJjGiUaVvRH72+QfLggrmUGSoqgKEXR0AmBxA5mvsrgj8QvXp76w+GE7
odZ2EBhXRWz/LO+u813v0+zyOi9RQMA0joTvWJzdkJmEGlQ27e2fMI4l4Ucy
2pP/ZKz71eEGf7BUGJOZdtUUkhfOFiENboIq8tHHfQD+C7I+9ugHnXTjKCfc
FdLREJih6BPPXLONLxs8AKLmb+Oj2/3PCcZ+O4FssSOoYu1RfMhjhifWHimt
GueqLvw4XJlu+zMXDjRDp8o3vZXu1W6X8nYdeIk93uEddEolKhDbccvx/a1X
6yt4shLLXodIA6Nwc2xEkberee5lD5G/+Uh80nWo7FtWe09vh1aTVukPl9Bm
10D9XCjwTSFLJWDZ5+TG7fXUjkjCVY5Oa7NfJQbdjSeBwiB0+Y9DvrTzdoZb
VoCKSDemmZLvtQIvvKkc2qyuYw0vIzGbN6sPzWTQ7RKadPkzK/0uGOMEDGvy
cp2yp6IUnp17pegdk5+bsET+0m4Dyiww1j3DlyVPCKF4G67nud8Y4jvqpS0b
7yN+SUVId/nQfEZ9BUEiTm4DrlKbF2Bgwt4QdeVzxpuzJbU9JDzgSv3u2v2c
6NxBnRR05Em5RlNBRwHXlQdM1tVMXY7poliuJeDXRjY2Bn1dpYO9m7CbW1oi
TFB3munKS64cDqKQVmQyQ5Lyyjpy1AVQwTNNFGencMnHY8qyqcqF5GCwo+6Q
Kn/stbFrLKrkySBKJIPXVXLxX7Fu34X7BcyA+wv7FfiW+e0Aray3Za/frdyv
m1gehJpfS4q42Z/NHLhinWPK6KiYyVmzPMfyO7XBbLC13U1F2amBDrsjQ04o
mUz3CwPdCAxJ9HagO/CWfgSBvMr0o4aFfGRzI8Pf5MzN8WcLi0Gym28pwlKw
kU9ID0sEfz9sB17b9iFd4D1yEl1WtMd6OS2Jew4k4Ma5s23hIBi6qWeyEB2j
r+Nbxu2buYNJ/qIQKS+4FffUcC4i84qbFB8ViD8EeugW0UhV2scJN27AablM
NqweQpFilqCSGScmMKPWr1C1EW7zOITljo5BJXHzMcEDaoCB0j+uveXgmMha
uWe4295ps2eGQuJJwzTwjGaK4ODhqW0glJwfVIy1BPdUbVMiNTZgG3mBy4FB
GY/uwfQS4ERuUHiBBkKJ/ZxkJaWU/BeuHKgKKqGCRdAn16VE5pEky7x8P1ot
5jy2cf3Jst0zXc5dUqD9QE4fpIUkDe1EFn50TBHWZuMHP8Mpyhe6RErZgH+L
0R8heYorUUdB1Qx7cDCnuvC/Lhn7g1yRDNvVvUFJXHSJAiqVoxtKNipxMMx8
C8SeHvyspZSPohX1DIihrKMIAleI0QnVMQxaMJFQDTFrYUnWLqX5EMIfGco/
/zAvYhKybXZ+79GxMQy7zXP3Nc4fSBfU6nqQgfavX66v/jLOiUPnw4n9EyHx
YVC+R0ZUtA6Bsbgj+HIgbC6j4FLbvgeh1pH77OHyFhvQTsrJ7HcOIWxZsgb3
8EEewvp0hYCXub5VocOlX9HkDxcTn7doHwkBxGqIkJXEAFKnW9r8G0xXRBx7
q+Ftu8Fat/Rd4VaXKnE+CjFwk3wrRUvpADkoHvetG8PUjoILqoN/gUmg7f3D
No+bXFOUATIwJM+nTY56avcM5kc9Tm+8C7bSsGVAfOr8ECQQuoTc5E4aIEMZ
0oBgIOsDUDi/nR0Ytgnwc+W/0KKdEpqIJ/IlxxeJQBpl/RU7lGqlJh+gHYCb
nCJu7ZdAZYuqS1RmRA2SBjMo6Dyl1WChCXzCYHBI5U2l/Bh4M+HPzrryAz0U
sHtf0Nn28lHugqDzQtWduGuIbZfPRxnOWGqv/Zdn5EZbMr734Jxacu+VRUW2
bSEt0royCNCcj18ZYMxgn/xq/XqnqudBysus99pGFGdkcO6C1P4erMVSwsaY
St41hEGdvblE400vbgfhKqpoW7s6doxI8GAmdNFdos4kGuhJv8cdJ4xu1Pdu
+qwL9TnoYGRi844DntWBaaaqqObT5yfrUBzj1AXGxyaU4h58qd8mTbHp4SKK
Wgh+0qKdqWyt0fsJew1fZOomDcMc9erYzqaWqX/BKsyTbzb0wXOwe3N1pC0S
+deJpfCclV4FnU+LJJM2HX5LVLAxZNi5Mw+bwJo1L+7kyYk3mYAoczRrGzWP
YliX3/kO8/zYcOdx6KfVqpAIKXlKIqbG1Ilivdjp5xz1ZxqjH9J3lDiuRh/E
XluJ0ZtxRdctS1kabagfjj53lJ7uElpiRr/54SFE4Xp5P+DZZgfPZZv3kYL5
j2olx0ukae5neiv9gm+w41WYrMhycX41Pf5JmgL63KxTC3WogP50n63Fg/DG
atMKIJvrLwbCumyC7YVyjaqIQw+4Huq4id9v6WEK8bgkE8Z/RTp+PoCQ+7rU
zBSQLex3c++gykSInjWobKorQhiUC+V7fnOYdnffcfgV4Y3sXQ5NBzSXvq/a
/nC34689NBM8G41ksLiK7AETnGSDrdqcVZUjfsJBR817yHlqCU+ZKIoKLGp0
GlbvtZaTxhAu9QhgctPaLKDWK0lDFgCszBpmH3R3FAVKzL1AAtCXnkINtLLG
oYkA0YzlmzyQ/6D3PhqYmhaVvG9z00D7fRtYoMmVsPQNcrR88OeCdLlZIUkS
Js84b4Qljen43i6IsXKr881h5FaEitDsRcrziEJSqSDt4LeR3HUMv3zIy1VZ
T7ExBCG9lgJobA+eRU6sAnEOzsD4YAMywffzMlOD+6m91Op1xj70ENtIfiY4
b76K6JhWwJfUtbVA3OGwWi6x0GWfKynm/BUwjfShjvVeljEUjo2seubODivz
8BDFT/c6CzeoDp7uBaXHLQpYLHiGWin61IbEO3sDVGZdUPj8fPm44jZW4gkX
WAbVXJhAEGHI1qmDPsBDVyh9G9q0i1LgdqYamOqAvF3SQoTOyR+ZBZ5W4g5j
utWmY/p/D37B/CmJCYI2mIggHCkkU5elNySrma8HJbTOsZLErUEzKwBRgxxX
bPDSrKYAhKX0F9ztxjvBis91P9+pDe8exJfmaDujKjnCjnCmXHMlYhLodAl+
SG4n17Mr7wNImAVSIjurgHZAs5HUxr8c9RvmKQTJSuXznAQOQ5hPU99Jbm2R
eWMSKsGouZkll/P54YMMjj+5ibMRPSRvOLOFyoHzHFm7RObQoMwem2QeNdZn
5Pte/6wK/Xa0gXv4iGYpilg+zyIG83RXxR/GHX/MvbluKOtqZKfIki1MDVFj
2uOFMYsFKqfQMy4MMIcME/8JKWbsMScYy0s4bG4AcsZHJZSxx4Wzz3blblaY
eVEhtmT0BZs6HsNUqxzET69jxuxr3Jo8jZTrtZLFLs8rrvSKdxOe2XTh9EWr
O3ZGbLrJtlvX5b9R0rs7vAjU5a4DbvccKNiRBnKBWuz3pFvRtzpiZngkLIYa
/UxZqPGC1oHD+PlVLk+cuAXxFw4u0nRu88KqgRzb8ZVduBBM5SNw4QVhXKJg
ihexmS5glWwgVUbBjF7Pqk59FL60VCuu+znpN53qYJ5jL9GXA6WDc2h7fWAH
6pZWFfHKKHG0eCFT+5eEnDeEybTnu0M3QDb4vVxXr8hKc6oqKX9kgyq6FN42
DatcNsymYXweJTwgIG2nW6RMOCxCXfxa5gQwOALr45AIP1vM2lwK4yiHkVI2
JM/qvY/cc6gfmQvfs4Ji2ur4XGiFbSe4NImsr8JgWJmlDEa6mQtrentQU5fs
loV2ZUMzkIhXFQb/nz6d3kCKU/y8vRGXzfDwzQDG6CmU1hMwWFCLCSTT0s2v
y+BXKGFiopZDOSujTUZQYzreWs4Ml4155Ha2EHlIJ6ulfoiGuQefF7owD7Ab
oaNlt1caQLR7wamlOb7lA5AlI5WJ9o6BNd1oiTfrjwg8NOmg5YjadJsJbmuc
A8QumB10ezTZCRPpqemEHiaYwzpAVYDVqDB8J+Knx2Oy5YF+xOl7kW2NUcIt
KqgwusuIRraLUGDud9xPXvTRNfFCS9A+qP86xqs7mVUx5AVCokAUPHBbThkF
meRBP2pZlwBWA4BBm26ji68s7NL7zHvGFtH6idS32+R2syhBzDJwVAorytyF
+DaCUx1guuJVSXwviOPBCEjgpiqcXQj5GKU0qLq0rRjSvLtzMxx6wCnO5J14
wHQ/Y8OCc6xqZKAFZkDF/ynwedfR/csyBzIhUjf9B0oF3gLdJ/8N9ywYgOlS
ulPPToexvjUH8AMhrcmLxTqzvnLAv76+Dw0s0bqVhWF7fKMdntHQhLAyn13e
+BIXK4xsBW1tux2B2ey26EptCr5Mj4iIh6/0tEjPNqEQt17o3zCFUMIT2pXm
Cqar0awFLTddn2c1RxVBgqYnznfHNHd57riB6126LyDNnuCI6etmYOyjkauk
44mJDn335mLdNeD/IzhxYoSGiHMCX2M5X0HXu1tdRFegw82alMTmKuDodlRq
SDrzR5UbQ1aepMObrGyJWSn8iCrpTY728zWHlr1MrHZRdNIKDXpbm8NSWUZz
slA0chbpUi6ETrpYrBQxx8nDaid626NnRGfcHTLvuyO22T5OLtGbEqLmfEJ4
1lKRHqMY+j0Z7IaMPWgdItdeR0R8Com7hsfJR7GbXMGOIDplOXLYBnu/ov+i
zcaLm88XmQSR4VCU+2Hx/GH1HaLlPrAVwIWDYQy8xjh7WqYZfhNstSz0BzQo
hLNWXw+L2Ul0OIgWdw9dTshU2O0ULdXxXy16j0OO9NkdIYu/MIpLCLdONPsk
TnfBKhimQuJz6vLDtZ384uwBehPRDl8phW808z+zT6fROtcpx22MgiQVyf0s
NcLM7x6i4ypo+cwW7fJ44t51hoFeXrhiGTQOfe+1CpOIuTWDuxz6sbwTknpa
/gdo0sYVln6RBfoJhd6GGDlItIycUXEKMZvPg5IvFrCXsMUXL0vnvIVCbjUg
doCUu3R7nzundbGpHAEU9RIZjEDBH+X3OqrRMK/Ht8h8YpYgYl4WvM06/HcS
DXov7zs7ERm0O+MeVYhRrkLG4C9tcrTE9nblCuaDPb+E4qdiG2/57Gaj6TTB
Q4YF3l2610oIVpBH8Op7ltQ30sipuOBQgcfNE0hnU09TIrrJVmdIH4XVxv7/
Dq/mOiH+LMkniXP5XC6v7mIFXGnzr2UKIYODHjROgOvaz+fUA1uBmyy07oSD
To2bRvqCwvYoZKdE25pifdX/fFHHUCnm1tQCOx2WAMtEfCKPz4/cv1bTc7iS
k8PU8jULZ/mBXlTcY7VTN5xbz3wYD5Z1A6EB3cAa72zDDu0sZ4d0DQC/6cEq
8r3bKHF8B4EM9GbeVeYg6ZkCHGsstcxB3TpXnZTvdFl0Q8h6XNCFSA7EIsp/
QexKffWfSl/AF/of+F2VqAc7K5iyHOzODIcdWnah2eyKm3Jx5T5u6P67v81d
CpdUYZIqSczL2mwuvZBbnEwzSsBIV0hreUIVAlj28434v3g87qwnWGij7oHj
h5NUQB2tbXbVxgZiowXiZ1TlSCXtd3IfrarFrvc1imSkmPkjHFXuwT2dqAx5
1c2USut6F1GT6UeDlWafmTmHV9DzIjI6Uj/ed36lZy7I1g8j7vocObewm17e
4LJc7VM0j/ydPn7Oz/coUb6iIqti8WGR/8oskYbwMNtKTctWq0fdc0pktilW
g98Yaz0A0jRaT/g3ei9PV/Hl6pDSC5o3KKN/+ZMy53OYCmP4l2z+IFNP/rvh
DqL0wTW1PxEGIaYr2KTirMs7Rkkbnzv5xR9K49SPK674LxQnEgOCIb2HOhbu
KpxA7camS1r8sFCeClBqUZCgV98/LDaBPEnzjNDSs0XkWDqguGGYC680G8Er
lcuMe6wmlVH0ZFwE8N4QnVwkQLGQuO2o1mr+jwIULJZLfHScFFfgpf00mnB7
9eatHtzSSmbOHPARk2am3U9cf4eSHz+1ew2ZI1mtJskvB3pDv3U8p1CJcBwn
5/9WVve2h7p9Yd71ih/yto2Nu+NadfE8bikeRxD5/mg0oI0tjhhR+kSCNpDj
SQukd9pTYvVnY9K2oAU35GN+m/nb5R8AIadBg4si6GWhS2Wu6oY2yTmcghHG
hWF2F+tB1EZpyXT3NwfRzsEXnT224tJuN0qnKeNQiqWzemW0bB+IVtF6wAfV
1qeA37cCbAxJyeQYjFEXNybLFBhq2tbUk1O82Pg0k3zEV2Y7W4mmCZ662UFV
H25wRZuo5BiU9Hnn2KN9fSu4IAUuOqt+tCOaa0rzhSwc/gSFNuZUnf2sa5uG
lA8Wnm9qYtJrlSGtrAxfU61O3RnXursh90Kp/RLfZuc03uXjnfiKutdKhakC
4rfvruQipDk+5CR8pX15AYuVWHiEJIXWAmHUMTOpjNWVY2NFA01pd4XQtefs
dj/HQYvupvBL8HhasplLcoTWaAi3LadlG00V6KsOEtTm7KpEdTvy3ArnrjMl
rv54unmtmdPp2ffGWrws5h1kZjyMm9I9Jw445tk2B857D9FipN5rZGhFhba6
9z3VClgyeoNhFxQqq7VNcMlbUfl7fc6pFvXixYhCbLMpUtYAL7TzlaJOT0CI
z1mTODUBVTZPBDSXDGCM5wxE7mMswJizd0KRmPJ4e0il+UuuxWJddogog3Wf
UIroh8Vg/L4lCh/m2c4a8us4RJzF/J8r53knSmtaml6TQuT3VU08fv8tdvJy
yuxNyKZPy3qwALer18hrL97EQq0KsS/ozoW7ZaQwF/UMSUrcGtXWL0bRprkR
r+zATi7BDfX+gm4p2I07rG/ULXivcf+y/w1RBUjJzDAFt9tqtuPu/X/sxthI
py7IjqG8jxY3mJCqtla+XMXrdL2eYCcUcBoIURar/2rg7jjc11e8QK1lpuBi
cbACH3yvQzxE0OIDSUOVucDv4P0b13uqe1S3/5sv47wJogDap7snTiuo4ZuH
br/uThBdLidRQbrg6gP/EruvaZ4/gfIifViPYFO8hYIhptddDqNm1ylxU4+f
6ZxNO19JK3MIU5jsc08pn5P4R43gvUTLaSVZSgVwBaVe9bYcWBgQuBDSc3+g
UPbdcZJ1/6+E95blvb+AeRfRqSgct84yVyYzUi/z9Uhftz622kKVNGNRETb8
tBjn7hjIE+7fmxHTb6vhpMetR8J8GTgNuReGN1DSjYl+PQfym+xLTchheQAD
a8fST/cZxBpopYI4GrMkLL4vse0kK1uDOftHe/StphtQ0iS+I2sNuUfW8CgQ
qXrEmx4bGG4XLkHok3gHa36I9iCX2Kw4xpLTZo3sKSsRENhJxHEL0kPH7mK7
QgHTw7OjMT9V446xCgokN5Tydpxt/EPNsXt+kXZavP/QBFTB3ZbK0w5Kr4Ga
xjODQMWPmS/+qYgeeewuoHu2cWlFIPllD5Wh5Rgw1kIj/w6avm/k2mcbuk7M
y9LCM3EgcUg/dmJ4mbAn+GQGOL09g2cL6ab9esd1FEH4KuJp6OIJpQzzd+6W
r2e4R5i/Upfsm9h1A8oGY2BqOrsy3yXi2uLruOaZgeZnENw45JaCC3+ZHlWf
4JQnFgKGR0Pv+eG+K+rbOXV4AyOeNUyf0GfvZ/hMX7k5TOP9ckJVvxQhiocn
3HBZqvBxtOkgGpC56XqQQ/WdbHiOdRNInLjQOgGlBZgYhBp2ILwHfhzKVGT6
A8NimuWiyeplPtO0w7CAIxmzT8dto3DF4Zk26mhZ2IgAwAty9MsToQiqGQnD
9YcEC3Bx8I0bm5FhUCyLnbwQIl4B7lLGxe3TSuaKsWbGC1xERRcamMEW6TR8
ErUubFj5h3k/kih9bMD0h6rbOMxt4vak2QejG54VzyMxckg7YeB42x89kAhD
4Cx1pdJM/pA6jUoIDJsNDh3MCrTYifLnkxy9D/9VRO2h9fNd50uPI1L8H2+8
xfOA9Ve0NJm6rQBRWVHgQnNxnN5fRz0GWBA0UdfLwogRY6dskHWTxevQmjRm
KSeTRGjbdaWQicMHWlwZfdKKLrcPgAe74JlhpWlSmAMZQPgD8R0bkN2SyK4D
kn8a6bVwDInlGl9VF70m9WviQSifxs7OnluJ9WsgMfFZaDRquDMNV8GFTdzy
94MeazwBK/1CrAGpV/CO96TK1XT+Ebo0NPPh0n3SQe4mJkUdPcFHM9LrBmKQ
EbUILlk81jRSC7XlpN1QynK8wJU3fSpyhkmn2OUGw3kFUYze1Icb/1OWiql/
BD1KRCOAFcVmsReSOQ5D6svIBNMIIt0treueFROp+IFK5o1lI3xEo5LujVNn
JvwCoktXc7ymGMc5UbLf7ftyKMQ9Y53qImeF7lFK9ibHiIpXKUuWTE99cM+p
iiJ/QtueDU1nW42kLRni1hpZ1bWLqLRtuloYLjFF9PikjHIsIkdk4BEB1Gi4
UDCNZk16XuKVYAXz6hdAt/6dX2/d3Mg+JccrRsDenEdJa/HVVQ6e3NHt/us6
z2Iwiej4BSXedT0v7URAi7fGxfipaiyLXOIGuTuR1aOaOpcyp8ntXkUVRzFF
Y1Xz0JzNEyTuCLW9qrTK/TQ+dfFDYVoo5Lidy4C0vWZ84ffmLXb00Kuofd0p
lDX21S1frPnUYihDaSDWIftouyDFD7qap3Oiw9bsegm2zwStqdz4or5f2sjW
ghUiLdMdNbZcGAZx89zadxrhd+/l+1cFaOqb7X6wm7BVv3MuSWc4dyq3DyT0
s+2sNT3l4bBGSvHVVpjV+hk9Y6bkgl2yQiQE9vxkQzdWJCjZdPuMIlFskKkD
PAPw9fn6h21n+SrKPOHOL1UF8F2Xbhf0U2O7tyQKaEDCZp28PHIXQ1JNN9tK
ZWuLsIFMxINFSu9iuz7opOfbeVuHSTxqHDLgLWn+HxzaZ4vnujN+VNC4IE9V
b+KuMvlrXDKApktOBeKzAagt/F4Xq2r+A6JNiRia2wi559lJE4gFGM3XWoYr
eWbQAqF+b6lqyuTL0vCVEDDMoU7QWpVLSUAYjdyUTnREUbxlSxxpHPi9mh2N
Xe87SzexIUbZQn3FFHySlKrWva6c21Yjc+d9Kg9jSWAGtdflXJEmcqVnSn9w
UQFt0A7s/IKrqv2OFqOnJfmLG2m/MFqvjdymNmd+LPQEnKuFdqPBd+71vlR7
NZOAfUqdvVN83+n/VfpLY0v0g+xixOFgKhg5OuCTECqKkLWx1pZDZhrQNonh
H3uASZQ6BI6GBVBmIvihV+x2vPmKrBO5lgZWi3Cp8zNdExnN2E7vMpyEItth
29pMhnECiTljOkAw/iWxrTh32+9HeHv0j59v0lodZ3o7y9ZS+i+vhMmpzip3
hVykpjjwfwJmIgKQqjZxtK6MjPCb1Jwfg6J9gscizvtZebGSJM3cHvFPiUr1
zOaDBZdQwIyXCKsBBydxivXSlvw2jt00IbCizXBi8Z2cJgbb4BZTmM8TFwe5
yzXK8ZOYek8NV4mxbPflEbrypeRraOrTJ8kexrDBhOx8EkocokTLPzt6TQoP
QDXX2QuDJ1FZxiTbmChmAi0aXYIpmxGFbuLZyJ94qzyOKXbFOehG+dsAerzx
8Udxo/zSBFj9eEiRyqqPCDdkhQS01cMlAAlM7xUJvfFztI/Viy7ty5bE86kn
vjOOnIT893Jk4PubBkRjNJgl4vNWU7333HKgCtdjenhAkHBDDwxTXad0QwDy
G4JQzTRUpjMKPL6OKZmpqR9vbJRSDxDHjmUi+UX6wZSi0WhFLmxFIOIcPBt4
NediYUwm3WC+kXCEmVi2lUWBT8RFdZ5rZ3tDhonCkNG2SuMvhqSpnvgl3ewG
FTLjUwhklk00xgT83aqY/1AJ45GxVv/rNEcauiGaUeONV/zZT7mL7UYULDn6
HOVGSDZefETK5+FESJudbbSBUDAj6lMPUytLwpHHNTSq7sT1KhR2H+3qdkpj
EvEJ2hUos/DYBItlUZ+b4HtBjpilQUaFzx7EWAlf7eY6jUxZM8nIoos/Eyoq
1AQhWOPbQ2o02NWWA/mVrcFVJn/4VxZ1ncO3vR+EAy/NLsfZKQgGpti8OCmZ
LovaDIYOdeTV7eH1G3ZnnhJy8orHHfeIf0kM6AQxUftoFGp3cseO5BBsxFzl
OlP7SYkyeWDVLIhQHV3cWHT6/dAQX3eu/CMBLazJx4EedtTjQcoXOVoGARUh
3c0Sb1v2OnEVVsQLFAzr84Wmd70xSFTj2gE4YhEMFPZWb1XO4RwpxgivGM+E
PbDSqesY+oYhd7XnwyCQVEqh10beYLlH0aqoDT6uGgTeeIFxZEejRIq67u4t
M0jG74OrSbZ/pKQM1TSwfxw0HcK09Zeid2x+hMRgd2qqNX30DN7kGs0QKVRF
xOWtzJShracv8MqvEPzZXsGZjX9T/2fNZazcMUJ7PELK/VqK8ehQSoem3Nhl
cevI78PyP2+SS4ebudz3jdDKo88lKAqszSOW5fOIlGcVrOa5FhtuB+wi2X9m
S6r58WrRUoThX8brU3HzvKG8gDXUmE7/494z2XmyaywXlaUTpKj20ALSDOOp
kV9H1PiVKyl2m6NHw5Ss0ivKcOwoIt3+H8PWK3psGhPBtEwVk9jKJOJh7pIS
PfunW/Rz/M2D6+y/z4aulbkzGpq+3ldFWw3ewRxwQ9Bv28pT1iEJWAlQHE1l
5OPc5Ep8QCnWsTH3YZw6szdmvtaWsJhw86tAU1fY1TxhETUFiG1j135/B4cD
iwmKstjgsLuZK2zu2VZxImCp7qbBHGJomA3Ds3At847ZaD3PhMHmXi2JY6Tr
/Wk+fK9X7MKPwKIVDSsQHoufDb+Ki9rqQqyX5sD4qAMVvJV4DS+bCcrAZukE
lYkFKzr8l2QSCIe++FHzqt6E3o9Co/INUwAp6RidIgNj6zJtFlFQuAMdKm/A
GV2goaQB8mpYL8kCMjEAxN0Ww7GlcE1niGynnWwg8Qv2Xlc4PARU4uOoK1di
X/61BPgfZnzDWlyZVW0qNuiY6pTTinlWb7XZLBGvYPS6M/T+iXQAGdHPBFk5
Hm1g3WCC2gvHMVfK7PGMMzG6GU7oNvsjE5D7x/D/W8YaUDykKLvQ98o4TSSs
pjITD3Rq1MRbhvlnvWb8JxqOxkw/6BSfgb+yvwR+PYMKeP2JWexquFT6XT8G
augpDItAb7CunPgUkr6/F1ERWz1+9HQkybtaylypoFa3mOZ3Yza9BZSdM7tG
4GeAldSa8XR1bxHPB9PTsy2arWm/viO7dLT41TwKmiRuru/bdUXDlycaOV1k
O7havxnMx1fcVR/z7MLV4WxqxDMxLVYRUmQbWtqc9DNJ5m69zgHl8bL4QTFJ
a36+65yN8nd/YSb0twN1mUkPDOe7WxlHV9BhA32XT4GlRvn72qrX5ZEYtA2k
8LqexF3Xm8qvtXkWcifXv7RniNYh3LKXkf8cpjtfVftqlcDOiLgbKm0uE1Sb
Bas/AkuAaASfDItmAkm8QgD3a9GEeykIiKJWzF+G0Wr+GWVhIkkSGZwt8FEs
qvN1NObwuIcKZjjxTlLyaJ0fGQwBeysxIczDNjR0wWFnFxu0CZz+tSkOf3oa
1gb12n14i9RJIs5uWqSzp8X4P9u6oo12ncDnZPEZ73hBiCDMcnXc0qH6IsuZ
MlpPABc91G9pvv0IXS97IYK4Sd7hH8EajJUdD9//UyrZOEKhgY9/jm1kpAJa
8z2VQjMQMIChvtLEvFAMIW/nfDPrF0l8+2G3jlDK6UYJ/zg8htNM+aQaMQDw
QeKgx22SpBIwE2DJDlWaaXlPpRqZUrPKW3j2wFjeo5x7HkkfZHdtVbzJfGkK
2spa2lDjp+Y+tiBD8TvC+PXmYWiqD1RiS1Y61r6R39Aj+4ruPlae9f+O8RcI
BPzLqXYFuUdP4SEwjvxgEzYvH/vVmmfuqOikAtZX1ve3Zr0NzAvH3a/FLb1i
ocyfI1B+V+JksEeZmxlON2e4icxMucEPbEtBlF0G2nyjDqa+rBacfP0Qb1cl
c1o4y/YABTF1DqcG/6DxzDWG2/rgpOLLHiEDk3R63FpKw+Tov2cIu2UGhzob
IYc35tIRz4ayONc725teBN2W2rQRnB3AmbCPwHLOjo+J25/8CikqG9UnTyq/
fxGBadtQCl3OQky3tfDdvCJhhdOc6auB0z06R9lYwSk53t+BiKk/xhgksGkb
YIOjRx0UgLIFbGf8PXulXXzbP9/cUgMZSSA5wgM7zRDG0+yhVLgzAdN+QE5s
rMW3vSUxoKAnZ0lfyck78ot40GZEhYa94YrbPMpcbL+7Uly2i1vR3o5LelSM
hdtDsrX6Q/TJolCjl+QsMUrhaAUzOd790RKVa3flUU4Dfii5q47EbjNc2JAV
vtTge4fnglww2xRBTEqPJmj3khHglxVrV1rN7PHCibyY4JS1pVtLwZQIfqWf
V8UDI4WmXFIRbNvro1g3RMJKh8cxKHfHoULAvDuIWeB4T1Czo8OqRF0zwjeV
jU8nRT/0oPPREQbQZl8vAeAmjqIZ0KIfX5MRK9lW/yXz0CPsrYLD8jOYgE9i
fzRyHG9uH3pE+UthfP/ElcJlreMBvuKmVehyogn7XRukebyJWv4LkvCL+sYV
gq08SVnWP3/HjvmUZnH4tSMrrF7QHZjBAni0liEjjpZKiRefaO2iMt9Xf0GE
k6VsFKOtzzWUKTh3WnUEViLTcxOLxKlqgy5VpWw1LYGRbxPchzGvTzx8nJrt
5iSnDWaVVxOSLdI6T6fBvLBs7C4QqLHMdipDpW2xPiovJpKbKnl+eFCAgt1k
YiX3uqhHqysZWKvINUzXXeloFeDxPyYYnFNwDbcH6myswacFw9sMowubwk5q
a9Y7e+ThrjakaqftKEnm8vqXpE0orQ0aL/qjnK2LfFvVzANf1CJjlCs5sUbH
xg1DmCtVuedZ6s+vSnkLcy5rq4g2YgEA/2jZbMseCzNHggpcN9HO3u0yWfDD
BUrPXdpLGc7H1ybWDnqiKgakftztd0bhJQ8My3+dgEIdPU+A/SJHbNNXDPvl
WIV3R7UwCW3iwL7oflpo1Aurphrl7LDjG9Y29i5E/t12wihqgQi8EVdiJx7M
LwiROhu+xOPovBZ0sD2IkxpJYy8QROd/XtUwPxMn0SKDfsj5AncOPU0k7HOB
HW/8PhNHZq7qht93Ahjb11CCsYbZnPPcqU8slEQNvjjCvynatnrrGzRLcx/w
nE5foFgoOCTVGYpAeLHrPsSjOTjCMSnM+RF8IZV9LTnsYW636ipori6CEVPP
Z+DIcaE9r3Drpl/DtuoyDCirfucldw6ZylLJXfSHOQ4YD8LbS7TPThPl1Q2p
2SRqnGkkGD0lpQZSWsV6C9mLYDywuwrj1K4Cj7B8EBqJDfaZVG/hT/qHx2sS
hMzEDi9x3u8NLC7S8LhLSG//T/Wbr95TNGsAlkqYh3NEQCoW4t0zxAVQ7EBS
FJMcU5+UjhQM7kD4zMcVEppR7HHxsaFXEeQroT765MnpUnGVmzHCi53lD0cU
j2BhQQg54dj8XBMFeBgPGPLo7QGltv+3rFqBPfMzJkSjVD4mQFuh8AsY9gms
SkzScI2/l2/rXcxpCYCN4dCgZWX1k6nU92USMpwom/H3ZPgsCOYk4jdGWsWl
6xdSMtS+gHRN0W2XSN0NlJEq9Ogq99J6g2XGCUiovIOwjDe7j7bNHNwJRvEV
CQFbVl30nQTY+6aLq6uFu8FT/ztis21OFCKDV0EpX9178ZoKcF4o2fNV5rdF
HiP/lgny76rahqFSGIr5BM0NxfL3XQkQbf/Slr0vWQx8z3v+wdMrBI86Q3J/
Xz9ElFykvhf/BDM+/gwRtP4T4Nq1BS069Kw0237VhBWtKFMZqs5iily3ETR4
fjxsEnTbTbQm600YuwIeVTIvMISVPmeVBn7R5Vtive6BdihLucyQRuM7aykU
w3h4QW4PHd99ev5dyh3tsUj4ttFGoeqHgv4dWPlYRp/JpB1Kl4e8n23tOwsx
w+NtveU95gCRIs5HZHAvr+I2SDqFSZtIYPaoc7D0B9fZAz5iORU2J/0rIR2S
TrcNf4Le/hP7XzMpThDDhP/LD/nGHFMWlxQ1uvQviQJf5xPhRf2DmggLDBFp
WVsOUPfe0C3kTmOxdSrUXy9+PIPDtjP788CUxlsFPlgDDtp+PaxUKxADCsV3
EIBF3qvPRguiXNZiYdoHUJiz2B9xeas2+thzhnGjZB1JLBTZyAJGK7zJH3sd
6uL0vMj+VJiaV8/6j9fLF1VZiqYiWhmTkMR6A2H+6dN2KKwaxfJi8/lxh8/0
a7WV9iN9cggwJcjcDmmiD0nLImak+tlbY9JZtPNXnbCw3XdJJtSWaZC2DuT/
xxu8mZqX49UYVuw5I3JdZxxmn05dkUWVXMvx2/4Akwec8yH/kIkBKMiO32+Q
hqv3rCfdgt6LkolkOA7SSpJjCInQ8kbdGQ+EMdfboNOO+oky+YMjrDXRkBLE
t12WZPdLqMf40jBOY5yX6tVfb/xnzL+YwDjIVVtofJHHuuNSjYyZCXrVEXRp
0rRYzPbqGPmv9poycoK4lPEDjKJf54tOfpxSK/UHUBAOhw+Ste4TWDWuD8W+
+uJUj1Vgw1JYEICzSysoo+3xRMsqpOFMEN65K+RHSJsZ0mWROTo44V8gm0HX
ahu6SzNWIH7WZiyImrCXwIjQ9Pzmgid6cBl8Ded5fIrudsZJ3/xDMo4p4tay
97lbmwoI3zmWBQoO+obk9lGrU2hS/uQlYcxHkBGVAQXvC5bCrf9mVLx5J8/0
z7XV1d+M3AQCxjn2Kc+4Xequ+570WwmRz8honii1OUFZNwdfp1xR9NL9Laog
05dZa9/91CcevJPTLNHrR04jxS+aOhriYj2/F+uCMeJ3Q4RG/m00SGvBHp4+
0hh630B/txaoJAanA9yvkkcjwpOYcD2ViwlnS5I7Vov1E/71eSrt0VJ1COdz
LylWlKlwXRixS0r0tfivnVA1sxEBJXYmp7IGBgeHTo1Cyg8ePOcLyme8vbz7
qyC4ui4GYJvQFcrq8BF4fiQmUs1iIEO+I7XLYkrjwXcO4u2yffkaJnzDs8mz
hDjmeCBQuuFKEWwrgKp9Nc9LFpp+0+Q9oubpZH33fgpeTaTBmWK6ERUlEP/9
IXY71Z+G2H2yJ1X9JJ1NG3wsyuwGN9Wi6+FfE3s3p8MSlc5C/XJY2jGH8bWU
EdVrVhsdZFT4v4X8S+rJuEaQOquwmwESmezXscHW0crAVk/5rdmKxwScVDTx
77vdLSgUWbtsctGHEA0uWo/Nj1mp6JPFbHfVUz5tpiRBvfkfnuGN1NzsTOwh
bNJ+DFdPoDPjLVQ/0KBv9rLph317Gyef8cRtJ+jLljbe8WQ2tKDgDGZP6rFn
O1uC/A3EnabDZb+c5vuwHr4EX+ViYiGm29GRNZ2esv4hif5JHY0CH1qAu/R7
1giJHj0M1KFsbefaMwbEtWL5pjgdbL+Av50gKxfX0qtr5AXCSZgUFhMSZKMp
X0dp/7ZO2GSt35CQkwz+OP2Trypqig6LEP81GUCWfBtpH0UL/OFymA70Fd9m
swf6oGZq0ccqfJXciPPm8+Z1hQTX6RCkrJwIgO3F3OddIz039h/ugNN3W0cJ
4mrqWcU0fs2Qdkil3wbwibT59zf3lnyefMWfbWs/ywtwn7E/eHr52q69TVr0
LXXXGy5d46PDPVIKwyAx25VsT8tnxHGMX4adYVSB9K171QsmTr4NUB6kM5xt
cXicvARMXYzkntIR5TMzcvBYFNETYQtvgmKOHs62AdJk5gmEnbvfl1maaBBR
Ro5ZCeZOF6bOUUE4NwahT1HZrwFCsD3g4tUMl+CJYcggW2F1w4IjyE3qZTZX
35j9I6yFDS/qozJMM2iDehJpqVGZyFxeOOoyiyW8aHeONqE0rC2gvZ1A7U2R
w4PjbuISVhWIc5GULYrMD/d0I1QVVe+VYiC1wBAvuXLNI00L/hku9aLWofVK
fBTU15dKxF6IVenJx1VnorVoY0JvGHAQRDczX4XhR4MYG8B71J7YKuMoekUG
5wWw5z1wsY6d8vMBh5+G6hPYw0wlZJLVIjt7y8RmY1zIthd4P85EEcfSZgxF
v6uIreT9y+lYZt0KjFAJWIiuPtr0DfughlqBbYRi0m3EOY+qNG8dGc83KaFL
VucBPk0oFFtSO3ReJgbScOBH7lbw3/kXCbfjtElpkZYeDGfVx1Skwl2XLH59
mJfK4mHzAHxg7WWVofkOdqIpjl2aYjOjJ3+czfoWeWaEox7mIZeUW//Ai/up
X0E8hX/B2PfJTWcnvqY4gqjD+SgPl9K4evIxSS/B8ZAoKpP02ARVSWk1I0Za
E0tMG8NeKsyI/3W2eDBV8QvJuyKjeO6g44jtm2CkAiRWioZMdfLln+qnqupP
ghnhRD3y7HADhDBevCGrP8kgt+/9NjVbn5/Mco48R9d4f/X8p4WT0aCz3BuS
MuZwJNDDpXi63aGy+BRH2DDeACEOzn9LrYPd5oHhxM286LMiDIfZ1ln98x2Y
pjaUn/42sAUYxqxkPvTsj8rtethQEAYxyCGzI5A5aeG6p0pSbsgAxdD6ii4k
nwtz+jiLrrPn4Y6KJJgWK5PBIWpIqDfEKsIiI58VrMOJph82ivUVg5yNyonJ
KJU0v3hXQvlNxk43cXsvI3xAI35UiJmlU8y+safLUNR6vPhsvQsvwK51v4hF
5lJee/SvFIArlYQCZVQjfTaukJWTcpGJsDsKpRBkwI6x56JVbAfGBm9mv7MK
Y2weTEoNCV8JlUK9oB9LYmBjR4ajPofmDpVF1hT9iRJSt+GmXPFy/0rY+mCY
HdAGcrSyCCz04bPCX6spH+XKuEvEe1lf9rEgoMSt7tIAtRdcTm4eqvkogh1r
HyqBTsjqExY7zKzdMQQRukxzsG3wKSW4adA7yqsuL8DaGfsZi3kmA5IY7Rb8
yo4h5Q+LsbilFv0k5BR/t5kdL3ti7Nkei+NXE2zchWGuoIQOXK21J5SBzO4J
N1Azk1cjaKmpM6h+QCsjuN1kigADDqiPzgfB+yWJ+Gl4YUV9TGKS9pP1QSE7
IgoedsgPZpPp6PGJjIiZP39fAszE8pgXgz7K5BeCIy0w0TFktjshEK6lHB97
jjP23SvShrc4LGBpcaOd6B/3kn5f8St2DQjZtnamPY2E1C7olnJm8WNLwVxa
LwQbFpDPeN1ylHCX/CfCqnHDVyJQiQvR1+xami/tiilIjGXQs+SXW+KUyxn9
VbBa2vHkJbdN7TB8WvpDgVsHnSmp8k58VzRXl2SyrUArGYV/6Jt2C4xMItNi
IZH0558OMynqB4eGUA6xecohw9tSNfyOaktLTC0V8Cji77vG6Z0eJ51G3TyF
AtdS/X7pVZPRiB/eIzVtBF6oubQO/07VR+nhfum9teUoMIoqkDSwHYvxPldS
sBcVsjbevE47iFwDr2mhDQQVYRVQLDhnquJcqUnGj/83GJNJ4Vfv922ScnM+
oQULMcFuD2Iw1iMUIc8POujjwo0pFQTbeupHfpF6l5EHcgNZOLOs3NaePmfF
nOJy39sFVxpSM4YuWo03P7NF/qPc7VyFieYV3hexm4fKqX1ENZgmLNv9saJW
uBdELrUf1VrChKyUY08nav/tos8fCeiSHlgigp6HlpImIzFGeRwhbgAl37C7
Fz69QwZquuSDe6jFKUqyhyzVmx5lhenj83dgFezmuIt7KDX5gQhYLGsCe9Zt
UdEPa8qFcVWECI52009Q65SATxwz5pD5p1BcVFtua3k1tzkHz+untxG7Pqbv
p/Lyp1FMdlcOKBuBHYFeuxXDJe2mQ0mi9yPrTck727OB0ZL5DFSeNgeUq1gi
UfX4qIuw+MKZ5s3HtnekRLCBfiEb1eaWKRettgUI8Jo3Y2S5C8Q9wl10wtHP
OQwnpsUB5DzgErf90HudRXJZwVgc3bfM0Jq0pDvCa6H5SqMmuTX8P27RjDiD
A3/IO0Xmjuwnb/SPwN91Rc4DOZUHmRxMxLEGiChefRW0SpcJFLfPcECuWmvT
JcfErSrcsIjNt3Cb+tuokkly1SzvsGRSS01rqpZyqNZSrbOKyxqYg0Kgxewg
PagAuZxg8wakLF2ndGcgneKMK25dgG9zZxoeRef7N/lu8nSDWXXqC3soNzdu
8OlMCwwNTJSuSO2iqDsl8qOuBEvnzNoab9hW8O5MjBc67aK0q7IyKfVfAKym
P0NyO4SNWtP1eJsofd/bxXLkNeOVAfVKa4iy+iTOmZVREOlNVuTbHPz4E3ia
+D9yALCytRMHcPiCbgohpSo7KQK1VFkqAGzpaWDDTlgdTJtxt3/pVe9tq4I1
jftNMPrqQ72Ve2mpch84lEzagmTFWYqaj5a/+Q18D10kbysB9jdTPdA8Y5wX
A0COyOK3PLfqjvEYgvYMshmgFejc47eirz5ZkzHR6zvszKPFHJKOeEeGIKo2
AoT8rQzFebJ0lf+nHTOuLdFeHrYVoIf1JdFamjWMx3VfeQUXiQnAoyrQJhA5
rptUlp6JUpVNi8BepytpsI+tyV9LXL7PPsv201Qr9IJe3/TeNQMkrOBtCP0X
QMg8jzaJof7n3dVKqAOctvykTDR9iTFYkjO/od+tWIMW0F0twjx29UD0Yqzv
cC/OgFL6LxQk2io26uyo2pgr1s/S9tmUbtlKW4fPu8DGXciQTy4U9AZNTIVP
Wf4R5JVu7pT3eFpc2MoU10/FM/Ph5aF8fb3ctuUeguJ9B+0y2lDBd+F4Y1vw
iIeAj+c6x60a/J0anfnaJM+6z9P4EQst960xKTJZtx3vm6Akq+d5DTP9wzID
FrzsqltVIGXyAjgJgCUCBpnkhQ9Kfan4QRvMJIPOQJ+wQajsvVD1AtBs7bTk
D+NGx7Ygvh8VFzd/1wG6wlNXKuV5Uzk10x4sVII6AodFZB2yVOnJeAtgXhk5
2t7zaK4dFDHEvFnRRw54FmGe5CIUWmQ6Ttcr/heObf713HYkhdfryw4WI1Uv
vt/1wXyDfEBCCv4mnOmnjn0axrDZh1GXjw9mU9gOYFbCqk+Ago03uKgwqGQC
meRsPPiDUElQPqqcgDvQUemtto0qLa23IcFWmG/rbWmGRAft+gFbZHEFJSpM
cB/QDN+k5vzG294Fqv1XyJfe/mjSy9yRC01qkTje4Fu0uEAAQgbLr3pn9miq
wJHHrX9mATAvSU5J70Pz7QxqDpgn/iArfzp3sVEIugibyjMr/QdP+QaKROpo
QuGZehJRR62YOeeYI3MmhhB48GI0l9z5YifUTNd3BMm8teNDUTtlwGZU1xPN
lbRZYgva093Z2kAKB7IbYTX7v/8PY5SknHYaup3v1Bz7k51PJ+SlGKyYt/zD
BLmPIaGItAHDBEVftwHQw19sfYFqFx96aVrjP9bs2i1evzjs1sOOFKJVYAhS
xc7IberYOD1hNGSW6+lI6pQI9q8xBCkBcMIUg/f28QL7VlX196YiEMFJ5Pb9
g2yCXTHapcy2/Q6EW5Um4pgVW1LZF8AJi2usbaO+0kf48rtKW4OBTvt/hR62
+8fEryLTeBHfvu+7pHXAH/0Kp4YT+xPNu76iafdiTNxJWMlP35rnw/5siP8m
BMWMONUjlX1mlFvsY6zRjJtbJ/agYTmU2h14VuNLgkMuwjS2LHwB0PWeDbDg
+93fiJ3lIhS45wxq3JiXP3YEkl08RJU02K10hvfQ0/q4q6RE9trAhDbXkWre
pjuwHvkQiyu4MJyG+b/oReu2THmMMbU/x7dENZ6xomcxXcW0au+NxgNl2Pon
Fmverc11+q5sYvJgNB/Vh7Vqrd2WEyNqeNmOVLYA91H2erHmiisdFc4kSUWZ
Kkt3qe7xCtT8ZaOCpfhm6n+rs81IwYSStqf9sa0p0Ly4/BiXAAsuboxMJqOS
FzJLJmXOjnedMa+UZKfngFz62nnG4OPb7o44A7SDzpnatYKaycKGyEIDSPT4
BQU0ItstM0L0lKH6G9f8c9fFq2VyMshcX210ArX4VHEuwWUiMLDP9bFIKh8u
lcH024aAZkRNV320rP8xBKCJbzQSB2QGivV8ClygHqReHGFhmzKdB1nQkm3d
NvIYgonRakBxBTPVx0nSsN60/G+MjESbT49Sli0wi6O2m0MYTPgQIVvt+iXc
W3vPVzegUGzO5SIY593qnvLX52IOXscpsf6/hn94dUdn5yig4CuABnReOQww
OzLYn+Qg1DsM6yBA4zeBY1sIf3Rh5M2WqbjPBQEbyCH0r3SStqova59aFhtN
nhlcRNyWjVmnP3MMTQ9gN0SZf8ueZAZUebIGl6YMr1zAu4b/fCQtZL/q3gFp
Kw2LXms9zPPmrXzO+RHVmnie0o/OOjxaWOdWvPRwe4u7fSk02S0Bk50tEAB2
pqV3sP9zIBUMhnX4xpMbLMhQY7YhlpLNtmt5zZBOszCTW0t7fHK1K/WD9kLc
JI1dSgCQMrwCiaSnGNQGM40zD5+AVhuo5BJm0Z20CrKAC8K92VuNuCUe8g9N
M98qZC/ug6ejZ43z475eI8RZDzuzhw+iCxTkV+n82rjmLXdwTukhbKaptjmK
XcbcMJo2GG9Yu+tu+KOuFFjzCeGke8HqJuE4dpRHT0lwZdyqt5336hX0rCaN
Y2V1vNED9rWQa7OY6kvY75ETkLhGBQBJd+kBoyHt9HshV8EuZa4ZzMDsmJRg
KC3J7B4Zn5ptbpsuNqREQk5GFlGdsAAVhaEJPm1V9uU2HPlQrDlCoG02nETd
DYDf5R19hD5TmJwnXirnGA1dmCo3+iUiW1/QDrx0r5TpcQyITUjqQYx9Rzxj
9wJGlq5FClir/Lpc4cCjnixxtV6F21DBDsEreO0DV4Wt5tuJDgI+fcueBhM5
3+h3pmxo0BwFNE6jGFxvBhd/DMq0hS4ZL0PPidvNfNgrVKbCVWOQLj11fwCs
7W6yqz7GmZakxeOtMIv7zI5BowaVZ8RmSEM5Nx1m8tSd9HnRKeJmuf22sj0+
gBNH03zqGdftQ10E3zUmY8jorNMW5VnwKPU4EJjd+MiOvFb+XeqOV3+Va1Ko
+BzBnK7P1c2J/6BIT2aPdOyPs4Nw+ZCAYqrOpEzveS31vxsAcOWVqqyUR8D4
qSnsOzKL0LOktiVOx5IMQliNwr5bxB3VcbTzfD0caA04PZU632CuZf4OwsMy
7/idxKO6sA8hvKvp9wwAw7DasBxolhY/h4k6fzbM/wl4vdAOECsqum/08Icy
TcrTQ0bPA6KAjJEZZDfucI+KXecONUdPxe5yRueiTeg5D4KQbRT3814KfwxS
wo2ft4FX+4sPponb6eYEhi+AiAxYUYJdhpT7zWT8ZHUlAIEW2+0DHYQshkAZ
/uaTuA9Sc6hs/JM7YneWtNPl45S4YMSgWvikKq8yb9noW52iHEWF70ziJfR8
YqhPCHTYDU1ykvqKsXRMJWsgqLXeUk1g4PRL6RitgCvQrhenhPWxzW7PteNn
xAztkmPC9kC0bexnRKCV3xpDmczinD+JJ0iiqJNyFeJNgaF03YgSEXOAF3a6
ZQbFUXwkurhnYb8nZlOjQsVHzh88YO+uYbIY1puxzlCMETjkZivt3ygScyiZ
PFhBIgulx7b9FWQW3c1F0X0j3xaaRNFNUANgxPyaemc4d5mxMUAGP6IK+bg+
ecuAundccMbrUzOKuNGbH19EbXjUZvf+T0Oys6xizozh04XrurrA47OGfLE/
rb33dTnNNhOiRx4j622rw9Xei9g94cQVgSi7wzdy5U/jM6gnzD1VYKendxu1
QmfSHkboi6uIaXvE/bus8x/JaMCLjo1/0kluI0EiqSM5ugPwBrMQUx4dpQg7
ewWPDQ0D2y14I8aLDEre7WDgIvmwv4aBfnfqtzUXL5+yCRAjatPkMTGbwhWv
Wf5k0Adc1wXaTl6nH2yYzUb8PtiOgu1MgNO3bAkDNst0Gp9eO2Nm/ZEKNVyJ
FhqZfrxOf5bt8WltGx2+2nUdQgkQ/yZPljH51eQL7LPld/vG23tB2tBkqM3C
mxkdlmxuQqLJFVdv8hIpz1leZucF+iP8hEMcWE0Vm4MzXXvchaLvvVgQgDJ0
s2GFI6IjMgphu+6iwpPyc9mVl8wmAhuyBRjGIt5YlPxVX7qjQXmeAElcgtkG
Fo4sn+anhEVAcLzbLLFPHisNzMl1LBrwy3PQoKy4CyGl3S9CcG1emQo5pqY0
Vb4GRIMkL/FpkiPEFoBFqowt9cnaGdKuEXlHXOBtIzq2bmsSmuhHt3QKFsif
e4NW6M32QJayt/1q6PbBnEnPj9BhJ1IlSc0sF9GbftlzhYIhmx3xCRi/tUHY
vT02OBqPUx9IHNits4QPqPcBEa5lMcF0RI29Yhc2KPqS5IdZF2qR5WUQDl8b
+2QkQaTU/3KMHrnic1gXqU2w/sEK1Fmb7N5Llbh73flPVxA6dv9UWvy/PpQ3
hOP4oQEWQmqb5daIm60MDqhTFLUbuHdeVK6B3ZfVtn40vVGoujkbHyuF9HpT
gCMUDUwDX+2xpKGsImlmHBgrN0+IpYiBUXpMYMvXdU+QHaqC5appjVsfOVVy
QCw9+61gJblMSHfG6H6+Fq11/rodJHwCJf6cwJlPW3NE5q2sqmdocdiaU1Ws
rF8TQFKPHU50YE9wSjzFG1P8gUUPUZlZFErI967H/fV366LUYK6pBGC7TlRk
Axeq+JPuVOrbXEHAuZc6NYpzYzvWKUvOM3gQOa+mZx94DfarM6AokYZkish7
CImJi2unXIpqfi6I3yWY+hTZwcOgibXbsKD6TEzWF3kTKhd1mujdsguXTfeJ
8+HIovj1vdNrUIE5PfQXbcA6CEKDt8mm6QF944HrMxQnmmN/dgwBWdf4R606
JcMNsWiaXETB4M/McjNxNfSOcCkvFoBd59tQ5qZr/8BLnwTV7DtvrNiQUqun
utpTTygj5XYmvRqrAhwiWH6Ui1REO4VG4s/dK3U/+Q9amVtrnYpaCQdOGKPg
/reiT/PV64EnkbrJqEFst0MowsE1P4r8gPPaEBBVeSWSdHiEzJDHJvMqZggI
XZ/f69VtMj6etele6BoiSNW0Mik7NRyhD3wxT4dA/A2ksftwMi/xpNfDElSZ
sW3yzar4Tdlvy+T+bd3X/ZADN4711eY/l1ZTDfiZXPxVMSYzUAtzdtyiEog7
zITRKrOYhpKRSJE+CSrMhc/AA/M0PCkInnYxHfyNvDhVRN65wDPPKDL/bY2h
UARdSWIRWb7/P9cAHezh73aBa+n/vRsJ48jcPyth1WRTkxW+UNGrCyCOGvYs
YyoPrH0znezRdWlh34CU6MivSEI+UGkbefFevmcN0EhWxGcYEMQFI4iNsO+Z
Rf9J7o06RR1OBguhZgkWF0mAhXZdNBIn+kCPALABtSCe8o+W4mNJI3xPLhrj
/FWq6IALxrrufVP+oTa3PXZUHd/F7UJnFtQaBM9IdegFGWtr6BwOOrgvTwTS
Sn7ktxWvqerIhsq5Lj9CXyGELScTxgD202H88Wkt92/TpONlb1snc/T0vTzJ
rw/l7lVCuT9hi5p6kNkRxCii4/L4MEZTHIB91p6LkWJ+Z8uQbqTKru56Yyiu
mFpa0pKyVWqEswqnulB3tYbii+BQvznAhqIociD80xj2o5MuYGiO5Yjk8GEF
QNR2Z8Pn5A9v2i1CDVoKe09jlDfvKX60UcP36WmQ6N00+DLFLQazLdSDqC2w
Jk5/81Io8s1t1UK5BuyrN28G5VAMJxbT5I6x0+T8d+C0CK/ZZuGclWVtf0/K
uwTgq78Exbw7LnswEA6QRUAYjODrTUPhk54Q9kSoltVYVoSGOZpawAKHkZCu
YXDVgDhZ6xJRMwUafvfSTbKjSWKGeP3creVfQ8Iecw08idZ2mY1UnB6zFVFt
ZY6qmlZXMHlA12nPf6cuAhLI+OcAoshpxMJ0uXYKDT9KdBUmm/G6aFn2244Q
8FSBIqvxm4xHIbCi6Z94wBPi9S2IsLgC3RdJIWqk6ReDyrBotAt6Lskr6LaU
WpJvz5yJJewBjZhjcnWZ198lt0iHhs9hpwGaX6cDJUFZbpAr7rG4re0j3qu/
Z4jP7VONZ3iTy8qD4mjUU0UG2wjd/qk0gqyr1TSpExx3o6E51I8JupAvvNUy
uo/vtGv8n5EBZTTMwwv+Rq9rIGky56xfkahUcnpXaJ4BGrcFW2msZUj8GXLB
cVt8K/38dF5FcGfMXGS1j9enroHUsO0uY4dhUsyqcV6cxXoQXvFmq/FmabG/
i4NUtUDJaiEv9AWgKh8zcpHgl8k2Ok/s1GONBO6u13MxzHOVwWyMgqC/TlZ0
sU7jbIqTrSL53lJlwTdE966f5Tknz6mYhcsdUUqtPk+3kIf/OI+8HFqj94WX
60wVKnXKR2rssi5bf0f/30helM+wps57xNwJunc4Cv7/CNwMogkjEXuYmr72
rr/aE7xvf+lGw0dmtWDdlPfPshi2OAti2e1uEB3T7oZgXC8URB2FR50joKON
JIYjirMzsQ1m0wr9rz95tdnz2ucbAIqUxSk73c37L4ymWQcuD+LxYOpDbYIC
Hcx5qSZ3w+aq4YYASii7zIg3m+9jKwBIJ+PrnMvPnXkLgE1eykyg6vb8ngUr
H+HA/EXgBTRmCkqP4BIiWp5bsTrzQ4syD8G5O1fEd6gPKOmzJqxitz5ISwyp
/QrcdpYSD+jfW1ZDLGdHzDqlhsj2VNgk8W+6ARKvJl42/VWcbJTIQzbjeXlO
m47ckDxBr7LGKqk6PEymZLEbzF0s71o4lUbZhnU9Z3pl10bXUabBIxh7h+yi
dl5Q/hL9yTD0ey5H1386oTLUg7Zwze2zHTpoXbU08hqdUSiRttbS13gaAdug
ej1Rx1faQ8onPSwo2VFtGpD3zXnSq8S5gC8b1X88wmupGQQGNt80gHDWCH25
TCq28vSmg1mF0mUdQG+lDWM+QCTbPntdWZJ4vnXRB2GJOw4ttT1Yh5B7y0uc
qZFw+WCSMT1MwzjNiVHvWE/SHa2XgadtDX2uvC2L4YLWlRO8j02RohMmLoQD
0kj3WBd/Y1p1UWT7Wun8S8HzSWGFxH8mo3KV37f+iMbxoPIIynCnnJ/FiI5s
fwIBOtxXEVx4lHUXsqCshFU236MD/sJZ0Q84NffBpY6ntdtltAMe2/TsJlHQ
peVou/uAI4ab2VREx/Uk+tvyan1OLXB1mKuviphXuPNA0dNga1vQ4ouENLR8
Ndw0TKPM4G33bqu7e5UC3eE+okh5xQKH4dTECVxb0rQQbTHHGzOxQMGPcrrR
U1u+SKgZ1mjl2fpw3w6k6g4gmH+DnLdvkidWxD4r4ypUhj/yjXct3f/CDZ6u
qDD51tFNjEqDoYgk9+M8DOY/ZZSdodVKCTNE5pYiizPjq7G3ETQm3rN/AbFx
/nUlcpy3yPdpUJduVcyXvjO32s1y9y56UnTnnV6/KebiMcL2NKzlOebxs/YR
pTMWrzMijsXakW4fiA+YTvm/J7pz6mb01FMs1DSwlyTby2MdfvfRIkXsURQQ
iemDXpyX6W88FZwQeAMxDg2oWZDhykU9wL/dxwu1z+QcKesmIRXbo+ReI08v
UUi0MBXmTWL+sw2GmPcg5fJq933E9+2Ds7vNErbsJK/ixky3UAJ1y9+UBw4o
07a/MgTGGNlA60n1uOOfclVYYHUs6t3+cNuKJXVKtjP1IpC2rVLy32PWlZpy
3HkzwBUhdtaUJ726dDcbMutOzO6Qx98isL6QcBT2S0qC2CqnOBNxqyyu5tFc
b8C5DiDZdufkY09YMpjYc1j3xduje07ffazc/oAkGbEb31m4JOOo7BvTz9sc
ON/jk7ktzMVANljov3dLRvlvOU/CjNbiDZ3OH6LCkkz+FUqhnhtftXKLugHK
5ulcrxAc74IEWBdFbm+Y6e/aouzD51I0TfZujFvJWfwyPVbs+a3l4wSbwJuw
T/k3yf/o/Fxs6J6J1bUmGYsBOVTs0eK+ifBotmyDGk2KTPBjhASzQlqiHQSM
IOUMR7UT1LCpHmlK162oXWDaZXrh0tGLPwwQ25b7OwJ+vc/f07cRCuOxCeJX
XPAJft9fdpL8y8IzbaT2oBwssmU8SEomZ3bjGeN4zdQmbU/PQAszTL9DBWMs
3DjXZZQbRwuEbSScIj5+tIkzXUOtqBdNUiCfzrbolc8CDB+Ayya5cA97YJ6T
QcnxSdEvu2Spy8xb+r5VfyfLdAEDiuyLmymdiZkHdQW6cJ64X6jZQqXoGIMj
IGDiOJFzCBD81Ct0f3FzZQ1N2AQdwCVeT7ERwzhiPMsglAmOrMx/g7PeqjyG
VAB+zBfMhIUB06G5zwA5lvF0BJL2unXHGL+TYSswoKI1CANPoaYHv+OHW0fr
8T4tbPsC3lvH29R0xM0kV/++i1GlVMCID5XjwmsN5N6lxoy0dIKEmcqGHJdV
uSlzxPOPDBQCjMwg0iYa1YhVzBN+EL8/0ssDuJ91PAQGX9DsAzEQ0Ewz1A5N
fg+SNM0F/fLQwUld6nCuFLhTNI7R1D8BOeCK4gsNPiry5EDrC81eMCkeh63W
vicjMt5CJI5GbRtrvHaTJMeDMpae36VU8Sd77oIySpmJC346WrAsw1dyKd0n
sEUupF0fzGhhAA0NEqDeI/+hGzVKkk01F0w59xUd/n417b9VSyaqpo0DFOMZ
kZ5iAsL+aOsi4hSF1MwBxViZEe2wcbxPOStIv7aMFz8fc9usifOsOihMjOQM
DmorF3kns1QoGcskP6AEXiItEiBRLGjn+Fp369H4lrd0Zm+LAB7rYeR5SV9F
arZt44lpr6vgRWlByVlkNiJCHd5gc1IaNO/XKv+HZkj32Ds7zs2NUFV6kn84
XinatysuHd/KI9tKGU8H/n2bu3r6g1Z4a+S97cZ6Qlyxp827CF11+Xg895bx
6+s2/KXGrJTarx3WAsGhP091u786B2oLwl/zUq+dGwbADXL2z+Y/QC5ddW7a
gAxNas73f8Nl6+enTp6ZIXBtw+cKwkwP5PiY7b4yx+xhoc2LK9HizlmEDhRT
H3wscgdqzmA3HfYPooyxyYTuFS/COkD55UWa3EMrwR7XYL6u5UP9Cfgd2PoJ
LpjaxbEmnlZsLAZ5M0xj9w4g43JTz494tgmO0VoJJ1DuIDinEIN560e5Q0XU
4GbZ1W3BOyyLBafLKsVhwr1WAY1AtJ+gJX6/nUXdMLfAdJBTVovxs1ijDpce
22sY0AQvEza2LoKersaW1z2jXb4kbNm5PmUryBYYd28fage7J7BNIDw4Tfl7
ltUuEia+IS8kcUvcefHM3a+uxRoSeCZErRv96gP6hHlWydAmyc3+mjhRIxa+
0BC5jIc2gDz10XGLZ0ZUJvr2ghjKELSQ4tJOO3IZr0zr2xgSaplY9rVR57B1
Zq7Dh/t/CIW+nlIoOyDnwDUINOKQBjhv+gOpOY+dO8w9DkyfQ+WBp5l6bNqt
uSdkhAnVg3HXQWBqkS1+NyDIVoX3AFd9mWOCAEmU70aHWhYD7gTRyFBQBQaz
ZM+m29k86INAmY0DoqSOvxJWV0botVCJ0pAYWFWJlEOp/9gcBPx1TJtep1Nc
9Uj6ztDoQ/6Y7zw0te3LKzxL8qffHYBwBawGIsEXzk42GAnSNWPEIeQ8xuQW
qTxF3JV9XEiEPlYCD4mXZ6vjGREal7Xej7RP4ZlwJHdZpomk0J/scrQwdnWj
C9sITKtpySmlZP0HdAcm9dMhiWpbuAw3m4NS3w2WraDAyeA/7g57DYvaXzH5
iJla5wJOs0BJhaDnCF73mO/lJwXL1r+A4dyESVNqJr53P/l+KVPIyhdxN5zA
Xt1bByedvBtWRm7Stk38dc4WgH6O75uN1154+uyGJ3XUt+WSLlsQSaJEpkfk
ckdH/v32byb+BKBjnIgFe6vuxn8EDaZaK6bA4llecX1IZxfQRx06awdC9JSe
WmvJH0oMPiRk4sKmsrN+q1orzf+9M9MTWdlsG+so81r4UQMPtWeQveWYWnCo
gMZDjRUk7eMpxX2Opiw4LsICUfOj3SVw+nX2GkuE0S/K/B4SQ9zLz8faf3mJ
2H9eS1T3Lu0JDv/psO20MJPJV4u+h7+umVDNrfC1cLzbgN0ViMVn/WbNJs7W
aLoyXkeENpEthaUw4c3ld1U7EvVxeln8KWSZqR2iYBSp2vLq5qOpnB6L42Cs
4OTnOQbjkhN/OT8U8MQ58FtqcXWEBTLpCcIzUh9cOdWMyR/d6Dwzd/P/IAEe
yoAfiwklmGey8Cw3arCnHkK7szrY5RMaPkTbO95/8R/7BwWejRZnx6df+Tl7
8A6fy6uBC3XL5TNJLvCWn79XMQH6g4WRLj/yThKqJFDfQxNEnvTcH1x2Z0ZM
hjrKBU+rR9KD9onciI/vO0ov1yiZHrb6Qf5B0jNmoCq6V2l8oiruSngv8Ac9
gYOPpa+RC/hhyZDZEdx4Ft8ecq9Et+telaQ2fYPYDYPZ5sSU4SxIt91JekqT
2B612+GHdb/QAIdTQLoD5lKI745kWslGDWn/SUwbe1UOrvf4i445V8EY3lrb
Is2ydV9x7EiuY4tHvIqYwEK0c833VF8CFEQPRutZSm2Xgozl220EtzhdjLR8
0Zyh6I4crnWA57iD+tyWD/5p+Fl7OuRAt95sWMEBuAjugSNDcqfVNH/7qQhN
P1uLeb5qeOJ01zUk3FOYxicYfFWyTq8+3k1AeTmCLiNxOFlI/6o9ksaHc6+2
BSp68XDdq2uJ6n0yQ4rzcXR+7fuByu/YHfdSqmHSHutuvMlBKQ/Kfxguizls
+Car1+Ag353juy7k4e3pLHMm1LFxYOdoHW3Iq9IogoA7qhhAhQeDNXK9STpJ
fGieXeAix9RUIpUsu4EHTbw2qrexjTMu2bokaIghL0nrvAE1JffxCHwX3RP/
U4z2KxiWeBC0e94wI4CwF7gEMD+Uh9z78gjHVUTHRziLAuXVazSlk8+Pofjz
aoYNXcnHS5twBGdoRD2Q+Q6b4afwApaEGldyPINVhEBjLkOMAeyNs1eDZd4S
YjpSovdt4jrnUilSoxdiA35dMAkpBkO9nnQyIT+yjKnYKs09m40j9g3itn6k
F575c5ywkK6PEiyenmxDyRbr77JXP0nAbAEZXVHbBlkwWNN/PpvlvI1XX3ty
a+pYnajgr0Q8cDBvqdiPBzUZFnK4hevnuNRx3zfOvUyzimiYB08l4E4ztp1w
T90R6mkYSinyB4LeHuAxuC7yWH6XuUwBmeB5MsPPpk1bzJjUm67L0Yz/lTFO
abcRQt/DEzdMF4KKKZhaaCxr2iYJDWHXrkBNghsriPiyRXEYp+IlaKZLbQJn
Mo8B9sbvzhnAJCKfHQFb1ahZey4QgMvDk6l7do9DyUFuA7W4/2zFnVR86a/B
OoUyg5aahZDYmAT28Q0W1zCLHAsjmBEoUdnhbzHn95qdrDYHZx8M3rZmgDZi
8uwwEsLsvU02ICwDBPerPgM8VJSsW2LUQMqWkzxfER529R9ifryONlsYaYYF
kMhDsoML+9MEWvCDJ31fLYhmcW47OBvojgRdVht0thP+OgyfNrdPf/5YLV3B
g3r/JGRODO45+L8hdpjIzKIYMHHqbjVaQCeWs3WemMihOC40mcd6gPlWiIx1
LK9Hj/5xiixnpJc2NvxhuoDSMr1PqpGnyL5JEf/yO+llwycDHkxFoiJiFkn2
i1msPV9FEaSGUnXS3UzvQ3D7hA2G7AaywgLm2hHHMBxJ0aFXZZcMmYx2pST4
IYkOA/pUVaTn8vPLW8bbSqI/JippTbICH1wwoIlaW10vnlLY5T/E12TOnqMc
++ScoDnkDxjFVBaaAnCbrkc9QhBwY7bb5LFNr5PYuDx3h9ub0+OrCQaJaszQ
HfRlnNdI+4uBbu5dlBd1ZyahSYIKah0bJdIuqOHJOge1lV7AurNSsDZ8XFP0
OLjkfldAVDQua4R+l562IJmT2WivfiYZEuqpWTOToQ/fdvH7GxebIXw993mU
Sn+VQutKtVkEeL63FiCO4r4oTisE4KSuSymsMOo8x+hJaeQh+qS0nnQihoty
hJ88gFn2XZDWZY4IrQ9rQ/+WXaGIeOo8D/daekspN6xygCGwXwGb9KECiIFt
UymZUsBPYQVwpRmzL1xeog5ZgHniiVIum9rCBC9NSUh6x/4rix1n7hw1Eigr
DPH4Hh2h+ZIGdOdqxWJLBSs1xpeGPXXNwoJ8Ib0CdcNRv39XsDymijkfD3lh
zO4TjPC6Igo4oQFlepFRI6iwrqoZTQCEsV5x/AFBHNLc2A16VfT24JtrXFJX
WpJ72csMBlV9Y1vvYVDxfI0qI8Ca0zVfKfB1AE73goqCn8P6dh3NcdToFpM/
cI/Qe8l17QwjuPuDUTiFnwOcQMBH3+jzcynPEzmNGCXMSRueDod47I6t76Ce
eEt8G3g/Wyt/VoJtr7mMQC3urjDmSl/8OpdmP4xAgdF/lvaZDqtIUu145g6Y
nRf1LycHYhrBLper1fSADogVfdXmTXmu5CJEnw6AVYpRjRqg6CyJLTuvXzDq
/9muAxWyPJexL4CDtKRrGMxJGGfb/I2I6U20eS8VThhE4NqZD7fX5u7kq7MK
dkN2RvTb1oqtQR8mEEivH8ZWCkMsuXXkWSTsmh/wXYg+FlY0uO95Qn7INrq6
QFcqKmWmUgyPC6iU4orKzFJd+evn28o9P3nkPVKLSpWeU9/+Lniu4w18b6lw
4mAmsYXIZ/mTfpgEmn6difzpP1gphJVOZ8Ybv2IZ3aF1B3pjbHrPIy0abNqG
d+mqsADfnM/jUrH+2hw6NX1n7p2KHzGW4Xp6gmwjwRFWb15HmAqrtSrGOa2U
Sqor6i3IcMw2lyJWC10QyEaHRdX3DfOdyxr1jCv9Pjktpjmt4bVS9kaSm56z
Ciwpy1lhPdk7te1bUc2aSks3sg4VS4yV8tARletlowrfh1E9j2tmzNwfjQGA
YoWNPEoxamN/cHBhQ98Uavlfdw7eng7WfQvnz3k6VD/kXcH9/IPtPtVtk4UJ
cY7vIBzxwKdu9tRTQhvat728DCoT0510WUbJvxtYtuVHZKexJCKrVgBxPQ43
bRywkZ4s+uBqV4ZiUQRsAt4JuCQVPuHTHGf+KnqrBh7F0ulhjgcKg5+uy6eF
5GN+ACtUyYDemURrjg7kd+xRiCbbN2lKlUsWqnncyvtcieBl4r+gidaJANoF
nHy8mnn9tLI13eCeexdjStebRa5NUBNPIGwTmuyWaebf6xufs+SPw4VtTVyi
yUZpxeqrl6vPEjOhEMi0/A4B7t6WFGoJwXbuVxjh+KBc5wrA4zU9apXstTJd
+4YVw4kwic/66URqPHryC4cAoeI2thcoFnhT6xHfVeraOpRKFgwYhcfqLz6E
/loPoddRjtbiv8S7HrL2uXhQmt6igosfhWGFP4w0dQkh51R5PYFQvmR+x+j+
eweYcOKKZlbYtUwagR8/n++RKvmZsNvSbKKVN5tPDhz8GL+rmMX/IKQA1eVh
5JKlcD7xBMEnSly6a+r7ORZytP75Egf2C7OkPAVwagfdFGYcj99/5PcvIByY
b7+WrnS+QoE13KzcjMErAxjMEpSTp7Tj+Gu/lDM2OrLPbAXvRL+qoz9cGDeM
ct0M2E+fl1K0fv2ES+iMMbh6AB131lpTakqBWn0QLyaOHcFAmIDfhaBrpsgr
u4CklFp4m5ywZpews2S3D4QzTFuaer2pw3ZAa1VV9HNQBN5zm8hCKFCYXeyH
xOGK7TqWEfYjS6SLM//0qhfn8J5G3G91necCwOWtUnIrUYpF5Oeo41eR5T+k
MWR0q2DewJD81eYcurXmFtAa5mpmsBx5wgY473gADLT5lnuHFliFCeW67PPt
vXorD4J1624chjnlCWcVq5A2/Q7+NiSFHExh2KTpvXeAgnuo0OHBZTdfQExr
7RXh9Xp0DyONYza8NvNnjtMoBDxTfUyZGFxhd6ztaaYzaSPxw+MeE3uck3Ff
DemEiENQJQRbFoe5f3XtIzNE+PVYyop9tampPHf335qnL0NGJiyF4ysBnlbx
5domXAVR8LFeVQ+WYMhYUOWy8ECwQ0MGa/FYt73sBGROg8uY1b66d6OoS/Cm
dw/gphsFDPeGEJfu3mxHFzBf7aCyQw4EFFyvjgQyNrgMWzKI7qqU6DkbieLB
YusTfa+EcpP4oHoAoI99lCDZkfRw2zVOA2hv/mcFSRZgsVdTNPXOIq35KFNp
ND9OKDQce5RdJsobSaeMvA6qR/3xfISsIuNBCsc+tIV+93F6iXUxw98X8KH6
fq8DHWHyqZ8BdGWCY/CDu2/6K0TtKfi15fPnw/YKAstqWTfEfJff6T9e6TdG
kPQZlpquEpHICfhFetTa63h3LH8hBsoGOeeaxYLUQiGBGZfuUyBr9Ek+s3fe
kvnWCQvqUPo1REBEmNCxqy/9e9F1j3Uwm8aUoQcfC7vf16pEQS6aalbmFZsz
CuBl45DqaEtIoOhK6G7689x2pOuhRRuCFqyDetvFG2BLFkeAw8aPJwyyCtYS
BscovFTHkuIF6nI+xCo0z6AqhlNOHFugxgX93Ol0p8/ICiZQblrEPNTt/f31
8Fsx7mL9kqWu/1uB+/4WOaYOzD0nfPlGc3py3b3nfZgSWMsmqH4ECcc2rPau
TBvZXrkZQTYBwNPdazhhnq2t8DD4JRKXnOT2vUNa24L0EHeh28P29aIRMK8G
sXhoNxiQ7eN6TSMvzFyCrA9Q5p/PMofl2PuNLd4ykKb3SkhW6RuQJPgbNUz7
xwofk1eK6KsdOxEHqqKJ/lbRffE2RBNa3kWVaYsmTS/NCW61MBHdfZyB7Dam
nIOq4AZW9oTz5zFK3h/ZsFak/Lw1HRfz4VfQNxAUEDitIrFngnnt7CsrED/h
+cWsttPvl5HVe/DoAjLqdGmzs84OOa93zzCzLVAmt3V+r0FGw60I1LJC0GI2
LOz2tpCOvR/poeXZv56+lsxZ+c0QJRB1oabHRI6NTbimh50RX4Ahp39v1tcZ
D9Lb4AeeZ0tRNvzhJeCRJjTQOyQ9pZ14pOXIWC/2f2tw7AtX5kM67rsMMbPS
voU89GSq9NTHqJ9d9cXkQo08Yj4grIF0+c0BaHeo4VBEfDTYnhUExKCO2MYK
OwEqGzNEp8Tkr3MgFljmSRSXD6NRoAMfNBQ+t0u2LPCIGSchERBe/cYXKeJd
eyYGhy/dJW0EphVqazLKaUUqcaN1ioM9VXIth5068epJ6NbWAm8YICiPU4to
zXlbPvuX+0X9w/F7t+acdMqVm9V1f+2u5gupzE/CYmxHHZ8Qe6aZ+8spm70Z
FcL3GZtf2S/45iHNcQznmFgfix3ZWqeiNQvk4ChjRQ336nV8u4/TSFVG4wya
cS9pA36Nt1eWBv5A881/Ugqb9pAp0imOVZIM8ekEOqpPelEAlbDXub60Zt+O
Nw4iYL/UjG7OUP13qMJcsmKn7IrX7d5tBJNU2/PWqOpUihpEB4wXbntg7L6N
ZK3kDCgbzDTGxJZ4ehXSyjNdbzqZ486ZUm/smqmtoLA8lothlEo1wJgs9iPR
VYA18o80hRJoNOrIYQO9wN9+brL5Ke0BfPrTeOibcbemLwH7V9HAIpVR57G6
WL7mg65nCsd5Y1wmxZs0+3KcU8MyKZPMKmAHM8dVTvXVhGZqqqbSn170YWVt
2Xlot8f21nTPjZTr7BMxT+66vB0CnnDNI4HuCYL1bKf9+ZZNxXjTOMCyu/kz
QeoMBOf9IzwerNGtMSLAndgIOLkhbOCh4dW3kHnExbQn8xcFlwSqHVro1Ejp
1c89n52VmOPqJVN16pCV+OKvEkofd2yLW6x7f9rMFsteTwWwqpAMA29Zucp2
TncQnlHPkWd3cslzj+ojUjSjMqcW66uTpJNLGFkxhtUA7iy3fKD/Z2Kh0Ejt
PnjcaP8n5ITAh03ILHhgJLnO59XhJ3z1tfTzFVR6WGSvQPdkCzEEYoFK1tgK
oTXB12RkBobd833imgLH3WmAAdDlhfRcf5MT+4c8/Xw+RKhz+o625jZYftRi
wTBzMljkAdvp6BZvAh8mbY1kya86ldsn++2sq0Q7z6fTzFvX2roIIcd0pWlU
8ih0Sxz9TvTtvc7OZkKaiqpMRbLmpBxSl7dFDqytnyNnPu+TUetppyX3Swgb
1AtOqkyQYgfhjAgZCtkMNlFtiKY55WCfPwVRWoXHCucLDD5ITYlxGjbmTBl6
MKwXh4hmw35yctyeOpaCF74C4u+PnR4eCwPssnDeESIy1kyK+bPw4f0bcisq
b+GxmZM9DQtGMRo9cmfnmbhiLLL2XdU0irq+Ciie53OlSgtobUCCQ3z8UG7z
uitpuz3SJusulBQUDnBeeH46EFoLU/n0tcbo0qE1+pDpebrjEdL6O0fv3X90
Z/U1cA/lcsr2ryE+wWNnu+fhW+mXX29ELstZ8utXz8RyFwVZd3HnodEpEmD8
/Ad6AZJaWrGX++Qux9f8xBVs+eMI8RHTeLLNfINPb9bDOgkD/A2yojQalSjS
N/rJ39shoqftYzSeI3dQURWxP7LJmhWksDGZarTea2wwVfd7zbd2+xwFR6WG
0flGLJxKiN7+FMsK+g5ZbBul2SEjwUs1ejC6yc09nuHbmDsSf1PmYi0pe6v9
CswXecs01P039ZIR+dPTqcdshooL7abNW2gJStdm5UHVG20g2Phu+ot3Tb4T
qYfOn3Ypb/xEZGKqeWsWDgxeIRdKAgpx6NgFp7McGxTAgUQMgoKv4oIXbitX
ea9BlQQ3oEojv5fsxZn6KwpcbnDpo055tdCpShu83nQXW2gIgPLXYHFtgzhY
Jt3yljv8rFgZMioTzAwGcsEHv+1GUUUBHKPLozn4U1Rin9Qf5wUGONFgNRXz
PwLnMD9sUbtyhl9HZO3QLz/kIuK2HF89b6WJHkTHIe94uBgzDuuPMx2ZR/RF
Ai9Usrt25TvoajomPDQM8buvvMwzIAkak+9wkv3ZRiRA5KSDg0vMrNdQoI2c
IAaSdW8WbytBo5zG3LftF6cjywN1+H0d6j3C+s04nAWV6uINIata4ZCp/oJP
ZrK5VjFEEcOhrL7LG4TN5dude2iMt9x1xkLFL+XaODQee6b0cwKcoew20Y7q
+bwbLHH97GPv3IMcbNyXPwiVSuquGudc7uMVty55IPY5Pwnee8KPDMfUUpf7
GocNagOPQihp7GhXjSwfs38+SUL5vcoBzOxoHOAuafH5PZI1JvH2ozt3GGJu
vSSRVzTaK9L16dLsyg8QNZfHZbbNVOOX7W2ddKplCRwTqOtH9neSA3R82+W3
VKcmwCssNzVyUiW922X5J016jV4O8PdaYgnEaCVQH3ETJp7DIIcT8+oaTJZn
jL3k/Xi4AKBicuofyKQMgwKDG4Dt6gqj9cvsCH8tZZ2/SDhYQUG6pBOTS3gL
1v4SrhVf/xQdXy0WXMuXH1HFuxejzWLh+KSOeiKNiBkWuYUImtmAs9EqK9F8
USnnewDlA8nRqibThbW3l4H+3IhGKT/fKB5Ff3QTSHd4CLcIkXlosaQFF0c2
+oGY8L8+7DW6Z+yhgs35yv/e6WF3nEAmvDmeFZ5XbetMM3ynpmOQ8La5QFF6
oG/SfTElCnvFceIBthTaaET1rAGMNONUYbjB+MlsN6dTEhajVnPjCp2BJ3GT
vc6GNBlMp+nVVQi3YL1Rmr6eMSBYBsOlDhP7vyMSH2O73ejlRm98jvezDFjJ
hkYEwTl/ejzykHYLdjU0EyU9njHLiTfv9qJ2sqK+X6ns31uo/wwMqYuRsVjd
sYBvazvqNJiLF17Jm299fmIaIu2a9VujqcDJSKaDO/OnT5MhdFtSa2Txmbgz
mSUpyPiyjhkE7L/o1dCYZF0ogoZKAx2mgOiOA1vBzUZKZbCNj4Y1JX3gkfEK
KlaD7WoCpZLPI3ZPMdMw43zlH9AoKQ/LXXsPM5Wy9V2V3+avlj/b+XQjDZh5
73XLf4XZAHdG0089PTAUZTau5Xx0uVi2fwvJSPPGd3IR2f2aoIXihCNBzTrf
wilErqTNMcmLFgD1q+Dca1YiMmk4q6ZviTCEvZbZ0/c9BHOp9t8+hKs3PI1w
7L9zbz539oVZAv/5zKUlqAFoGfsjJP/4jd13pHjSAjrML/bTw/BEGgjJbF47
F5S4JwmwsuWbcZrCqFvXS/rT7WlWmYoiM4DNJs2qwxzW3Vd2SMWvkGPwQTII
B3gzMjRchiO1Lm11ttgDIstfUINTKayX5xLPdWBW8xDbunBo1Zyu1KAdpVjC
FhkzCCAhmuZTbrhIioGE/9QClHoyxpQ4ezhT46A7kHCI1lNOL9lMXdE3qncM
n1ISnUhuv/FglP9XPUlOBAivUwAAlbbMinERiII8fNErtmarIGgbLrIDmyGh
HA9IhSa1AF2xrvCG2bOYuZLtmSfBiAPOWIlTrQAyoc7Pbm5xPkNlEYWozfEP
E0DOK+cC8Ss3i0mBmxZPjCRQ5rCRjPCcpbA332emPxrNq6sL4tB6Tn6iTU0I
qv/ZrJa/uLcsR+oxsPyYyzIMJgf077YTqn/397YcTcl2W9MI4GSSMX24EwWa
XlB41QzjRw2tgCzsndYfapRsKo2dXvn03kc6IAIrm/JpieS6MDdC6vdyw8/h
sRcY3hEksQ7QS2stgFNzSi1UYuSnmJ8hB0LmV2sT9CZSu665/wslSA5SwXFo
1BfinQydgKXXCxHnUKCS4htmTvx9UISGezdGuSGUy7dqD0f5WJNNjmkmjk9z
/qMarH1pZSVhENHEafUdgdJ05a1k1plyMmo+rQFO+PyUCZ4T7T9LZLzpLo5C
WsWX9oanw6c6ELEgwzcfVRFibMDjqlkIVAmb6/wfQ3AmSN7aTkKfb3LCmkHY
VnvGf1GuTqw1bBWy2d7TgFqSyzUtxGxLGFiIH1FpkDGCfkBC75Cc/KNRf/6L
zP3UObU4N3Dfyq42VfbHd7PHTMttWGjUQ2x4IvVv+FW/dHu1ZucH8cJizQCh
TH5wnLDG0KBPn2l40WmfOEI+6zZhz9CW7kTPB0AeV0Xzk7Obp8Eo+c7S1oxW
JdLXzuqS4lLLRYHyCdRGsJLVty2la8Z937AHGRcujW9RbOQbPqMfTAzRt0B0
kwh8AMQRwVToeflRfmn+0hCoJZwjp3EUqhRIHPKL/wVA0I7gFUARKWc3R+UK
XprezjY6Y6Uoc2nG7bf3cYuVaoYjJ4lsii5hHz6g+PVWp6hUnSC5D87AHx/m
HseUy85D0ik38E4CDNzePrTG4vqKl4f3ZEzRz+KTU/v3876clmGiEX9jl/U1
2fTWN6PvMbsalFlOftXwj762jFifOzycv5nxOK0+T1WVYu9mKYlF64Zj2pnt
Jv+2FGhTUstrs4l1qUDN5PI2KUsohVErxzrWmqTRvWMewjBs6GIqMKP7cZdt
Wb6NwdaWUkqGy9f4sfryj7DxL04IsQt0WikbQfWHQgX0AJr40JjPpEC6vFYG
ylgKAoZniM89MYamfpGqsZbMD7xNyztDj0ikRZ+eK/xzOWjz1hRQlgpIE3cZ
br61RdTyVOvvN74J4hFNMSIv4MMHdSMKU7ofhZhlVTZfW2Hf/7XguWbxsbmp
CgYcbpxJWIzNf/NQPt9V/wJuqrVf3ixBNfozolOHAoTkp4I4gxyJKMd3Uk8B
CEDh8gsxEFfYgZHi8pwzsKAt57tDzHSD4PCjTSvitdYpLMxSqNsXVzD3bgoa
aiSEHs/t+yPUu6OrZy1+cC0rOcP2PKqE8J30oqlpoW1O4OGUXQj7I04HOiLv
6MNu+4OT8igzrTOa0Am7bO8TVXomIakLY04EsKzjUKuKzgQsS+fAocBGnuC1
FmDRxqISAq2+d/U7mCR3JgLu/kyerbFudvB6NqEM/3q6GpGKXIrMfvhqkW3p
LTwto2ohHtfqGXVQYXunN6IscTF9O9VIA4zy2x3XPZSoWS+cnmgjFt/sk1Pi
xvS9h1ls65OiyN0W2qgXnngmY2oX/8tGfTtzQN2AKmdnvXxOrSrWj81WCaDC
+Sp/9Eu6LVxrxsxYKVomf5Y11gvBpzcBqwd2nGk5tLfPiKcRsPEF3z8JlM6g
opuzh0LpGdKwVbDeN58ywCjfiwt1O18PSzqhWpLbQImTG+KeTfpVDRiddAqH
Lzp/hz87gE091YWOaVqmoyZVVm8fvbik6goQxQXrTHYKKDgh1ESmPG8bytWR
7DJjojfvng3gBCcnHajnnkdn54t3gGa5AYDn5H/IB0GbMGyk4ogS98a3CuKE
nk0KgL005DApobQAVGDEswe48kKzLyIsCp6mdBjcA1f0JT+A79yivYLYV/KT
04POtNYxyDnO/9DcaLC5mxGCSorpjGAGcKC1WKYnCCJo3VqYS6hrhFpAyhTX
OdVZ9Zr6eRMh2K5WEXNla9Cr7DCH0tA29kJpPdBySACN2assg5E54y/K4L2e
d9Nhlnzo/4qmSrpxdk0HXjO6wMEjCb6QL7Vesb9tIUTs4ft603keA+EEHsfx
3GmRs5Og9ZnMUZbYFFoztnjzsJGZRPyfHsiYeMbsj3BShTHz9z/QzO8oDiIr
Ueis4JTyQTtv++OfWhmeaJ+MTp3MTfb7iwYQa1XUGwMfGAjA8Dcwl8CAureW
f4WA5Jis7Dc+rpXESgrmqQxmF6BeLxs2SK9rMiDcgKNTq+mhpfRxO5iZHb/2
KDlRMhn/gqdVrKBOpviRnEY2MUP75q7gRa7yZkrLB5EpuK3lOHWLtUVfrR4q
gOtJPqWI1GQI5r5pw8jCGn5At+ixFyN+iJZgI4fwcggGxPfYHMOPmG67Lv0e
xXI9s71M0noNFXAUkpedVB8G4TCiUOOkmeeDRcNQpdJw7RHtuxOEgiQ1BagD
k9jCvh8fF0d7iOqZm/FKpiMJYdCzoQNRvETKCNNy/taYlZgj/X0P/mFs8KnI
aJjGT45VYbH8TgwzAf4uU72OrycsO4gX3OjxS4YsCS5KKmfVO3o9SJoZVohA
vwVYR95LI76bPcVLmiFEMSMv/8ziwLlKJbPUlSs5+4znBXeP1BmV0+PDl2V+
OhBSsTpGdFXTexm6WbUjFYIpCXSQfxqouSedTAYyDgplxu57h/KS/v6l++XA
bYSphLFmKX/oE1ZTpQYm3GismFBtNhZ/JH+hsXrbTAmStrcw2QJ9jLAvidna
MzpHPOPEv1KJLn4y4fvATt4mf9M+KtUasaQi+Nxe1N1tPHVk/7ISUtqL7u51
Dli88/78aDU1JSuwU3XaIN0dlS70Wud/4N7qHcJNRAGRtfag6cVUTxuacvFV
0hWdd2ZAow9Sv/jrVEwV83ArnHZOSrJ+DK91R7vbT2cP4V5IJkGKZzkqgGMp
ARDqwpzBOUreGUUOfZxTkW2uxBB14ppoejvOFYDmyo86fB0djm1Cx/QLptc9
rK/z7vZ2xt7Fv+DoWictVGZb2OP9LnmujiJiRyLZbH0/UyR72u3vHOpAl93e
m51TbRB+ZzDclCbayHvSAHoD2ud+gDqdAtTJte1CkE3qrWbtCSyi0dzz4iiR
Z/dCohDXmonUWXwiiWveSvidlYdomz+5g57gOqZIUpywjsYuoZ3lcU4hOZfi
kBzxkVldjFk3utRRL6Fk76UiqfZVD7/19fzBueTklnKjuAQJZDck428D6bTo
pUH63CzGEadrR5fuiYEtAs8yKuiO5+ndTD2SpqIYtMP5IQP6n8raeU6jNzUE
rHakRPFbfVQ9+xWBsKJU5wl2IIN3icRvZLqdIzJXlR8YgRsLmjcQWtwfIQ9/
UbW9WlJZ8AUdP4IhFTlOOkT+WQ5yfg+aHeOLpds/S7h0Fn0QSBChwR4HowIT
f++Rw3akU5/D8Y/McntfX/4obDnHZaQDTqo5cOk2TL9ygKbyrIBR96n1ENM6
AM/aOWaofZH+bQPbhiGrysCYqI7KCp/FxinCyrHOUax0ZZRhIsZWm6oM85ZO
kwQPqOp/3jEgl+kOt2PGIamwN50yXNqr/hkW3UqEKR/R3PYv1Q09bJHgp4eQ
sVP2uoAelSVN78aYjg9WfwcokhgaZbWEbz/1muWC7AHqlTVMssgadi0Rnwha
xP20kF1HtVVkjQFb+BQJAtNnQ+0bjPbFtoqnQNwY686cG26BK5FyxAFfc8U8
7RrvlyQaMD6eBUX25miNwRIP+RNE7lRKrheWeeCvmVyv8sZ54FW6AMF3bWDX
YpRc4jAsLWhIJE5ViQK2CwrGXq4Putim29wiLnwzqdrPqF5trwGNZZgnxXXZ
vrppC9l8uPDX/6hKbA+QPzBdibydbkgwJm8EcZxnviA/MLfdID1ry9PFHqPK
eQfAMPsvAV7kQn8P3CO5aLY664B43oxY6lvQcdsTD8D0rGrGhsA4xIT6YZiJ
ehRKjZqlmoJWOPyMxB8eLWVVb7ZePt+5TOJPtFImY5jPJcKNYCI6mLcs0TXW
tjDyChzGEY2ZXsjgXaD9mmpuapsP2WAVjmxsG/FX6x/aX/Kc9kzoj1sMvXn3
leSlxs3nF51o31DAkmxi2nsSbVcN3LFdAJz3qVTjbqR9LDHMUC2JKt+QNyJ/
9gPtPAPo0XXW4gLOucq7nblUrhOJaDN2REhi6OJaNF/z+6ALkCR9BuIv3+ZF
lUIdUF2W8F01DkkBZXhLzJsaFhktKYrNbL0EK5gNRmNG5328bVyz4QCFu4Df
JBr9cbil+lmg8qn3FV4+vic7h+hiqAfTPW7RhIEHHeyM1AUyX0NAcOGuaXad
bxd9xwfOI30mSLlMr75KbnsLrpz2gsfpOzKpicUBz8qd6J5jnQBQ7aqz2wkA
PTsAaiBKAQkaV8DiC3KIGcMZk1TEUpyxQaWb6xa0DuxbAwlOXsKaEt47P3fv
QKJ3L7CJCNwF4VAS/Nce+EybCJTWx8nkMw7if7k6HpkRHE45ag7SbmrQzms/
H7lYv6mljcgpwiB8iYqsXSEQXH3DtVyrt4FezH2krxkg3MlhwxddLMNCnDFk
z8lkQJWaIC5dOI6foMn6SVrZgOY/+HOSvpNjxOQkUks6gZXKPlXT16VMfogD
aJ48UdFEAhWS0hogl2ot2WPoq9tdhKoS9Ug+xK4Ip0cihMHxl/E8A8Hxm/Wz
CEoFimdm7AcMGPJsOS5t4N2CiVJD9ogj88ndLVmEqcnMS2QnvEABE7n4dd/V
o5WlnXpSa+2wQi+AMPhfqWRImRIjsJx3hqiPnv2DcZBv1S759EgPK8N7KepM
Y0I1daXhcPG0kQZdGwtH91nlsWw4czk9aHp9ub85a+VBaXvKz/WRZ3mNxKB7
2xqcQ9yyAkY/XlG2JftqRv0dXm6yzSPccXJYUk1Rup5O6415v/WTQ4nTbCsn
7VS0L/3Ogy6vN66CqhReVr1UifQwy9NeTQQI+QOEiHjDJWvTeZKDEjSqw36/
sXbNForJDPr2xTohCOnT7i5EPZCWWX7bYzOUjjXSW0mSTaf5bqs/TvXdTjsJ
QjNGFEUWeqwS6mYLYsZEsqRKHDSZbGKiq0damNc5tdUDpymoO+Ff88sSQlB2
a5MdINhFbt6U5Ixjr5qSDkRCr7hhnFaxkGbHLtRuzBkwJMrwaK3FtMCFe9ls
OALUP17JNkn99p2K+GeDia8/fB0Lpm2tp6dZ6qBY6xwxib6cqf5URsnbLJPx
RD5xBq/WO0N2YvJ21iM++Rq6vgGBHh9Es8IEDdX2UjY28AZROiPOvEtnD1bB
n4/hmYh8qZ1VZ+CyAPF9zSQt1TDh6OEwxJ95vnnA45di894CMtx0OdqdKxq+
PhsUOeXK7+c1Nrtdm3YPEUYfU9IF5gBNAk6mr70hAtXRRpvxKhGVMsAYtmT/
wskupXNQZW3GomKd5mczScU/OvB7WTfFEJgF+cmKPtDNq7mjD52ICqXLopNa
t2EeRwurpGcEu1eHI8qQsV326ZLe1u3heGMxZTpTGkbsGrug/OY1G0hemVA9
zGbGQ+P6ael1URuWEXgHJj44pXIdYOQ/UdbLY0b5eKb+Z8N0UyFh2IAqFWDR
0pL9b+LWWFf5LVBa8JicOQ867RSI5D1OVz7nYeF80fEETTiuPePDOGy3dYzT
7fUa6k8tRUfjQVzYE3+8egkZI03qav6brppQPayfXuU2mY07avu6tq19byXV
wfSwunnhGC7M8LuSYWg3CWYBdqldiuXci7fNWKkMUzSAu9eoWVUFsIP55KfI
IyBoJMwww9jAuz9aQlNmbFHLfQHfLDDrHkP08FGeU1Mt0ZfQ4f6pNKPTirVU
h8Ml7WM7Zr2pI7/iu98nLz7ym/lxFQp59FAQrASGpv4ryBlsfmBQPyca0J0a
XJwO930EZDCb+s60cw14dNeu7lscdU983LD3GdF/9DFOePKHIiOHR8KVNKyA
AU7IkiGcZSEFgoRoMIHZ5Rn/+5PXN3VCAwF9ADXUIod7isOR1p7GTktW/9cY
JR/ElFb2PFvXYVb5XaeynJxrOBXpsmVWwopRw0j/wjId+wxewVHLVU4/fXIX
BQ4qXnvIeAsxwbu85E4bmQv9SdL7IQjHiKr7h5NLKrRGtks9YEYktlpbwdUL
AlNJhsm93v1VIHOjfydY5pueMps6ZVl4LqtYnIESIG9wbim88L8WcyZaUNKX
V73QK3Q6Z2bwdeUVcUSGNJg57UKhiFivySg6JcqJGZDd7DyipTiM+BjzScXy
uPzUKF6Q96Ys7Ykjfl4+/+jJXolRt6bw3n3V1g+zig7phDaoz3XdAUcDfDOy
upeiwckZrY50Txv+yMgXdJBQSJlLG6eAU8i+GfToSFV7Msls6mtX37Xcwenj
gdUxLjpDZ5OUitQ/RR45ncxAMkSLOnOMnV/s5+JrLLccfFLDOAETqr/3zcki
0QsJ3imUx+gDcyazR+vzjuzILo0Botf0nYL1BCxuTMhzog5beVdqKruThQfy
qbUNRyW6uY6zqkb4vVjgFGFTKB7Uu8kFCPAkqTsG8w5HwOilWeUMcaC0sjF5
wJm5z3qlxjgDBCVZB/zWv602Y3ZZ4QKEglFiuswLSnOwWBckCODutmiyIyxa
PkUphCq6VXhhlBceaUtXbF1xN3Edm+tsKmxWOW33jGeKjg34IHHg/KqsgttM
pdtFO5F7cAMA4cGK3QdFZUtGk1ft6GTu+b1P7buYZ9erI3xz4B4iUXRMXmgN
Ym2dpUUxrfb8boPRvyA5pAo0lM5DI7klPNCwOYiW/hoyZxMVL7fR9SJePOXJ
K3NiPqFf4uVFbRKmXe7FaW4h4IN3IV0rvUcDMosTddSWk+bLfPd4uprErJ/F
jq7m1+w9qWHkYKrIWF3kSr6QTqIJ9ilrospkHznbOABt8vHR2v1sXimYyy8V
jyUerryp23L0MKo6ZD3PEI8JXd4bar9c65R8L90meNB0xE2EQrUd2J5xebCi
ttbub/vdZ+V/fM119LSY7VDmhg6bnXWL/i4POPmXS3HuozSa9I0WKYpBiNba
8aqHBtcR+XWThYW0tVkAIh8OUw02G/Uf0wEtqOcCCnJIu6h/Mj1UvzFkYyvt
9Kbsqsf2evWvr1JGm/DKHbBsDPhQ7pKi51xkeUCxjc6BEDhej9B2ER7e+vqV
WBTywD64/0o5C82sSI3fAVoDgIb3vhmeKsab2YaDchcepBsMOpJxhpgfUwYo
7H6rAqS/km/9hJYhKtgwtQYUCnXclinw/EFR7qCu+DhpXA7uYjF+X5vAOVGx
g+vPNO62fW7r5UxQGB3UayvWjFSYsfy4vEcMw6ONxr/3ek3ZBS9AdWl+TGCW
DSSOoWAr+xQpvrfEVIaxM4fwQNEDUDwnHFoflqR5VIQfvd1QCE8l8alsnDYs
uQaFNAhq5Tj4MEyjOrwSdZnGGmaUihS8CM2wsrrc4dQqi5pJDCbCJnYB2n06
PF880hWz6gwn5FO0rNvvYrsUYlH4PtWLr5NPAsnWizP8y5akBeXKc3tXVEf9
FyaIlIDlwxlwp42Qzq4apZvLFkudFIolR/pavdHGHDyZ0K848CcjJGABAuKB
6EPTtiBnxaPKwu/YWhL9Jayn9XbLcvBBXxlvUwn7h+Hrdj9gA8xyMWfSxqSP
hMqIushSMleGBnSqAcFYXzrDoN+FUMqh5ousPpCDP/snnRP4QKQ8AQ5n5ShV
s8sytMdlffw1N9pcv6vaeGwdr4SOGb2U5gOv1lMg/8tulPzboHb+d3GoisuR
CeMhx+UuZqSbTMfPTBlHjc87YOlgWyWJH3cxoUY2aUdahgBZ+Vq1R7zxbkjh
CyxL/AYnsfuT/sHKvH4jJ6j5fdfZM97ksJ2C+/ymFWi2Pu45xSpxKSVNVLoz
ZQjoXs5TwmDXJ7FYRFKHBb16E45pdO4xxlRiI00dzb7div5CcSJFMsfjxnDz
I6N8eGwBAVzUmKFUBM3VwJBa3Wf9ibkBePbkezcmyBOzkKgaqTucTAv1N88k
/9eqjMycaHhSINKVDt2XibFBldes8vrnNykIubKJy8/8gCohe63DiD74L6Ws
Oi8ejtgwjk2GoM7ZNO6EjtZKhTdWinelg2meCf/Y9br9p5OLHNr2HC38p2ON
jRFl52Ugl8it+WfCMbakNU/98D5L2mm9/7Uy0rR8Q4kp5cOSp1xaf1/D1lwk
CI3UjigUfc3d97Y4sO5zUkFJr0gvWDXNIUbSMXOCAzx2mqrPe780FbDEOGS0
fcfL8cmWWmGyE41M3/I9+gVmlGxc5h21Z+AnbTubNjvdepF2cSdBPQ7cPfZx
aJDNssD/XV8iUqC7hbR3n5wm0PTWZVsPqPrqipSoiL/EmdWLKc3ckLAkVc+9
ZXfNtRywkNiSnX1IqLVAD/vXz5aSZvov+U3Dmk9sAsnQK0nJvvb3WV9uzM7b
1cYZUQ28HExFlBkmBJ3w9NuahWBCkgwRmEPaMQCEwVF6Wb75JMmZTo81AyZf
Lkj4OWjYGFuh+RqsZjYN+FCc8IodERor41pd2+d2HhPZYDVgMERJQhlh8E9q
Id+mu4iHPWLdhsEeGL3UF1g2uJ26uC89XPRIzO/0VLYR29jbXYvUf69iXycy
G0heLt4DjHQ+8lCyqsHrr4axjL/Bmd6XwbKuhuO3FE4A1rhahJDgUHWLcsp+
q24X4o5zSYvtjnTcnv4fzYDNgR9mo7tNdAhT5DPz2v+eWkyYFZ/0ihjjNpKn
29vMArc4jGnmAMvjrtyi8vsPXjlL5qSfyXECTIUh3k/naNufX9qkdWWF6br6
trpOMvuuq+AYDxhPJ5ElDrI4BYTatMKSIiNuduZOfyxN7pyV1Q4NIuQm+7Fr
zfXw8mUCRsMoH5V6ZSH++5lyDJNTy3TvvomXeFcvVWNo68XBSitVACbh28RM
a2AuQpv+ooOXCFnF0Jz5677rbBkmg+GmkyH30CmldPaHNB/BNUGgRmxGB3JF
x25eCeuPFpw8sPSkq51oPxDnxYAwHCaW64YvS3BSh9miK6FxDRQZjKo6DZfg
8zBOU+berLNItNtNvwYXNQ/MktrnPI20+GzRbmvTsl8oeg5N2O9blaxy8qs8
tZazXpdQJMcgYeObYiDo4tf69Ks4t2tu3/pX9lvxq5x3swDiMPtneZn+pA32
pxQj5y7ssrFomH8jfvZpqjMns+NrqrQ2JKy/fRpcshIFRtHnrFgrLVe5c5GM
tHbXfBAvKP/qQkJOEz+PJpT4YKS1fsRXuHPxM2Ic6V442h3NTCLnKAuPd6wk
bhFKOBTmdhu4U6WY6xhfwoqc60D925AFFeZiszCGbtDSV++mygj/KQoO7316
rqBKqYJOVzirwgU0coGDhyKHx1mycF7jLZ8O5j0P9Ha3ocwTAx6MhJFlxu95
zvtRxYM654Zw33/SIPr48X99tuS0lVtPvtqpmLbfRaJKObK+T1j/OR4/cd4t
uVld5QAh2tW6DbEk5SIUL+CdC7EEHT4U98CLQAvsplUwXcs560QU4vAt6qhR
NvH/L7kjKJIdFFdcEawgbPF8g7wCrq7adl+nug9BuHIsq9SwaT9Ynghpi51Y
yX3P5IY0/3VEDiiT5U1aJkMcEk12HZUjdOZlhZnTakxX03xCvyx0+Ow411VX
LQW56XJRkE4ix2m0tO0gWKAZN0W8xsz9NtRdjJ92hzAgN9lV5wIvLrBUH+8o
Fc3aCLXvBpWDQyVVCVt9rrZz3eJ/tht+kJ1IxB8owojOVteQF7Bh6qZjeVtv
6iea9vzk0Manfw/fSI4MpeAxiVEatigitsymUa+6b1xKSbYjQhog1fVR6RqK
u9iKmrHdIjJq9r117edMdVBoyMxXni1+z+5i/bqL2wm8OIouCg24L9VhsoPY
7z9X14huBMtehtu9tKlRCLCPphf4Cu/eNwBSrrJfR/HJDeH9xCQ79DSMdXMS
R2bCM6p4j4vHHh/EntNz4PxEiaTO6aUb63gPads7E98HNPvBcOsMs3aEygBq
SKBPpJKmI6M2vD8VG9ZuoXf+EWPUz/FHUcLJFhLseiqPU5a+aHgZrCVRAHyB
/SNqhlWS2Lz3YSdyQkgjmn31A/TZ4l04T4M94UR3y1SBBUMsmLO5Z8E7xvP+
ofF60VopeEgq7JkaKO35gKOLpvqxe0NLiXIZkBF0qsyiPzMhWFi+JiWP4hbf
JcoAK67h2hJNs+P5VGgbR+dnWGf+cNMctBY5RsMVsLeSSS2sdAHFZXwd2F8G
uCTB5YsHskcsR54Ef8S3ppaYD9kRbaygy+dQM0TFRmpl4FzBacj1F64oYYr4
03sxUE77M3ZRSZAY6u/pQg8wPA/XuMSYTYhTUMAsdIEuwnKdolooyoZdbo9E
GDh8yBo+Ia4vNSmhK+d7iPULzjo8D6p36U2NHzxKM9g45u8r/f6RBLbfFt/s
dfz5nLepTjr7uCPmZ8XuAm5+aoNLpdr/m9o6/HNvqunfszTPAE1b/ieyrx92
reSl1v53HU7JGm51XkN1tW5iFm3ed00T5mCGZcCW38eeMBRUetw7UJjC6kVk
shwy+Ult+LI0VdRgV5++7dHPPkL9UhEqzuWOhLrhcPWMH/EpEGrdznRHb+sh
US0wY1dUP1m+nEXVLaN143IXIJoNEH/1Ed3pAzUmU0xezuo+yrMAS17/0nTH
+3+a9O2dghKyghvX/Q+ksIHpKGTUsV10Gs42RtxeWL+I8zsJI9z2Lwr2fWaG
ghfTWIp+8LMr8cDGKI3TE3kdDHUbapsVSUU9VpxahqQDXvLA1IDRjMK5hiS0
0rHxhqmkhsvC/5y+K4apQHpCJg9ABk1MO/Ea05/vq18HW15MqVzhuK13wdcx
3EInG/iVePVBq0++XDjsAvD6U7zjkjVmPYXCK3v6oCPEQNUOdW9sY6SGRjG2
0MyBUVgw96jUEyzUjunDO+tEbEGmzd/t+gdMYG/oCbMC+vL+hlvhrJhEh+AA
Ot23DNzPVfl8OIt6p/O3PAQtdv12yr0FN5OAPyJLe3FX/YJHddN7fvWUisBW
AkkdfoPOUPQ6BWVkwvd1VsUJ5+lAmPQDMzniZgioP3+8ml0s/bDRmBf5/Wgj
5MZYUGrueHsfa4I19cEF4INFRZo5dnN/UbchYfaybmh5Jwut+3PaphBMPA6q
LUHxqgjwN6SUbe17eD6GDguB0WTtLuWCnc7xTxGLRiS784k7iA+7ZG+8Xig7
NQkRhKjHyCcPNI2pbXonr8ougrq2kPyoejkDH8OfYs8zky3/jnlSMB0bzTfj
KFUsfdH5cgaJ84YhtEEJZ4BnMTl/ktAqoWraqgW/k6l8W73Nohu8SKQRmaqq
SEpDLNFmphcY7a/6EVn8i2rH82f9FbRITBjRCs9UmACeLkzoRyxasW+5Tf1R
H7xvzqyo8aQlL3/ClrWXk8z5hVEO0Mla59wAVyjDvBJ4IPPJRwxJL7roOXn1
3KcmFFHG1Lr3nK9ndC4j1RKCFIa2pMUbV2GdMp2wQrSMM8gOF0n8HuemQFF8
sGaFy/+tAwVWU5/oevSY5hTl0Brot6/dCnG5rmZoCsP9iGujZNXjshv35tiv
auKvOnfsJsKrV5TPK+1426MGDuwZkQdQmbJBFCeg7LCzn7LSa1M8Ryov9M0O
+ulWGcd9AA+s9SVrIKRPjjS1YDYmswub4NFXcfyMsU/A0O00oRRyJV3S4GKL
gveKmlqBwMgHz8Rk15YO+KpUuoiwvrODlRtdWRapRWix4lA1dRgCVjKwjpjB
mHaa1khtiuP8FKkQf986LdSpJbSWox9dAANG4EnMR4iUDEcK220Cw2CyBioQ
wfrY3PKVhxIDB7+MqUkVlGRBj+jk/NYya2oTtkXEVsmt70907A9PWZ7+a9S0
I+S/0m5bSgS6IIzXT6PkIAMyc6jgIiesrk1yMi8PRrF1/fPiurtvBgCQmU3D
4VW2z7a34hjLza529Zs5ccgeSawxg3dGBr5s6LFELpT+6sJndtvbxKXWNRB8
9Aq+3BvPxyZqjXeVThN9jFLVPojemJnz14B2kJiGX53vTKLCaAB4WTUq+3P/
DIWG4iOYHtzfAWqj8CBmilY2xZyLW7mL3gE+LbfAOQNKvijijBHfKZfiEc0B
p0FxOnPVXJQTikgfXysSlOCBCK2VLI+0nn0EBYrl6/aw9AgIcHuRJjfArki1
9xAeCf2dMpow/9Pdy4pBxiExvEWn1uQWyQwrjp5lbyHSG+sRmD8qjoQEjeiK
I4T+Lce94g6lONMnK3g0xe8Ql++VVPysdhNvtFTV4pyXKSouyAdpejO7WqGb
hvfhUYcmWVYbPsYYFEfzojeqE9FynGnBJLRZ1EgzYZ0XBYn9XRtomFmjRwOb
6aVllbf4n0teFSjb1djut1S2CFFLJj3kemdQxGhixh+nJy+a9NxXVE52Yzx1
RvavmysNMC8/4YvFn5bJaJNT0NGkFuesi+60JzccNbLwYxVz4hSR+hSn5ObL
75MbySCGvQfUfOfoyIz9Xzh234q0EAU+ZIZtoXIqyFagChNPdqgVJEdzpiFh
VaqYF/y8zEUlnaBangwRDVahzJ8msi4rznJnpMRx7RITvlMiuRdQvtyE64pB
Hy65Vz6t0WiugF/mSUv8OCNipYPhOnXB/2I+OsfkzK6uok4TyaC7GvkJvGHN
uB0qGZq0wSd/2eH1uepxyIw6O82t1UctCeTb1CME1D20KC2GxZeafPauv9J0
Npww0KiorAqGRBldS2Whwd9gaX80Egx5yIOGhxepmDlpkLZ6dm8C9TQq15/7
3DA0IlsWucbI3HPZ7aF4TrcsbwhaAKxEIFLFzzFFxjpn1w+hqvBP/F1Ls1re
mViXIOKDv8s87WP2TyRe9Nve2p6tAxnu6At9SYAc42eVmVyUznHgC5ZBdWiG
0aHmOPbgw5oTMBbZqkqpPzamiQqalWTmbE/GslwzIufUh+vXaiLE4fZUcSaU
bkqaH59UZGijwnp4v43Qade8x89o3M5sidGAHRYS5NytY1OTfJd00yb1MGc4
G8+vNF29p+5mDqd+kG6kvcnG0IO1p8edJmbLDTUPzazxhPmmhseXaEz6TF/3
xhRornYKn+H3Mthbw7wjHTOoJEg80TlHx6gaJypzYW+QcV6S3zSziiYyq6cR
zzLK7QXEjx5yyicfrF7BWSxwOjjqARAT4yM/dsSfOo1sJFBwXLpSUjQV6Pla
nxBCSLiskJxOE6lBX2kFMA06ABb6xs4ANU0rdfgEFeQT8FcOh/iu+WyVOJNp
RyZG+aG38Tijb82blJFosX+unjWJ7yOAKS3827l60aWCWmcdEDbgm/rs1UF9
+0zBYqfVeDF/fRYwY2C5aPtf948hbsPD4UdA9maibXB8AzWzcszHEJ+XopL0
4jzz1Z26FodShiX1otYnrL1xcNRB5S2ny76uf5eSRYWbpFsqRzA5QVUNA6Bn
Sa/Qz4bW1Nb+6UDUuVgKQBiUw9TYk/N/rtqE4o/G0A++QTJIp4ICt1DxOQpW
Bd6qgnk3k1l17rFv00YkfwbAGqWVP7XlDzxRoLeJ099Et3o3Vp216OKaiDyf
SumGCR0Pf3nqwp+nqqdWAy3GN/1N7BUTZ15lGlSoQi47buQVJWMz+8i8oiyR
CCm0G/rsmQTpOsibKk3S3R7fYgWtZora8gFRqsHgU8jeLitqnNMAEjjAsAp5
pKagqAwfQyo382iUFMRSDWxqFwELBoM9rbMpsqKcNWwWJyHwiK6yNzMKTOUH
R7mKO5kXt2isExPo3MIF+HKC6+s+4XHG5gLX3NuNNCSVv4L19OXBRIV/6oeO
cPOL/VE3UI26JafmGuxC4ktLAgMrck680pJaSldIcKEQg19sFvRhHzer5uq8
t8anK7aCGt6BttOXa70PkIyHAR10KlPjfGqGvy9bZV3USFS5ms81MaHPIrWw
ScDWWECeIA5/K6svT7qJ15NVSkuzmRIq4uiz8tDQsHQ3FzdTFPO20gVqECWB
ynXtsIDix21gbXlZ0D4zoMQaHmoua8wOX3TiNwVsy/7/Uc8RY1x5Bte47ClL
xDU767wGBuYWPp6bUEF7ZX5WFY+cbSrTHTI6ozJzohgbZx4mhR9Bi05JCh9D
YVEuC+SWpEVcTD1zcD9cJWeSx9tvDV16mPH2xLge6B6AKAEN1TamSKoeam5N
oboliGgGxjJaWIu0zjUez0X0LG3pg04yrXA/7T/O3tzy+Xs/jqa2acWD6Orh
h0PparAyqh0if0+u9zivm89QHvC+qgh6+21jmPsojUuj1BvsWMVEmyB/DXJg
BYadVMmoGFgddDjAk85fnVkPVBojM5npXEEYwaGNqcz0bpdA6zckRa/kUR11
cDZ29cFHe9DpERSvFpa0JY0KhCHY0nKSTTAvjm/q/9l8kKgpY/dmIDmy7vf1
cfZJ151hYRcbMd/SDvevJPyGE0fDZccH+AmObAgIamOlkLlBiOAiRqps8xUb
VBKQ0RZ21UwgRzrFpvz41GRIM8zJxRX0Z7/gWoKTPOOLVGOqTDgcbqDzFi6S
E9TsKRpD3IsyoKCcz57Nz4khcFdqr16Fbvn73NwEgsokZy5Sf+UpCrJ57XVU
tasf4O1Od2QK0YwlBkWt8JhKJ9gXtU34oCVmXS67xWGH7yDlZi9n28iMJ5Ws
pFmeXghM0mZe4abdYzdqvNoConYbq5M6ihcnFxzHw4Wk+wt0IEAFOWIKA57H
DDBtE1+8qTLUO2LJhra1Hrf33KeXWR5Ji6ROT3CUQOM+4mzooFl6voeMTh5/
QP1fg1UaGW3ZN8XQOjBjWzNe+8ZmNapZCEjg2hDkYUscAK00D/Ak4tEvW4/k
hkPrwNjmLmA95U6D4aO9LpHxnOW3hE+i7dZEty5Gs6ExPgKL/Gs1fm6doLt8
ShfqguYFj1bP7zE5ZJgyk6XlgYFK4gAIVMA/Oo5k1n/4wEEN95+sFIoBf2FG
Dq8x4Jk7ls8GRdwZYW+bBW+V0uRzatpqq/M99HlD2EsDNrDB5FVp2PZL8OmL
zBVSWasDR/m/pcoLY+ykMic02kR6SaN7lFzk/AYeV/b26qSqLT+LR9qGe08S
WopDPLkkXAtr3G7j+aPMDv+oYX3eG9PE+Tv1ZKkfFpLT327Ho2PFAI2N9RAd
UjJ7M1CQZ2a2WCXdlk+ozbyQk+dnWfwWaiT8kVJTV4Imv2r+xeCv3MvhxTjO
XH5X81BSuuC19I9qVzgTaQ8e/gkS3tko4wS1LVQyII1adUek1i6y7MiWwAr6
9Z8n3Eq/YZPTsHdyIFpdxbRjsQRYs1Mz5QXrb4kS1tOAVa/2NYtAHPdmRwZg
15DANjnQBSlJjQ0PKlSQCzWXddsc/u27rQ7dFm6Mm9/I+cW6wTmh2SMLaQxn
ApiDHNdgadhBeN1KK9/bfy2AjkZx3PZISwOkGTseWWAxd+jwSbf5arQ5zfU+
NzWi0iddt4MEvpIrbsoDwVQ6Wo5iz99myFC5bzjjCzBXc891TArMaLRZi9uo
I/ArRqfnt+i05fF3Lt9N+CSBkjnMhpwI+DzMiWMLKOOF0sJGfPuUkxGFsAF1
0lU26KeLiQhu1yohjTBJozHfZwZZNPRH4xGwLjRBjp8cB/obekNKDPTR8Kvb
tn9H7nrvltOhj3Nm2Io7rQetHgtrZOk8RxofuZVnJ4Rtdmg+nn+L3Dtfjtd8
qA22J/1GB1YU7eN4YHuVDGu725L5ARCERCtq7u2+j+ukbeQVsFRvi+jfEfeW
OEKTBQaywzcyYqibA5gzv3Qhr52IWIj7MDpFzadHR2F3/PHX9hzFxxsg+BZR
n4gQtKB/rXqFbrUtDDIA6Y9nQ8xXWJwLQHmJbSYZQ7fgPTnpFdP2ealaKhaY
QZ42QtF+jU1qwvPPmvvF5rFeqJ//AXJ9PvAlLbYroD6d5ZxubZ/2AjzloBs7
dhYHUajzY8UeCScvxU/19o/zpJ9PMm67XmzP4fpkHRn8tyXQQ8y/Q86o972v
B+IoZsTVZtDbvCGiFkgtrkKoBbf4vRtOjeJYOc2WMxGwhwmDbYr9TrWep5JU
3WjfqEEll0uh1ibKMu2cX4p5fmMJFxP0vB9yNLN84aD9y/clzOGyGL7XQtkU
R+mLweOpPgvqPikejjLHJsvcAlxoxxUwKpD366AUoQmZ4p+WrfmDpq67zlif
f6d0y993SbEvIdJ5yjrNuXQQR/on92TiA2jOGP5E6AH/MpUNBDhZpGevxDha
S0RWLMXp4uf9KrjdzetMfR4uXO0mQWSJwAAHkNhbDQEL5zViJJtlk1llT+bi
2eV7UrIKd3+x5S1GW9/1+YaVeG9/aHcLNW8AM+r6cNHVBU6uofdSRcl5F96g
BsDMnpv+tt2fPrJt5W2ayGMXLOvVYd/kkwBv4W8/hhOZABt7A8TlrOBtM447
0JrsPWT9SbMolrWO8++d5148IAUA4yCAeZSbdMEo8w96q9FFVHh+kbXePOSH
YfJZDOYReLseVXk0RBAvf+pPYZ8o7oYZ9gVrAAG2d6ouDHkwUDf8l/XJCyUy
MnwQ4xg53d53n64DsC1ZNE9Sr6zvuBgK+gjmW8XGUNf9EN3ZpG0ovxoKlK5U
qi7NojvCgrqWbxouVf6ID6D/BThSGEFfmBuIeKPYXuOVkGquMH3A7kDg8vDy
yNaOK30m4beoyohMaav+TZgBlwaH/yjPJ9+cqUW2YoGEkCc9NkJYtIqXEFO5
0Hrbrw5+4g1JqA8VPmTHgYjeduvj2F7dd5LwvElfnGY2U/o5WugWUFVNEW3p
JN3NoEtOXwn8xePuXMhdebAvxCJyhgFSyqMq1c+/M0mKz+0ZRPMbmdY6yOYE
Kkw3xzZxoDs7qKRZ8Tqgj5E4BabHTpI4Nw/NOB7diPy2PKAa2Jaxjmw6PUu/
HMiXpOFiYTPzeye5krDP3hVZnAfZsHQO/4AbQNzpPtwCADMK0TFV7hldseON
alDXyc0bwrq8J/VrEZLTHemlJnLWshfhSxNsh/ppet7EpSR1h3CJ4y4rs7RL
W0QzVwHg7hR7gay3DIb0KSfQsi+88GUhwdDuLSQMeIJxQ3DLBjKp7LC7Gs7q
Nvvd/e662hG2UGGVg4M42q9zhEZM4pvwkxUiZq8M6YQ0Yv1pp9U/nDhi8uS0
OMjTDhPN9DUuxWXJpqLdcfh/ZoBA1cbQKzpWIm8Hu+N4v3MrjJD+Zlt+FG96
5mDZshaoJds0n3vUkoDYQvP1kP5s8z8mDNia7EC1U4/2MsmAkOOgHDM8lxyG
kvCXeNhDYSKR9zIIczhAOCPLANJCRXHGRkkyaL3o+BgHXUnaiaIu85IOsBiF
MPmYfm8vgcj1aF5Mfmm+e7NhAKPa4jk6wCwkES/hOSKziiiE9OZhlLUGS0Rr
O/aOp4D1fZV4AzGJBBhiWSqS2nRr8d/HxyDqcS+F9LwwpJFsv5wNu/uVNqYm
BKiT6mWGB6oT6t+/y4SJjtPuQE2nhBfPd/jTd+guwTW85BNMw5QT0xK1BgV2
6C389lZYysbe1d/i/csZcTE95NSnKDXqRLKequrw+K/1PT5NJhP1FDRjZh4J
eAlxQidRMzd0rd0bJEMhiaug2u12FBV/SF6dApJRiQ1bGZNYL5tWAhKx4EEF
h8MXkioCo7Cq3n/UPUw9jZIefe3eXkpjmRlo3vTJfCNblmeiAOlB0HxgdN28
3NxxariAUG3b99DWsCiqwnc80DNSmohkPM5EqufOsflKTSEVea3qXLFZSUXp
Zx5OLIycG30N1Cen48Nt8dKnUIfRjfm0YpaVApZO0Zj5LsaQ3fYf5ZOuEcAf
l/RSdA+suxmKxQfpWtKAQLSVWbcnii1OjlO7zu3CQykEF9g/mtkIwSFsJjwi
GS3AIdCCQbZvwHvhb8kGCPOtg9CkMO2V5OD+mY7lNvsr/S1zVqbBdVKGzzK3
qpOvwLrBJZ+/Hpboh3ZYEhkbXLtAaIHDAOWGj/aCP/s7P3clpQ5iZktmbwJ8
+tuwIAHWCKq2HXqU4d7P95EZCM8lgfG7WnuLKu//q6FP+iBYfNIUVH24bhdY
DfTVWB6GkBINyFChWPcAqPjGD8YNouKzP7Are754dvvL35VB677fj9VFM78P
4Ub7DrntkzaazznhGw/SZ9hyqhIOd356E0D1bZZcqEWqAZ4QDJL+M/GJhb2h
K9jkLl/TZ+z0rHMF8cJ8d5saqdAHEkBMsgm4gRJ3ST04t35QRdY0FWoN5U7E
9S4jSCTiz65Bn4E7svNRXedz0KUu5IyJsesdgKIKXntEXswmH/B1wgKdMmgo
KDibUA+z5T0Z4Sj1KMgYF3VLiXlSb8YtKg0uZ+VIVMvazd91/8SCG7KYJn0G
27/TA/dnHQvruCG3Ax2WOYFuLhGuuKn2XcSOXtZqKGwDmMPcpCsQvfqqrA/9
9FHdSG2/R9X0kstKoYiE4LYPn7ZZSogKE1aLVoniSfsw9tY+JTEBhHOeFLNl
SwrV00OawlxslfukrYx2xJHKQxi6PfNgY1BWNDnYecRurh6w6EYSDWr+jtev
tRys5xdhW3mGk0aS2oKlAn5G1hA6mZ2iBrY6qAdm/CRCYUmAqxLg4QwqznK1
1GXUIcyGjdjuNnn5/3cWNKo2XGHlfuom4Al1sGMteuDQuHy0KAjoBnGsFlVM
Uz3TQLCQNnhp5i9niS1won1VDJHWBjjDTnzmxm8keGQKpxxDQQXS9+hRX5Pa
K45Leca/uNyLDigBoOqf/8D1NtyPXNroD4dslqbKh9ir/fW5wlqKgz280Tum
+gEyO4Vt95yn1UZnTrzsXy64PEt0+Sb1GQMS8pT6HRzGdQ3e0U/M9IP0bM7q
/JJgz+Bs1NwRKqGL/WNl9RRMz6VWobS1RL3QkNLj3IuyANtRmL4a10MF3fXZ
zDHZPUC4xn6rF952SL0TKlKJEZN3go5+5yNTcfnMgBfP/c8zQvfIxkOTOWDp
t7afmzaPTuoNL+zv2G+B++HUqyOdanAf2Qe8yXQNUFmap2O9ekSlckplMryA
uVTZCL30GS2NjocEoNiyjwXyQ7Kdlz5KJErEG3Kk9Nt1HG9fW76LZW6VwxEW
w9C/gRSjbiEkv7gs/5ZqGqxveFxPW6zo2YWhYnmzggv5hZV5Ne8coRgSYbqw
UM5at3qbrIj1hlJYdg9vDBKjDgKtoe/iko3GVGH9xJanAGNHSIsgu9mFresT
iMZUw5piR81jFosecH++k27hadIKfdtYP2uj5FNi1F3rZnblS6M2S1/rCkaI
4rLTrKGq5PnrQAF6RcnpzxW17gOeETlm4DAQp1oOezueUOV+B6bOS3uEdB84
alvoM87xLcuVogkeF0PNTuKkBIjVNVuFGNri2G+uWLCcqbHOy1cLN3UTPb20
avpc6nPOCkZB1rN4OqICCu+TDmR5o/89UkYfjrRyNm6zclrU7w3fruDRCbK2
naKsqa5fK0JKGfyvE87+6u9t6GaEqRCX1GEbWbZwOULjp5yExZzyNIyk/bnk
GfV3picdfJ6AZpXQOQQk2okP0QxIKj+se78Cuj3Th7u9Udbzhl6ZcQm3F98e
kY3E6MAetawuaOmTBIaOcYTaKmqlJ/Mp1kx3Uhpy3GprGfhbFZnO6GdTInuC
Ir0KFw49Pr7BIdWxdHWNYXisrURL/PbEl89ou87AEoywEmzmtxBnshCQVpoK
YtavdhoC3iCAT3EdvvdEEviL8m9B2Mk7Ncjh5giTFEeWQ0Mmoro4tSnjKqU6
5a36gZtvWG1LCwv7ahrgFBnAvK0PUQIknUxHVkeegz6sZu8VDC0lDjfIlfq3
80PlkJKISn/SGyfvQQBnFFW6L+kNXBzmcI4bO46R8SnchNTxY01nNOHilKfT
jDDmQYpDr0GlHbnnuSXNJRDACEHXu87v71WOJEF0Qxtu1gDTooPMb8KabxAv
eQzTZQRdFrtAqzZrksNMlgnZTHMDGzHq63yx2WhSiIv2nrPo/XUDDEfvVwMu
uOkoXPwlNQR82gAdDOKplGZPxzw8zgP5pZKerSu3bmGYhvBpPZ0kcRjxJpkb
HLGiLYPH0SzcvrrLACy9Qt8fwG20s3rDRqAB2cKZ/ajbY3Ad4JmN6N1Chten
Qi3rCf9hx4BMA/THULtwEhMFWROsj0uytKfm0AX6Zy8a1rRJz6zSQ2WDjp3i
Ope8J5N75rU1j6GqvHCeReX/WOLRCF2R0fpFPwX7x2204NxDIaS4y/+f8je7
Z2350c4vzNEQsYAIP+y4p6gFcI3Sfdjhej9k5YFdehiRJuKPK5vbbAIOS/TU
DukmJqixZdH6U3nLgu7wcz4nuIBZ6ne5IkUYc4XtHMKKR65vDRd0zlPTNRl3
vZj4B9zjIy2BQCdw49LelM2mIs8dfQmM2a4VHZx3CBwQcbtupDoqRJInEihi
8Ym0/Tq9bZdn5WffeM3gh7pzYPVSYILVKM0Eh8NZaTkg4KwAoKWNPdqSprA5
w8SInqV52s0xFiu2wVrPLivWFcxYNCzuIKpUlnZJyXkgrssKB6nJdYkyYfEU
IJmCoKp0k0t0NiQoMvSuhkGfNQJzMEOi6lcqREPwy5JPyHZV8ATErPiLGgNj
2UKRIDUhA5gJZnIBcgJ3zCgaZCOGrhygcIUDM52tIU85F7xlrPOhZDIfdSTN
VDYDA+Zxx/vhA4HkDSDypWJfRcDxnoAR4kDqduJDBlLCvdNWyw6EEHqavJ1V
twQKM4f9I3FcLbH43XtNVV6dfzNW2pr6F9eDMIbvoVNMsahfYAwSCsCdt0Wa
UGF9aoRxPQytjWUh5DXxOEb+tFdFnJ5ad2z5SeGlWx37BDpcxqabQghSFAWD
AVPkS27Xl2/DQNtuGploDwbiTssNc5W3luU02GPiPduTqprihkNzhxWkJbKL
5XUtwsiUzGpkfR/IG64NR6Nc5RrlPUnfo63zlNBildb8ZSmRJAGjFhzajecx
2BhKFwPjE+WjwDt2fU+Brt97Cq15E8k+/6jvJjY/caFreLsBhUTpVTbLapbu
CbackWxhdKMwHcGhIneqav4Dk0Anpn9mKw9hG8qiIO7I3pcz7qaeRPqKkd2h
qgV+2vwyiOJJe+Ikg9oiUypd+cpoMEbqZUC66712w5sP475tKIhKhKcjm5Vb
VV99/WOJPGg1oPswhUMID0QrerjthwijCCOVBnrg+K7bbNFpVCHppNqmrLdF
ltz/VUUkB3ejrchrVTuXxZ5r3UidlofhzaVv365sbOoB407IReekwmcZt27h
EIpBMAOd+lW7ehvV2/DIfOpHm3cFSzJ+FNkOJ3Bnkkay4Vz3dx2TIRt5AVyO
jOR7ZyaowH5dyaDeqHcLsOgHhvRfYI0SWElmpDDz4x0sH5vIErW0HISg6Dg5
vdqwTgrPVjXhmSNBwXxdIRLA90Xj0Ni/+JuQ2VK/bWh8ScrjSFqPMrjRvV+7
GepZ6ghajL7LbvVHm71ZC3Fb79EsAfF3bnWbgQMlGEoPxflf0hdAEqkmZlvX
+cWQMOllssWh9zLrQqZvX8+oztSeKhP31Kl993ceGrIdrskDW21qQKcN5GXh
WRCN7eQJOXtgG3NgEO8iXhatrl/lM4Do3g5QTGmSN9v86SXWtrDuNdibH5e9
AwlMZ6dEI0a4HMg/csi0TZ4whWsgarv8fvg/IY1zu0iguV3xYFH6LzK36ugP
ripHjZWcTGInz5o19qWM8/xDXb04Pu2tZoNrH/bnt9VWmt9G1UlAPbn/WEgS
0dh6l8IRjDTAXqr6eJcxEzXg2EPxBmMdYWqAczXdNdbYE9LY40L544UQD3q4
RMlElAKkF/Wf+SUPDlcdF6lxNTzS01h3jJX/k40h68ff7PH652ud3Bor2iFx
EBkTMhKTGjAl8oOvelC3gZLOffrSmvmov0n17emsVm2LSlsRg8gZq30jEpul
UGwwVSAiMe1BmB8htthF9r6dMporTC6iWNGcZlhWivyg3txcsyx1cjpVgC9Q
bdb3QAWT5AG/3pGXBJzrFNChu+h3ZIIX0q6DuZUIBr8Itrxz8G8776yH/AKp
H1+jeElKqjFvYknivD7oUW2kEg/zlg0Cm954HzhJxfcUdTCa/4mBl7dsjofE
1Hfel42eWFtd0LDUCogDdsUQiHUUpuJsbXGwdxAWD8LqLpVVwjtYP08Icmdx
Umq6P0QpWxhuJ2jofTR/WEMhJHRCwFLrZwdGjy3lWUnpxMyy34aCsFRhm9lm
UVUiK2eNGOOtz/7SpMn9Y2KKmOP4R6rOiHrZ63GFX+QB0vcJe0hd1bpjSCOr
EAlZYNLoI47JslSwz2YFcA8bjsoRVtVEVSyDHppESMssN+SN9PxQIf9yaFwz
SvC9UYce/Rs4Xou4Lcbdr/thIBehxS5HQWvgawSuRwLJfEJjI/pB009xDoDj
29/QaaZVyfV31NfupaoO6Rb8JAT+mXR0LAUgQ+AQZvlmngPuztqmmZ9+zcbF
JOFAda82PIAKpPO3ydrqRzhxsqMfi3GCQlf9rmKHmSE5U9hNFkWx03vlx8Lt
xF9pHOxdX8gbCfrKTCDoPV/vP2FEiV44KTo7sePQeeaYY3S8s26gU3b2r65T
Djh8fXxvaHNT+wyAEv1eh9GU0/CyfpvXc5kVOH9iaKdPyKh3U/QSYc8Khf2r
oR3Tvl2Fn7gTRH+DQa4k7mSlrn/fZ+kh+gYBOAHEhEciOJPh+VFpJayZUNy/
I5LYJhpzCXktbNs+rPPq++R8tvMfgPgbKgOczQ+MBFPfzq2mpZ++i7zgq6Ky
AxV2dvyCdFyriSoKBFLZz1bEFZrF/+7w0Kjv0O0voNXZm78ec84e1k/Ulf6Q
UGV6O+2pyPUFejfvRwsp5jHPjZdDhuGtOf2ND87r9XJglkT9VjTAI7PA7tx9
4uDha3ZK1TiS2BGB8hjCHb0uC/XEEOjDGtyMSeMi0W73uyBVmxLBZVT2nzKy
NXhtZU0szWPpUCmmujBFqt5r6LL2HBspzu9kjQeXeUtOXxDqwxE942E1TvWb
RH4b5dY4sw6t7MI43ihq/xfDF2RfwKB0b2LP0RcWq63lWta36tDBFFcBLHk1
xRPav/axnuaEcGNzgYZhYeDZH/GCoJeAm8m3FxZ2oEjeSlFIIJGNz+rZOA8V
LSX/wOle3e8mandUFju588vO5en0T9c7Lk5SU9ZGuaYyXb6P3aK59stYGUvx
cbrZ8xaPyAMwZYWNNS6gMUIkGvH/6NxCFgsmvt5klI8kdyomUeT4kjY5l3Oi
mz3yNjq4wFBm9aFbe+zSwL5rRgSLtGDVryYUariXyVAdJUis/qGgXV+GMxjC
pVNvfjLg7zYlTe874Q6+NiAjFmkCjQove/nEkzG5Bfv5wEjiNcYA2M+Q0Nnq
rBs2EzwQG0stzlFCsyazO74ZHWwKWkHD4a6FrSH+dHVgB0NsEoCYJHjCfPHK
CwX/1JXAhs2uJGqnPfzPlcCUwR1Hlli2M6/BOF9Fxfbq5pQ9LPn1z+pPYBOq
ykHYQwySfkTgakAiCtm7OAcfuS5LSxdEXyUdIA83Y7jjxQ1RL5BEWyl0egaY
jp0NGoOvipi+vmD0g+SmyQ3kivQ9zr3WxXqwbFD3rZZanjFwvGfxxXMyoGl9
wiQGn7uDQCU4np8T/1kCe6uTAyJtgTvkH5QlVbSq2pcYVm1vJnswtiPYQey7
HebpiPFkJOMPv8QAZmtdBVlGBP2LV8Kw5Q+cf47M5ttb2znXfeAAFtJTw6dW
pUxzZW1iTMP/yzls2JednGCSIO9u1OJ9vg8bgz25qdPuJZxBDCIDEgXjW3K6
59v2VEOvQLghcg9ABldgIR7Zt+/AE4PgbOaqB2b5BRBM/QSpYbyoW0RvkjFx
ycDyN5R0FGwngzxGaedStrVwAmKhodv/VD8mWb/kBqjxsNoQMN3hWwkUGfDE
4zOf13WgTgqIHe8hHN14e6GabQ+7QlNBThcGdjdKL6XifBfS9esPWRaL8+kF
UvSFxlgM9lmM97X4hjYDbOB4/+mVzlyBwPF6Lky2iIYKFw94d1phxNKNlu1m
gtQGN8pFaYC4Nd87B22tdqZfTIdezxBqyqXI4i+2554GYMGTkr0lsaJl/TCt
jjNiKCXPngXEuUDfEBfh2SE7VbnqcG5HG/i1xFq+3bGfbpxZs2xFvpaxDD/I
wSY0JJny2zkYQQVBPtPbZvarcBQNf7wmfws8gZvzRtqdN2gf0HS/K8lHA+tN
nmoTTuF3Q75HpEU5C0MULJSWtbzUKG8PVOqvleMO4fpXbq/QOJNq6mVTJ+si
s91D7eICsGmea9PAUAizu5qtdcZcKTtvlRtCEIpBhpDmpp4CsGjxZIOQpGHu
WIdm2IOhujk7UFbJnEaTB7WCR+Wj+gy3NES5CFSiKEPJXPezUzaGx7PVf7X2
5f/wvAlZXYKNvAIpgiiHtO0scCLTtFFnZ7tzU5hTcesAPvy1EWtTdMbEEW7m
3iBOI+jelb8OFSe0DDd66eG9EXksv6UTZj1CtKysn6Rf4dIbTFX3lyfXUQIl
i7+NLM2c9fvBU5v0k3h7vAha7VnpJvui9m3Y6FphRlNH5sr3x9PbeIC50IFS
lsh9n50xj92LASqkqz4Ob/6KzwN7EH6obzAuefy37mOakNt5uJkutLFo144z
Q88xm8kbr/Qbv590vhCaCVfAGrSdDQsAZ2B9yX06uJIRcoGOKqHI2KlBc8Lv
buTMQUdOWGYzKazQspcylv+lUqSlFkSkYUSCnZCbSKdfH6+dsecI4XTDca4G
9LePSin2bODtX7sr/CQ155cgSUm3//YCfcVH3Us8T0Oww5rT6JObzgEIQ/Ct
9JTRGjewx5ZBPAID50BoFBaNPrhixJax3y/ZRivgs7/8i4hO69w7ZrDwFOtz
hJRgn9Zl8wdR0BZGizY5KVqyFpHIdsKgICvSmYreUWroYDc/UWZWkkIv7Q0B
qiaKTEgpmwQeE3Q/g0BxoDSkyf37Qx4hbSQz8D/xxhS2B4fAvtn93UyFOzFi
fb8HryBcSggXVn6bnlvtI8cfpIbANyHpRodBRJ+jQ3wG0VfCxUtoC3Bvzjhg
Sr6BDQg4CK39llCM+bxSKCoTvO8f/mNnXSreae0amVoq/ASDqRxWfYzJEKT3
BS9togR0oi9aEfiEZMq2O3u/f6kZgppTr8KL5zRDXn/csbMjB7jXiqud3fAP
qeuEmt7KjXEMtJgOwyd/ROgw88WhshAeSrAv3JjkkuHyrK55IVYzDTwv4ouq
vBJLvu3vbKo1rxIEPCFVgY+xoIF8WOvtrRoIqMF/+DCZELA0ma+wtA0JmQUB
RSEwC4o039eZ3d2B7hN+dJQVxOqXyF4izWb9LL0RDV5BgPjTo47GppvsT+fx
xPSZ3X5of47CFP3xnyRvmW3rezaknNeBD6MaNvnNjdHtxJunu8rGx8pPLo6Q
ZqBeHlFNkJQpYviMwVDxcazeLYUcIxfh3D3epWpNnXtmoYP2Cg2IIsPdTAVz
ZsmrmoSZT10ylgVD/eP29b+BBEPUfLinTRWha9dQeD7jtBLvZ0q6aUhC7yVx
auZSD2X4cFWkvEYMcHsEG4fR5FmWTC2SGJZDQidmp6IOhbammKNzCWmaVwum
JKh2ffROEESrFX68iPdsN6QfMTaZpMKLwP7lxVIWxlEHmxf3o6y9PqXnTCMc
793tMd+f2xhMBnjWBxwopVHiRvHAuQVddsy0whMT43jCH/3oY9w4LTGmjC0P
Juo1puoBS2Ocg5SfeCKnDt8eW7BTsvuhOJXSYa/g+OXumpFITetN2xxbppiR
d+mI+vTDbJ/K6TLeS11CAfZEMesfe/fb2e/s4J66jFxkmZM4uftqk/lUevH6
nOMeBtVT0UxnB1o7tSAZGYRpU6UarildcuTOmNZNgtdR+Lr+NbXc/79d3eMQ
UJgaKULKradsrRjVUYJW4zEgkIbwEEDqCxVqp9WkxbHQLbj0jtcktvrHgYwE
xTcvvTOxFE82AMMsqou2Bx9PcAAjnXI3r+/CG0eKSz71Pq132xBDnV4Eq/LN
WGN1cR7vyn8mueR+n/UkGGay5EdotJ7uuTV6+NzPS9ku1Rnp6oCOQyI0m11b
dOE5QBawg3T6MWcm8lBqcCOXgp1umMe2spe/nk9hBpjkIjo8IY7DqpL63XlC
EyJWsYlRhDITEmuwx/ZU8fY1Ve263xD/Vaox7VwRbPgZShiQp5Z67OKY/Qkl
QZIBtAejVUq0C0zXDcxfpNSTl7tdHWbacUXLCEFomcEMQDjx/jv6/lNpN5Zk
BAeu8AjbFoaGYcSRoOW7suz1sRrl0V/vcqqMJTPlHDtwp3mwyHmS4346Lmco
KkuwoH1RQBrYrxnC2TpqMGAauCG/g1ge5nmAyaBpOWBnz27ePZNNwh+BhD4/
q+hV43UjfCixUUOyDYFF4FoaUlObp2z8YKnFGtTd9UReRikgLDqwbA9eDEss
Qgt7w5RNUBYbAzRddLTA/FMTM2+Hf9jX29cQ3Xp3vHZwib+TfNKJdw16fUxP
fbfg9NbUzPYTkHKinLKxBlGiDRoacQv+Vmc1+KoP9rMYvVWatrBH7Hl+DR1x
GkYmB+LmYVVZry5aWSSM0vjqPjv90z0tTz2x3mKhkxR91D0BPzTq7wAt4oN7
rqHCayKUB8JEw5zUzKsG/vfdUeELaLYMu0mQt1aRlvluEbSAqJJEvGADnZCn
op5JhtZ/cyrTR2Qxag02GFvfdgYIS+ym1Lu2BN+eGSuuBVmCZpDF0H7vxwZt
qOmazK/hiF0LiZqdoqmn6KR0N7wateclL7Mz0bulHcqxLkdbOo44o667qAx3
xmSmChYw4CFG6tl8zJQKdeawf49WQ44ygVPFKpx1LBk20ZimyKwu//AlYSdH
wlPEPsqNTZ+QyDOKAe38Sxnn5QjbHRhR6tujIyOlPBFpC0ojFNrDC/82Syqf
5v91oana85hDc5ETmFeUNCPS+XX3zrVoirkTc/yLqdUEfCYX5AKjGsTOyJEf
OcisKsQdxdOQ1FBf/hrjfB94dU0dVlvgf/CQBMQef1vJJjZm0R78+jlFuQSj
S7xHYbymulGfEHn834Ikzs2SFAuZWKxmxBfFsAr+1hZoNbSBvVp1OYQ9SD1V
9hsdwQJaqtUqwDKcxgpPQ4f4Q6jOunKRfp+8imv6xIQi5abhOQ+S+v0CWyV2
bXdmuaVXEdWh6zqWau2J4Ll1qNZAMWSAVo29q/6T76EqoZ7roA3lSXCInYEo
yb7+s8KSun9C23sOHx9oGaFDsi064zkeic6F1V/YR2J6Ab8gZkuI4+rSaeRW
PXmglWUWreiXZzYlfGf78/AJUVzvHb+F9Zn2aemGi5f/Y6k9yRvwXd2piJcR
78lVj9Z7f+Igmk1T69DEyZJPj6C4cvawl3xOerHytOZFc/XFOpgOV0qALi60
pN/osW7Q0AGcW2DKz5mZvaYpcnDWJd2lwnZYnWJUV59qSoOy/ievJHzOQYfM
0ah42wsinD9ShzKi6mOI+wygpuK9LRyVSnx/epmBNJrF0xGeblfrndwrd7dS
D4dZfi/0Q3BNHavN2zaYoW+FBjw7yeQWtLjFAM9PEB7xTqcaA/XP5N4JArbS
CowfG7pUDV0HJnrtlE0q0NgZn+MI5sbNYmAoktjRRkBrXD8sqzDoNXOAKyL5
VQe/kgX5okLdmCqEKwxvZi729Qm6m/NoICK2qwsAiI1SZO4AQ90TFau8+w1o
E6btsLcJfybN/prWt6xpdDMyFfbi3NKCbHXDuMjspuWohI4hreHeSCs4Giuq
4BvT9BnLQ1ntHNQbpWZ3DHYxbopXaBDxntwVgXyZ5q31rtShJnByJhZRsZR4
IS5tr1pWpazTe0T70t3KJ0ADwuS7kxzS/V/b8My3DUGm3SS788cRsbzPbbi/
30La/JuL74Hl6h4qerc7ROqKRb2geuZ1qtJfkBcPh908T2ONYzIXY/eGTj2P
YzI7t/VnuOJc6WGcXiq4Owm2kLtkq+NRv1jG6cc7xTes9J//ka+MmgeXn9LB
8reLODxxWpZZue1YR2RIj7mIaenA1D837DQgZ9MKWTqBCtnyhmRMMRpWItyf
1a906XZtGs4x433LMhXakI0K0Bq3YgHdhwts29w8jq6Ff/YxvmwdJpVSSAS8
loUnaCSM1Uxk0dVuyP4WYOOmQKGpLIS+89p8/MFrzhw7BYiGK5oK62kVFqar
C6pnOsModhLp8fmn1i1PLElimjgwQ4Q5DJfriB0qjtzQE++IeZOA5XPx86qE
a5Qco5utCX8O3z8Q7j3didQVMAvoBNYlKGJn7SWCui7EoOnGzD1m+moqubr5
voD4TlIxZszQH22oeAJQezijheRFsBOZlyMX1NZhOJ87oYTDTPCIMgldCpLh
H+8pDkmCVc0fIw2QnuBnsHpXAcSlZYao4+jON+jBU0ugZEoePkxW2Cdga5N/
1ga70m1BqFfNssWcTfTtgtOvAXpJqTEbzdg+NUyKQACPfv4ZOaDpNjr0YPdT
jgIFDRwn/Oy+orJF2+PTg+lzLdrUqePzqHA1RnXxD0Wl6s9qQj6NzBHIFqYp
pPFjemOvYGnaJyaDjSISBvuqoW5QPuuDdiUYrJ367RCBP+TiDwHLjYx1bBpG
uGmFK/pwyxbJOiblSqnyby9gMStTOUWLcbCjBJ9lli22AClIHcjAp9yOueY2
a4Xrgqv5QNUMnc/3DP9H9XmnrXnpMQkpwmsuGQ6pZwlW5CTGXH9hCLuD7QFi
1LTuSgwAlZqqa3zg/hyxOzgwLvZDmPtOQ9h1Fr0gbKFF/qShdcgxaKMLHpVb
ZTc+SvZ4pt3uwC4LZPVPhPgS6egzZWjYNNPv64KENkRacENJmeeOtKoYVdNg
F1qJprAQOaScdWyA/tJl//k+yxCBqT5YfWL8sF/G0h5ynm/xt4uTAaxShtiM
ymIWrQ0d2kN4Zmyd/r/iP/+Sl6FLkfEQw2ymJZNX46rrYFSdoODlbIW/zBCC
ijl3A6lQLvrIUK/uz9R3mpjbWeiLyEG/OuInA2n8XNV5po1JuJX/AMIOuNZz
Abb9pGq7VkdcETPDmBxmj9etSnKnQPqppxN1bTRet1mXfgZoxo1m+JQi7VqT
rjJg5TpHtyRWZ+EWbPEh/hZh3lVeOBd1uGqh5r/b3nbRJBAP6fW4Nl6w51+5
m3eV3+KhteC5GJth4npznyLmeW7IxZWEI09+0u1MLYBWAedeejSQVrTJsnJ8
c87xzE3Rbi8/rOsWFtexSsg97EgycY+nTvfWxsDDu/kboOJH1SpAhFSKPnlr
DtL2fbkqISfN/E3k/WVU5XkN35bEznLDBVQRwuaF7HumXw9OibYEuALFIt9T
XZ6+xqYEJJxxUkzkljPc2hZtWKf26JVYle95mWCyyJId2cv2QgpI7YzBnscz
N6ptJuf1lDBFA6cOM1ENdOKFX+cqvfTq2Tb/p2mhkzzdeIkQQkZIxdJpD3We
m/LNjI3zDtIE8Gjj5CnzVYdDjFTvUScff3ehiZxq3AwqKgdOg/iDptM03X49
weCbjYaZcU2REifkzWQ4H0asxLyXh4uDm1D4N2pzJrihF2Ub7TjSj1318ilf
Mu7nsIrEynIkYiSXPNZc6s562xOnp0gnDdogSQchSWhTtkITi+S0OMKtXayP
mrITnaY1vyDdI+EoZwIwBGDkn+PTzN3uukk4XkYxMXMLDkZA2sZXaSF9ug+Q
oSjbvAKMN/K5VDYOuaJ2cx2+o/Dtv0IcEvyM5qKQSRfZMId3SVnLK9T1q6GX
O8m8nfXW+lNMZz45oedBRz+rRgrNYG0OMOfC2l9QJjabwMaNBfe/W8ZH1aor
dbKo7OmpIaYuv3jra3GKn+cuLBZbxeJzW/RWYSdJpkzYxd3GLVre0ZmSZdcD
Q2RChkLgXyKrKyqTGIG+NEJxopDLGtLXV+xBUH2Olq7kSYwGlzTwEjF/FrQ7
eMlEnCGgw1MjfoKlAtnuhJaKl7kS/Hgcd3xuCOZ8oQpCbCgBomz1hANQe3Dr
srnjj8W5hM/2e3VRlD+fdvORphpaO2lp3IHDSO++AYLftxpe+4ZLXolUrolZ
faA8uK2Nmd50ITSKBcm5QVB1UsO3jOBWxuUgGs+KGmZ3xZtjbZKDTXJFIgTI
TM2c4xtX30zWWBrZulzWAiHXlBJtiDl+w1szu7AM84kka4xAbElj0JBm+Fed
NF5bB9cPj9T2aP4k8rD6iEXcxCpVEH3pQMfNwqgvPIfQYx9TEEgS2nz8OTAE
HUkZnWw+JDpblGjoZpOjK3DIbD14diQUGtGLCK5uOyNHlVAc5vqpSyWIjEzG
FXzISna+MeRG/bOTJHEhO45UjQn1hU3x3H3ocFP/wUml6qkSakKIJ67UgudJ
IXRBau+0Si7zaON6agUIHTf1BABBDfmdv+Oa+K19n+ZiW3VxVBXw6SGzKAw8
Ri7RX4VyIhgf+SJ1xD1VmT5qwARpwVRVScgv8U4gxNbaojyU2FG8Wcb0kw9l
BlBCjGJbRfHTuQQHTpsJ66WGwIcJDlFlwHgpvut73T+mYoqf/WJgzYi0iTUH
khTt7abmmxHrn7vUUQAc3Os2fBKMbeY6aTVJyNyfZDNdzJC1MxfLX2HUdHYk
TN0JUI97n0bj0RNix666SSGQpIxltCyZSnSWdghZ3v8G5YfSdrPEPZI8YUnK
q/7d7CCb8IYqY/t29u526ATm39uSO/VL5IcokUJ7nx6aPc6v2sa/5uTS4ka9
bfQTuYjSEa6jPdVATW6s8KF98ukpOWYlyx0xNouw0D2Y7InQEGzZvEIfhw+j
HEkxGFrBlTEmBjGt7OJfiuFIAQa/VB++lIn1CBIignFFCihspCQUQyvazfdv
zkR0Ns10GrzXB496BEGOTwTMC5Vd4q8xJTO37O8K5blr/LTgpZAPycroQx02
qqw6X5xeCGlF9fF8OoD5xEnZOQiEmqjIczZ7mYVW6lj9/7+CSqjeajfwQFFK
4eZgifHjy32xSi23nOivaDm5XBGr7b2p+5ktOaCuttu39IbIWoA0IvsURyst
LOFOy1gz2lhJ4EEJPqA4k3guEj1nx/BapSLa6SOkLpppVy7uMPmnCwkvcKw6
pWTRQl7yGXCEvuMSjHnnTqCVdECJroTE9MFEbtgKh945E/zP9XFmT/Pzv+KN
67UJwRswS3YkXX68KEaKJmZhboCgXvakLfduG51X9yq72jhklLvJtG5HdU6R
m9wTYJ/R3P3Wy2L5+NAFLEvopxkCrDyG3tJojpIIrnUWNeWvMC46DuTppJ0/
MsCUdbsTQOi0JDXC7Gzh9VjbIw9cqzRB0jGUouC9+beSSWfNWJwZc7Qunnvq
wFheEefG78jvTmQw6WeLY+40A+fRfYAZSNBWOmBPZpYOKy4XdIABgmC0x7FR
tpnv4xCAx0KBkpTQ6U1j5kP8ss9b9freXmjgPB+xlH2kxYHpBo3+NXOitFdS
cbF3Mn4cKovQaFFL3wolE3aRDb31lbnTf16OVxxkJPGXhnfFGcdWjIZIXCKq
izQACRWdj+J3UjV2hAkCQde52WNT1Es2UmPh2JOm/80R0qZ1Vo7Cu3nRoDYi
p0b9isy0WBIrlOKykwtytr/Pq4c1v2xfo67KMbSXafhcv65U4PL2QTRzYLB/
7StTJRw01w2/FGoTrjyUYnaKs2JirZCVWwnIj+/IaMxipPUaptNAjjZeC7RZ
Nd6Pyv7KNYVs8UtkhAmJazfyAwH07SGu6lBgELsw0DYCSCpsZdy5XjiJktWB
N8vptclSIJ/wKkC7BKkhHDVffChgCpUZWvYuWnof1aYOrm5nCqGn3v95sYml
mc0y2k2nrhzbadlSE9g2FCO0C3BMqWBnT7dt3IvoMOBuP2dEMbBe588H9bIp
TgmsEIkNWU9T+9c72ndc9G6BLFZ3q7gy8WbbrfOPN1MMwL1CLPL/sHO6PfJH
j1bdlMlZ9ScWQAWpp/FgH9X5h3/DN1Xd8a7i4c1Cp+fXJHn52MBqCi5Tj5Mu
5StBsIrLhPqoqojf7PbPxGFWvJyw+TnfuqFtLY2+QCC9tbWLsIgFK9pUML/s
WZeWifu/3AN05ynUCHRFjG9QeLlnIzDJmUuELc15PT1Vhu08x5mw4pRFDNdf
5enL6ZO9CR1ap22+LSlfkv4MMjzDHokuaVsy031y+8OkhGzCnHyjc5WOg5Nu
R9lHH8q/zWbu47GF9WfFCzKKuhnsepi7s6bIpHfv+rVOqT8TyGWTUh2MWpTK
y38l9y0qMAPdnykTwipbsyiCxFIHaUHbcL34h7FrGSGMyT1nJ4xRR1v1NAOY
qy3s+oKU1HSluzrOoU4frmvAhRvSpq/RRjuqgl1ECrYtHn5tFj2YXDoRxmk+
gGLAL4mqTBCwG/akV7WDSc6EU5KiUpmaivmkrZOV08fG6A9r3pYUfC1wRcYa
UstNg9L7fPUEC65Z2R120a46Y9KZ+7V7ORU43Npcd7ZdIzzaZCfc4otDxLU7
T+wmoDnY1MfiCeY0EPkkdl0QJpm5hrW1yGsa7O9f81OfHqVS5cmHdJyS6QqN
5V+5WTLctNhKLG0SFU6gdKYevXBffncpkuZpi20sB51aTwLEDheaIUJiYj+0
P4rfr3rtNz2TFD3gJRMki92DnHYRnQq6RSQZA6D0SR9MrxnUht7uJfvUlyac
fN9DAwbDWDKtpBXPcmLY6HbN1PQ150YrHvFV8zsda8cvrQKz/RXZEfHdKmhj
DICFSt8y9HFi6EyrRzOZ+T95WOEvNIAWkdAb3gVKgnKw2xlxAiSRaeey2F2r
0aCUbXG0VZelwYN5ubosafiV+I5BJ9Qpmdl4bXklsylDAhNNRgdLtVITmWFx
2WR5+dpmFkyg08BZFF+NA8dekGeT+q0Zq4FzwjRQocsb9v4ba2zb6cGOaV+s
TbXmcuTll8g6O8w8j2pBqOkKcGZjMM98n0YckPekIy0t+lKjjJDVAq5u1ngM
I2S51+oeuUA5dlBcM6zD/rXgOhZwQ/HzG6Phds9RLJfFFAZRbaRYKqyvWsb8
qebHY6V8JX9kcqFG/aPjfwt0qiaPPf1YPXrJl6IusT2Kq3bPX5F+F4U8W1vK
IJyRg8fGKvc18h+13tTuYaAW1Jd4mLCUDCpq2cvoavYgPabIQBPYSLtsUFfR
G3cdozNZkmPOVAQfxwIPqEy75WiWn8cq2sBF8x8rwUchOPqepr0NthmKwHfL
zypJY4jBvoZeqgYKOHG7rLpe1rZBzx1MUktHuUlz4vqn0W4IIP8CJvdfzD/N
S29nvqfw+mHxKRuQC/017QWlw2aWNTHeoM/f4S/ddjN3nn3u/NHr9s9vuuoR
wyscRDqFW+cxp0HixmvoSJy7v/velUlmCrpLfG1ZwBlnEwN3ludC5v6dqlZV
dTKtyHIzQSjK4w8Ti4BW7n9TWOSSpBXilnouOiy1O2MlZ3UrK0Zp66t+Zk3T
kxFaAJqerg/h+W6ASs5hwt69fS8m1cKZlpeZlN/qewwPhtPcO6VNGIwEdUTm
VH2l3X7P1eV3eeCsbdIIaIovvL1iYasBGwcY+dJ1eg2mVy7md7Z8N0ZQuSkC
G04eOFXXEo/NxiuhZ+pzB1cCvq6A26S5EH7C6LgmhLVq6MNA3igDcB55DyjC
bZEwPv3nH0SeY+F2/NEgkOL+cYxF6RBSMdqT2axpCMzh1Knl2d74kSRnFFb7
TbheGXMuVbxXiNHpcvK/ODMs9tcPPPScPTAthCt5xXUkhLdIENCbIClRATei
CK6NjdezhXaATllckWRQuLEuED9Lvtppa0bJ6rYc6zceCBCu3J+5BXGWC5QF
+3BtJVOdlGNFS7drVvN6cyhWpdkPL3NNYbIMQ0t75TE53DlsnidShc+S9CnZ
SbXAg53ZOxdVvgsjGxy+bZSCXRtK9ge4tIM5KZ0vTXdyugVdQBDR1qd44GDC
XL6zozAglxzSAyBPAH/sTVfoQhHkw5i7ANoclqDsVwY614qO1OLuyLfcSX16
FBysna6ib4oLJewFOU2J7HQrUTF8ZvcB9+2u8pIVCcv+MR0YVX7Iv33jnTwS
ozwOJ6jc8ZSvOXS4Z1nyixLX+oKhh3ixUkAXtgC+KrzKp7lG+RCVpE0zOVP7
ngYvYPlJQIhQtC3NfDSQpBcWWGtG4y/E2oE9KZxBVN8MGDw0gqUac0ydqNwm
1hYjmKGGaV7iJnP+j8Rq/qWcXuto8LJmg2ZWMAS+WT9ez2nTuiK1ffDcMRYs
kgdnMGy3oTUAOL1PHatG3DEA/pwnhPsV5Teiy8i/0hIyIS9dYptT+u42+5FD
Q3KITQx22e0BBDJ8tYR2c5aFN1eqlnD3XkwK9UE2B5ohEAYciz/SG1ymU1yK
kT3L0+HD+LcejqhzaVRu5PLfXmbLqmUuqC6yIPEkCwMz1C4IEBIBY0D8x5td
BhXIIZ3BJYzolHx4sB+p+p9fiensg89vYKxUtGCGqGACYkiBwpzvwZiEZfFS
w39KpLTg7RSiwa71nTHXbUCc35quUp2azeprFBcLDTy1yJ342KY9H3J0FMIT
s6TONXcRgyEXhNnHQyILyj5q1mKMsUoFg3NokI8INoOVR4X1qLyy+zn5ATmv
R4KPS/scbsCJv8NtBcAf//XYP0nyjQYLBa8PbNjNmOxJsoPaEz+OZpb+XxzL
RdMV9rTCRBG4Cr2Va7NqFeiIifxq9Q70073bvip0ltqtTANDQ3ZOPMqfmrMJ
lVarK0LdBRsQNumqFDcVoksDK5CiUUhk/LGmKmViOK6ooFMmSadIixUVOiv0
x4BZKcnMTwifN/PXifcnMwvXhZj9zzp1rVP1oVpnSxw196hzjRkIOirEYy2g
AIB5YGA7qy356UtbAmbc6aam0W5PlEl3L04TuEhGkj63ng7UUOq0zFsnpIe0
KtfDDFpcEMLm0yjZrv7SjAwZMvlv77LqWyZxqe29RFBlnsD9dehLVtPMvkbY
WUmzjGuwJLc14E4brlILgZHzFKl39ddf7BgS07gRb4nqzm8oIRMdp7ZypZEZ
XHeaT8W8oUPIkHbipJxwcpejuuEUT5TOaC0cpjSAgrx5JQyH9xzUK5x4wUTJ
8EsSorVbWXrh/STUlSe5UQUcT658rT+LxcBlyWv3ewLFHt/sofxJoPXp8Lsd
ZWyjmGETUlUMqEprO8qRqUvNk/U5Eurri5FbrwW0DXJdRM6Nk+yuHB9J7Ivc
Y2gVilbq0x3OQeZPBNmD3kNhcBh8mwDcKhSBmZ05vuCmmwJZvXdJhgyx51q8
RWCnUhiVdOb/CQMmbE0WFlndNPTRxOD498TRVTl+k+WfgTA6WTy0o6CQg1vZ
TIeoWt/nR/xf7kzFdCtOyOvhaOLvNajcy3vDMh1xQB10ko+8ZEmGUvdd9a5z
SveEzoTXHa2MQ9UOu8S3FQN8U+TwItjrCcofUApsqEjuZNW6e0PdOLezV5i5
brJO5M/4E31XtE9BYDvd8kN/OgRLkYpQQG+tdvnRUv0xn/ZBoBNw8JPJcPuD
odohYqQlujqVGERaLU9T82sfWxOttbGcK1x1Gw3GUdgb7jD6zdeB4IHZqBj7
F6RK8ArnarQVQf6xrM8EsAJFolv9DCzj3KtYUaWDLXZk/2+Z8nYNtv4pTUEy
kdkMnNi8+2J0KCaod4PQgD/D69Aq6acTTtzRfTXDhI6zu8R0W4S1q73fw6F6
wgMM+FrBH5JbSinh5yw6/amN9q+4I/dQdf4sCYTuz/rHurTA3KNAEDR/dWaB
lTqaodIBWIyW23OvkRSzkFn92qZVm+dJ5H7N0lo+Vr2XOWqNjfDTHJ306ho3
oeMVqre89XFwfC4DbUVIE/yy56os7jZLdxCFAb4AsuM9LZwKc+vAIHbcEC91
M++kgpa2xo7bzQOTShNx1LDGGFmg/ybTK5Cs1se2yQzSImhie6MBWYLKq4AE
ddyYPu5ESVVNaHctKecZQvur5r3swqe/eTGP0HnxZcFvLoWd9n/urEkurWx4
7wPdLE02pkah5t8LrAZpCaM+/Aw7XsBRrtLFhskQL6ip/udfGCRoeeHDVgDh
b2QJSLALMlCU8M9Aqzd5UJzEC0b6rdfgufBHZGA27dXbEGUEfTBC7KlsQTWL
gk4hzEeLMutun4ugk+/OuJvpROT+yyEJGuNHQf+YcYrx0Ux4byfjAyWp2M8N
OjM96G+6Me77uqOMDYcOtg5Lxp0xvPyqRmAZ1tquaIkWPC5zd4iiw0U3M8J7
h7mdT204Qy7UsJPLRUUoxg9TM16FGKsmVQ8hDCpLTscJt8mzzHAoWtKWyzNK
AcTWMh1gQgnlyDuldBTMye91ePagTMGI1jv6Al4Ii0DpqMMhYrCbtm4MAUWK
X5vQT+6w34ti1WC4+KxxGSCqFYh+lxSFEgry49/t3HvcjPlNt6mbHRU/aOxu
4qSN8gZqIOOPEfQxxYG1LuGRpXwiR9FO3BlINDvpLrNWJ6i8vppb0QsMkoyp
/gpL9wZEusoj1ZAttEY6Khahmrvok1RmDwnuMhUmdY9ZAcsOYZAuajAtax+b
N9MXejaA9UC0/X6P+XL9jeF6Chmtm2d4sECBnpkytcNxkMJO0QJuK+2VaSHb
2gEnXeLtNWiBnSu4lEg3+IENjkXFciCcTrX2T6vfrjugOkqFDQ99l6GdBsUh
4dupxHjFUWB3f9dKU7X43MRIe9ltfsujPl34EwY8cMXHKCu6dJwIOQAPf/st
Dv9LzwDqsV2oGkuPyRQYarsH9bByJZkv7hWef+0rnLbK7yqoeDbE+sbm7co0
G6n9KE+IDyWk/+70C0aRrAUO0jSCRK/IQxdMS5NE8gmI9XYkz6gX+TKwEL1Y
Hzn0RhN1djVnid3xEONX8+IJy7DRAaZLsc4dpJhe/zKw10xAbx5FVXh5pzAt
mLI8DZRvthuq5XBsz9gcRPZGJoDI9qkhR90lAc7AgLhr99EpAvS9Z/3+WMUI
HZmSW1uC9ezMIZSLguZYX6dPdP57pawHUFvrVTqDeNQxsUt7q4llZGk5rNrZ
oygbvlb65Ik3+tYBjUoFooe4rGFeAWRAz5uUlJt/WAUXOv4GaQsiCaqVIdwx
yHHr5eDFBiP3hEC1CAXFwLnge2EW/0D1tTvdz4T+/E5HkWJplCEU+S5X3NQI
onVSkeszJJe1YVamjEtBBFzYBN6+4KzrFBViza1BfuDKZHLsrc7lbFQCJrTr
9Fqy+jT1svx4qsA0RubUT5Qq3BdGIoW8PFdLMdHVq+0jYf89e5EWthMgtG3y
QKcRoij4UOhqNGSL6aKaX5OXmLAQ534ntrHlnL2xV74+srtG0fA79scbddlX
3flpQj1oMt/SBkJALYhONDLYN91L9mCNWysFsBLRgxTzLz6K6BM9EUXZicqO
nG/eCnFrJpUfiwbPrEA3hbSEqBu7uDFTshNjJsOt+K+jRa4s3TnHB6NjhkGA
LdpbGcbm1qkoA/a+HB8lqAKsOrVFes3/AaczVzocLhFAt6r7QXdlm9AWqZ/L
NGDQXc5xxsCcH5xy+vSjYcelZ05LgooZeinzizDg5ON76CiityKaqKP0GhtC
W+m7djfIBdtnzItPjCFl2bgME493sDgvSQd7PC/VfDOUCw3YdzjGlNSxfEOl
9N13cyV5dWETCk3oHnJMTY/sNQq9xjvxPUixee5D1aWNBzkJLaoi8OHH6nnM
S6F9UN9zdqcPW0mQULHRSZK8m8FdzbKs1HSo7FKnzJeEmbsrPvZgnbyeWNmH
4FeCLzdsA9GVYASqBBCT2Qt4nAXCH9ZAt91tQInJqw00iKb8HIjdrgtPDqfm
G8l3j/AO5slN4hBtCzfa5ZDtVZv9gLYD7/bZPmHY54pk7jlg4ZrmSNPe1y7L
+YeapT3HeIAZvvmtOu/qOd01qqhfupQKodykYUAt3ehpn8dCF4vmgz/Ui0rH
vZR9TCs1DgmtiBf1mO1C6XFlmiXUA8KN2G+HEyr+NcG+UJ3XwlT9aKKo1IWS
cRoCAUM/7qbUMv9LHezthsjEY2dw9rL7lHspsKpAPGYoLu/wVPln3Xawf/R5
YO9/c+7mv6N52BRn0ZIt4nJ7870/K7kb66mqG32utefTp1TbISiT5OAP1FER
DMQu8fVeF6AX5zy0WF2WrjcUJTgLjCNo+NWmwPEWfkR4UqBnxMjf0LsCIdgx
onHYgERtWfVjyE44HnUR2gEJmjVlbqJ4iv7TlBnJ2VGFXPEOcLS72rLWVSWR
vX/oPqfTfesS+qGPyMR5JG3DRFH572RKCj5RwXsTQGCU+W0sqJ2vo9y3jZOV
goiIQBo43A9daBNyH29YSZSUpESue5eeJ9h0psQtFgNQH2HvPrhNImsjT2ys
ubmWNyKOqWruGw5HUMOiTNmkkAL+T+ScoMK+1a4RP+Id49zce59a+FpYMKRo
Y1zyjv4ew3Uu5DdwkUqw9eL2pVfO2ceKpVn8sBvR48m5oIK2UUmjuLAlZa0t
p7QgLF3uRpdt9Fg7rmFkNn7FRosrtg9VBfs3o1jTXMF9BHSXOVP4tpYOp5Bm
3NouSRIPWz/i/Ns4uxkg2UibajaqiK0MEemLnnYHQ2ZBkmIzFJWeImPAUHu5
W2g7q05smAIWOEsl9sxERgnYuWhMGuEt8oUgZuxC47HDcpSVQbQxlRNkEozn
bCK/XfrP+Ta0G56AHHuCDnV98Om19ClXpzSJSF1KUA5w1mqX7fKKKICGYtiY
Mm8sJoN2pXH/lgjniPrdvnjO4aYbIH0cQCJS3TTTc9gad8EHh7A5lc0JexbQ
QD4PkjS8ZxJvyRwPS16EEWI9cD4tER6tH7jGrAoOcXZ2o2uce4VcwuGowYlt
FbXA3U+NOeWQQGVdE6nGYhnny2mFpnJB3FR4LguxHZMVgNWXj3LuWvrM0vZ/
vvv1FNawRstfQeZUceRXXIBGC2m/NQ48IXTp47GaJsu8eO72eK5gmwev13tc
N1Q/AKKarQsNMyrMt9rmkbJd++CS3PZmGnhSBv8ntwGeJXcXJYrHfqQlqhsp
oG/EqsIBuT1w/XuXMapYROtGqDOabLtJN6TBnoKab3fC8g//Sn69TGQU2XQP
BCai0eYR78dVn8eLBtBVduLfP1eOg5R8dspaO50gVbgO+2rzOvV7GAytzn+M
dGw5NZgsh4eTasYFpG9n+SQQ75f0jV/EXpZNTAcm87GuuHr9ahUwuRk+w+Pz
QJULXBsenl7I0G2xNskmDlAulrgTiPi/WIDnFYWHghOF1qI0xLO71MfhqdQv
jV6L2to6Nsff8inMoIYkoHsiN9azOYGC0CntisEFXeaezpToeZJUZXGZPmoB
MYXwAwUstiIJTQGHAuJ/HKDPlLG1LIWWfZ2uzc7Yj5EHyrsc3x+fGKzA0wYe
k3MtYFeuU1+O4Ymolfm5799K4SzfOyyukKCVktaKDayDyvSodZDQo0TWVECp
tClKP3FNdzvxThWdDFLM1Sp0ayo0cbx7sgxBMV+DM0xk4NIoTweVCAdxEC6B
3BgcXpFpEylPoUcG8BaK1Ohr3eechGS1jY3q7D6AQhFNGalp2uzWeNnUTI8o
oGYhbi7gsK4UBrbW7Be3rtFpvLQqFq+mz95OBIE7vhe+/tkNzIIj2Xp3y5nz
HaEEUAZiXlI99YJs1pijDTviI5PItgUcv7umT9jX06KvLYjy094xCV2Wb5sT
6N3uoZ/cJZxAsqvbn3THfKPPWpdabUV2+xxeCW79nax5y8VL3L5Yh4aj2XAc
VKkXTzK7ceQ4HVIm2Ut5CsBnB66J05Kas7AYkxX+6B/IdmsI1ytV9Z3hqiC2
xtFNuAA3/dNGdp89J+ioj7KFPwDDPiWbvbXJSySuwkjGde/cSOY4BI7doNYb
LIQ+RDlKBAP9e/koMmuYAQ6idVwujrq5myu/PIPMo/AEaJd2MjtWi9TQZlKT
BLDUSAM4FtDSDcNRljFA0pUvMv2gdRbVIyONZEayTG7vSd1LCLlhGHpWtcn1
6c8uUTQG/9HqccQnxgbdXrrc/6nqKpBFQRIohzMj+O7KCMPk74IYmOkWtblH
/d0SdEMBFiLDKEgaeAke51+Us2uvHGtJd2fx3mntaUCzQAJ5KKRppElj5pfM
yq8Da96YNz5c+joRV7GVSD9C2pfXZ33KUB4f6SYgU7Jbj0xSmOzTj/PKurqZ
BeQXJb9QYvHsK2t72faOIojrAOnxQ6Zi6jkkI7tgMJgBHzA5e3ZFC26P22Dn
xhg7f34RY8HYLzcIjhJksXZTO4IWFyVclHtSC/U0VFCX5OT3yFdxK6nzcSUZ
DugjtHjhXvzNc2z2xM9TTnQ/zHjblo7rQ5fTdfkFYKCPT9l0o/6hY/oD0VuN
3XdPFfY0R9S6PjDn58urh0OF7n3r0Gt/Keikv5gnp1ZNqm4RwXtVByOPE9Yb
Wn8MU6Yw9Zd7sulybWgr/1b3ouSZyRXPX2lIcS+N0catMg8buHGuzyvtzeJI
U/PUC9JTepFXXmhYxx9jeA65sinOzK0j11v7FWHGvzmKJRzvFU2LztPKzk2A
Hv/zSB8xXgkriF1FoJxe9o7K9F0syGIOOQm4rt1Ex5Rmh7fhgUr4dZd/eScI
CHAhJg6x/CRMahYIioO21TFHUC+TIQfDW3iZLlWu+5CrXq7ipTpr6RrDsNFM
36lpyYOwP+LahgoPjcJTAfNEtc0PbNV+R8K82kK9G4roSRGXA2PmWTfIZ3Rx
B1fLpH7W9T0RpmMtGeqF7ObLf1rszsTWsHdtoIeez0QvdBGlc4i78XaEwBbz
tQGXzR/XbZ4gnTjZQakAZMLEAbN2nBOwe5riWc/8zmUfO8TOXcsONFemZsn6
sedt/k/SHQnAnwqznnP2N21yIoDD88wlDCjlO0qGtX7vg/k4mF83hQJDrlR7
utMaEmMkNeRi6oHJ3Yg7rTE+OZNtak/9Vy/qDs6BTiOxoaZY9Ot3UFuaXFYh
dpo6GQneCLljeL1YpKBXqe0hW62WafpjJC+HARKMpeLfcS8moHcu/NSrrXP4
DaTUOl/0530vKvb0ILmcqz6T4tWTPWtHoxl6Bj1vlJHuZZrE3MruRucz/Tsf
9baF+j7v9fVN/+WxYcqYb8ivc5ff2kWo9bDxcmQ/F+8sWAeXuH4boz0n11mb
lLvCg5phgZkDfWHoD1VfZ7iCalKbOQLfIz6X+1fvZ0v+dSgtPgmsZ2ByOWg1
kcaJCOR7N8vraGwVEOhSkpeCr/GvMU7lGKPakZHcgzJZSnuMBBUdHTNQuFMO
LIFyuu+E4QnSnt+W6K3T0J/4gjmd3caWJVpDmy59IouvHdA9+7H+XGToZuse
8rodC1x3JrJ+thnZSeGePIz2ZxknWv8q0GKzRC7I0GSWKTC1+Hw+QJf9D5ID
KE0IOZWDqGBD40HOjqu2IFOAhdD504kx3nqfxM0ONyN79IJdf5ziKqFbvSc9
eLH1OBwaFR0d/bTD9rerb5wLf6py76riO5bYfwdhl/OmiRmJzc58kIIggxfj
KZGL7qfqfvz4TjV04xtTC1XP8FamYNTyuy0uwFshX0SmGWg4vnT9XS0m6WeM
UgrQ8sL1TVeMvTbTXETdB/x6TUC7WmXpY+dvRuzR43LL6r0ws/uf2n5d2m+O
/cxUmAAQSHJ5nHKIqjDMHtRv7dq+faD/cUv2g8DZJFVjPxpT+8ctUGeHjbmM
TBaJnMli3CdJOggBlCC3QSbsEvZZwX3GLdmBpLMV06uU2MSzht2kWol+6rW8
6QYju4pIMmkmCQSvKfNgJSZEAU/7E06dqaYm81ibZgIGRKah7uxeJi14Ti2a
uIo4NDi3JTWm+N/+yVLDTVa1JFOQXkKSZmSawgpYfBREWO8DQwpS4iQLCuzH
L4Ine1O/rupimQEcOIiig0X+kc25UgY1O178K/yXlb4SNcX9lD6l4/6XQHgP
4TgnS2+HfO6vgWZ5wxJfj/mudeFfiwfIvFohNnK8dhyXDU7ZbP9MxiNzHbh0
4jD4Wf475cmjurNpbw6hiURa6xvSsv8ogqASPWm2w+tB5F1i0w3yfqeHTY0W
bCTIWHLirBS2P5hy0Dq1Bq5TB5Ed3oaJMdgTzgadptyaz4Q/HAukm+R6vTjE
+Q6qoznXwgGWErQo8ob1CH/n6HMwEE9NjmRKjFtEqz7Wir96B+dFOlA30Hnb
2kBH8ve1/bLKTwgg5d3gTRJGtsTF6uNOW6rHjerP3fX91+doWIsLvrJUamYW
6E6AKz0gV0AQGLhwYjGAj8Y1U592XZhYlhKi3MevogETuvGnekIqlikcvvoG
ULC/0PgTT+nqted3XuYfBVjoPMs+AcAwpgHgbgBHiQT8MtyJNnarNb1QMBGJ
6ywSQJdezoks7jpwnkEN4LVdGF/fErjyFYcOBOH+cEZTEoLqEq5VEHy1GmzJ
XHBwyJySEPN9X+GOx06OuQCCckbNMH2GCD/1AmOCkbMricJCWb9+xIAQ3nfi
vGDu0sQJvMYO95aUkIJCUTsKNdaG6TntiOi9/s+5HSkNnGkQFHwljs6P1GMl
KRNhCRR9h9MkjvwdyBQG9TezNQeq8fBIY25W5mjeUbjPI/RsRSm+2ExGtoTo
NMxvycjKHPSfiW1R6sOQ/+UoWtoLsfAES/rP4X0xbHa2RtnVM+rbdOls6IGr
muI7TZi1bZbiXNiisG6VNwshWaK3r5qVaA8eFbMd9s0LaUktNC6WUD7CkI0M
6tgW3dmS3Nx01hcPOJ6edttAyxj9xQAht9Em1hoRIWZcB9XdKtZ4osDoQbWm
hhjRjqHxQaC4o9uGhn5iuxrhvt0P1ywVOpDPEGRw1Mo+MqGtO6Pl6jnObSia
1K0rGQeDJmjW1F3glzYbjl4Z/Oi16a3ZHuhLgfEmqE8xJ0HYBZq63EFMW+ZT
tDD33/cl5cFTx1/H9wmM7rCYpGGK29TZsdEhEvGpBtm+jJaNkOtJsHIMfa61
g1Vn4acelWqrjXZa1zxUVHMMaHn3xyPMg4ie9fUoN1L7hLlo8eszTnL0S+fX
jHUc3MHqpPB/Eot+aHRiBanFWwAX2nxkiPEmWa1+1jNC0IolBVkZSS+dTrH4
yLGovBxFPkeXS9z+/tE05JFJoQeyQ3hz9Pxj37xjewBnzo4xVipARXwCg8Ze
2OpGCN34LUgKO5qc0Hk5wqMmyJfUfFoBPVKQEwAda5pYUd4dRdIHvu/Xzcci
NNBCFmJ0Zhb4TGIYEAsaFgR9TNdNZS1+luv5JM2bo5wvhCNr/bJvva9sgtdg
ZVaqAfyryyIVNXKWdqQAOVjM3lOiFw0Ko8smYwfr92g7gza+GDf3oJeV5ibL
pN3hTrm/kyiDwpd36Ay3SqtUFWrgPJpTLj4mYIyBAibnQldy08kGLsnxZEpJ
pSMjRATtAbmUzpfb+CanhRYjHdR1mtUtn6o1nUs3omWbiwNKXaI2xaBiS0sF
o6EbBgzJz0OKF7U3WqGwL6C7voQ37fKa5tXnheJGNGLekKvI9jZJcZVVipWj
wUrZELNi3CNhHl5+3YCuoS1FNhLzZ/lw7UOfzzEdV3MGWc6r9ATF8b56yOOI
Jjw8FCUnq989oCQM00XfTHcKITim5N4WJhq0SJIldbwrDaXUHNa3R4rLwY49
G/YYXqsa4NJvvChJtWm3UoZFUeakw/4G0w//u0Vww3EviICnNWgKomcbHU3T
6OTvRpErmQoPBg7H1fJ5kuPVPi+rtr5w5B4mJ8F3iPuBc8AF8lLvrbolGpb1
ZEHg2Ri7i00aQwiRhKNqM+VapfzDAshipGeUcVONGMJlQrmPOnO/Kf3j2EeF
WKOZJMzLorPnUJAf80sqWqw0HzaDRP+Ctb328S4TI4UJ5oe5sMOyRT9bgwCw
wYTWA2KxknHae+S2Sua0Ua+HzgTuyjjNUqltQAPL1miMLGmNK23XjyvofKbF
FAaCU0jQrv+2wuDBV4Un8F5sLwYBAn1blonxdH9PG9v0+Qf1/qV7zIunNAGY
+v1mwAfrsMVIJkgYE+QeW1wakw+YFlAY3QzbdJQl03ETfyJIv0unthfFWGSC
ihpA2cpqYCXm52U0joNlYEopijEtgFUrfgHeZKaTpJt2P/vKfHHkNO2rHRRK
9kWLv7qBVbybqKimYrh4fzcMiz+cpJwwEp2nTMkjuEDSjbcMwSqVZzClUMPy
etQL/7rVpT8c5BDxGNmNWQ0wBp3oOOz0Y44h1AYgSmcFbSc1v3efp29Oacsj
PBkJkkxN4IdDYof3M3OGaATQ7VdnWzLVcQM33a8sVG5gwEFmG/Cg1cKV0R+u
f3xmykNgwR6IyZkVBSdo7dzvYj/enMSt4NWU+/OMIXLGnX7vDPDcopyg+3s9
5TsZvGq8WfGQC1Kj0ernj6WPFKIqZj8vqCkLvRF7yK6csSKt49iFAyS8LKlX
CFl+tJltfIfrLiSu2R3LCSXkCHp/uCSeEY/zDob86r8fjE4KBYCNxFIBrbvm
m36VCjFZQW3FYc6xl9lJ8e7DH2O+m5GkwIcCIWTUYbK2mFDRhcJXHLCkXRBv
UQKdp/VK/sdsqJTlBDugGYrcg+d7vt+vC23Ak/h7vmdxAebssaBQvrVe4ar4
MV28k79wFT1QB4xiM0g6/wHJM/F6z8am3NAbL2sU2RbvwfT0wMUIpSR776Ww
VCczFOUjXeEq87VSjvR9UkdjZJhpAP4WtwYhZMMS3nQbqzG6eE4G2S7cJote
scXMS6Oxo+lsvbt0iQ8I09RVhFSd3QN5fdjBotcucrcI5rqP2eEKleYPnB9F
273P4/6RD0XR7exZ1JLdSNhe+ZR/BaTVvYEV1zTthM/ju6llAfegTL/QpD36
mMjfXB6mgsUinbIk4CTu/VqBRvexQMdj740FUjRp2w4xg//OZQ69zZ1Fs/3s
J7G0lFmgXAfrs4gGxzRlty9sMWbNgk5fuIgVkBkZM7HMoYFuk/XSxv8B0sMI
T5BL46cppPcRBDIm1vpD72PM27hVLzDKS2MyhcrJvbcC+Ee0TZylCJFLT14l
Op3wBFlI8YkzGkvSNIow2jGjn0AHA4e61hhFs5aSQl4vRD4Vm5oMCbpmMLR4
KGigIpf2d/EW2PnpoqT1HHb4rxRJ+rmrBfLDAX9eUrNxkf2k9OIxPF1f+iIp
a3ZMulq3QU2decolasMxhCTwkgy160bFssAfT+TSV+6Dk1XhtXVLtLl5N/ps
Ki9okj+xR43qnNnvPpoJqU+9YSn6H153lrJ2kO7787I5m44NfUsg6APKatla
lGHnBNy4JLMTkGDNpFkmZU0N3Uhk8HhyCm1htHTY9LaPcUjMOyMULFWdx4+Y
pzORE7Kh2Ac2pX31xjLUfZBOeNlwxu4EqcSDI/XYpaxHz5HXmJSODB4G+Ms6
HkRcCqHPFcWsC/sVndn95DjCacKuyaa9+Ks4B1nHP0Vlpx33ixG7kz8JxAAi
4RkEVgTtZ7Nby2+SIgXvJNB/GLxRj2Dib5XnxfYkY3ghFh8WFyPDg//ygmaE
TiiT2QDejZmWottTEa1XwpN3JSVd8DRHiHpBCvcLWItuPgQbbY0jKDtnl8M/
423fZOl9Vda44EIZsaOU4TRdAetxlEUgJhNQ/k6CValOIjAjvJjcdQD4PSpZ
McYNh2XYWD3zWVg9sve1htmeemml5JM/Vje0ROjwNdo+5cuQosrw18hLSG6e
fphqzPL5zAGjeVB79Jen6svUQ6sYZco9nxo3a9oO9QuuQV4LNFseqPJh1fAd
odu2+sgSOKIotMsjIdytyezK4iq977yJWGKMKQ3nzAhiPdPH9BayBGDZ11LT
LmA0/Nhs+GIDQKCIPwBC4Zcxd6gi6RFbEdC79YJt6rvRd7Wl5N8d5KrpSTxY
DrQ5bcACE1PtaKFzcsOpJqhRWdDkV8cB37/KRHG1My3xzwlEw22MSOaTaSXa
8+kDuKUHcOrdrI8Z40Bpv9eAKJN7HSne0R0LPqjNLP5+50XELiAkAigUswOJ
FqgSbdapIQDzSkItxIv3qvzJN+cv6ik/Sv4GQJcBig/dXPHk0oOSyEsDR7VA
nHG6bN7RduxFlmLZ+tYdIfjXljmlNO8W5qAlhAW8AW1vDOdTi6u+JXzm9Vlq
wFMB4oMtZ9SCL7Pw4d71n9z6KGS6f1djyNc8XpuXsh6DwhMpsYpDbfE3YDar
LZJ0ci8nA9+/niCXGXM/+edkipTZuiLG6UmdSDJyyuCAEmmVXZ0i7yKZtrET
wpQW9WOZS4EsyWhkGK0w6MEgZtk8SuDHiydr4+XMwiNBhkbswZI+mOvJipRx
jaCY+VWb3pxRbUBzKJfTJd5Qc+DRUaOiNS0jyU0knt4WjjrOahPWg/Go5PtE
ZKOkgvgIVrBE1jM5EYE7nJdVEZXVjonlM1DlKj/565uQPrhP3YrMR0jQd5XW
xbAN5qa5F+LaTIlQ8mFPhXQJs0SiUZS4uBXmSB5jflHoOgtWbiSFXYO7haIZ
fu1vjyobz+tXq13vR/3UFZ04ErajTA1ucLe9wqFdah+m9d/nIThxZaIbTv4M
GS0dvnUqaX9rqJ4iemQJHUzfuEF+oYpMY+M4r+x075cnivPn705XkQszePnW
77EXJbuAn0AUeoIjIF4yHPsb3oBKJMvAjCKnNqS6xRprOJSk2V/sKP2cOfcW
DF6vMjcTvAMtKqoCBtnpUZ5iu9WuMAGSmQnEE4Qp+q50rY+3r9l4Vj8Yt1WH
aFe+lG30lgT2PlKhRz5OIUU/cElqGZjKLHw/N+yg1oPitLM+SK8zS6BPHdZx
VcPriLf2pVp9z+G+fmNPRtpaTvHL8UjkTLjL81s8te/inw3xR8Clby+BFhod
9cyo52INdYfMICWWd1N8LMdQz0saz169UQFsJi1CwL3fWz+2uZKWqwSwDyi2
zvurs9bQP3ZAVSxGncxGYI9hX9TUbvvjXbymwmkzucK/YWNqUl+dCvYGxO1a
RVJmEvR20O+jLZ3JkIHXikX4HN1H4PayBkexmQXlFPqhhjGt1ruRTfYmJsXM
666RpvMXeClEyWey8ePaRvTDRGdy/7GzToEVAiBqYGxFcyB3YeB92WNDjtUf
XbeQ2en+Hsf2CvcYPcTb1Xk8/5bRSAxbyGYjxJprk0un5kAzPLkYj2M2r8/w
V1G1DpMJjs9O5t5Qg721L1hOPBRlI8IOd4Xwv5vTEXDwHlRHhFw1XGvO21gv
vkdSXdPn+HUDD0k8jMqWjHKlqz5+YPHgJLDmnqJrxbs/86U4hIhaAcZ6iMxo
x6rJLNN/TuSZiDczK+WZSxuzNf7lFZljTqRWKuNxk/9T7WdUVFKjqlJzb7Xd
JAuGfJBJYeLX4m6OJ1mxRDD4BTsdNPv2CrMXhu/QoYa+yS+AevDTFZfDY2p1
1LGC7Mt4wx6SYS1NfN0heqygLel/6AB0x7MtqO40WvWwX+cuEGyktWIxr22D
kfmgKrsEt3I1buuNWWxyX4ky1ykoJZdpHQmqm+qOVgN39dH27kIZMYBpvyl8
73usv69jjujCk9bOcB5gLpZw2JFJlowjWg/3tnITcwnn/jCY4SgVbiY2OfYo
0pbgTVPwFtNm6g98+qHbOvXzlHi+Wu4fEAa51Kbt/U/elZLna7HQqWHju6Tb
B8gfBxARche3RpOj+tgUpF6R8pafz8p/ZOVJezwZuf8HkBqX+vdSrY1JeEqa
0n9UWt5hGO88KXEYyay3jrO+U7L3YwNFHDSMA8bAh3MO1zSKHtDSyKTmWzDC
Mngm79GcuHSaxOwDFNrQxM56aAaTWRlyN87Qdv9h5Rhv99d9qzGu+PPTLF1t
9WWY7u+bSfbwrizOm6vQ56T1e5K76EA4M8l4cgWUGRxaXJy0mvjtbp6McsXL
wNJUEx/mRSt/brJbo/K8DLrA87ZCDobXkOyv2kfsQQqBtvaW2HZ8yw9kBImj
E1M7lLBQJCEIL3EBf3Hd/G/Mh/bvYSKDqh3X04maGkDwRT6MzQ5XIRF1Gk6q
flgKn9XJ3UfPt7rxpmIykYroUrCbrb7DHPRst2fy4X+G8VTCApRawnAxyNYU
zdACfdLf8+1JuzST5cgcXcNaqOEzFnXTKZVgm62nzDG9xzosQkqZbm+VSn6C
b96FB915Pnnw0BSrlJmcbeuvC9oTAd69nKawMFN66tFGYNSEqOLE+G1xKd1R
yP+vVU/+L5y/sMn5xP+hzEUjblCf1ftoGIkF8T2nDA7IllYlb0crCFKWDfi1
WSjUEzg/2XeS6Fmb+keErHbk8qn3bxRF9llp4KQ2kgNDmn6FxaqO73Quc/Cz
912i/rkUyOaBhWDlXE1djkzmZtZpGKfdXu9uHxrPeBrKm9gazOEu0OMDiKpD
1O6/+vqdRHX3cbmP2j6n/kSuxTvL3Q2X+bXpMmDpOfFzdIbulTW8hFyj5Ljp
UpfP5B+G3XZcBTS2+4UmUjKqnF8Kk60wO0G5N/YR66hXvkuRLiMAuz8vmtIG
WQe/Yo//UN6hfWugYrsNi0sBbe96poSmQ+SwuR2JI4bEWqqU3I+veXTaKT3h
c3PUPI1ltCKvrJIeFKUwh/tJI082jeeqZTUP9NVws8cf+qKMcd7WzvtI6xv+
GthWB4jyXxkCvjxDO1wX+3BTQwLPU10csp7382DrQVnLWNObe8Gma1TC/v9Z
t6sPZM3TjClymOCKJ9cjyl7dUDI0rGUaAGbutkgxrgFsQ1v7FWqUelrIB8o8
YSArHXSE+gjQiDE9OiiUI/MJeLc76+HAvQBIlaaQyZAmeFMrCNDsxzoKxfwH
560ZUd3cpj0mDsfBEwKpWfzPbQYKpHXwHpyjzONq23z5ywCpsw3daiWYBZzO
uBgHrO+A8mE+cDkg5cdSTgD8/tYVysiT7qc13vrTP52Fso8myk+FLe83KepH
e9nfysRytLwTUxf/HpPRpR6C12wj12xtRKUQ37X7EQtTBykoW2vgN2Lw8ku0
qb0j//bYAZwLcXEWIhzF3agiaO3UF+/EfXoIJLC2EYT1JlKViCSgyn3z25FW
YwWU4BQwFHvPbfvC/HqOqhiRTFIf3qR0APP/KoKW7+rORqYwT58CdQSwbzd0
MFgcqtYIfEgrAzirQlq1gztHvD+EPLNVxiUT8Itmv5Uw1H8n74+FepBh0S8i
sfAYFN4+Oc+zzF3CKVvWIvAB0SX7VVE8FHjz/r3FiHJQpOTYZbY0Y4XoEuy1
bPMrAvl5U48tiIEz7UEMxvw9FOsmIFROX5cXuLFmoq9DJhzkFaKSDMUeVwQ+
U1JVcXGTdnl9GHJBxBNG2YrAUmwZzgIIHkxnkfkC1djRxZjqicFObZwhMjEK
z7keIInUvB0wn5/xxY1ycA4qKjvJ3YwrCbPfCd+J9hZhX+8klM6hNR285Lep
vMD74bM5FJ3cbhwCI0LmduCSHvWzg8tuID2hcAq2jHjViSoeXBqghByQssXE
0GwRIcVTWRA8f3VutyINEqG4wWkmcFv174lzOPIo70saHeXXH1bqfmU4KYMN
JmPoMMQtO7jSanSg9NLGYBE6cLwgZp0dA0CP6vtbOSN2TzdPiPAAj1ajzF3Y
kSsa4LZOww9FwNMYf9dkHQo/pppH6clOr+uvpzAN+VpwaT9Za+4Uidpdro3W
u4P4tWoo++a0thisNiKAqxi699kAcXShTcbIat2AWlFXgkw30P5DoFPWTk8c
6QB2AQoZ7TpV2YfmXlv54zowFmy9W3dFN90TIBqtiWGEbkoA7Sa4V9c409y5
i2dfgBrPabwJyMQnDz3ZP9G85ZW0yBEmK4LdtUUMfIrl+BaHQhQqDnCFi7Qm
Z4QCJcEAa+4b6pvpuShlYLwXV3SW0TjdTlJsT45DUzggOMvrbYCgmzjakDDd
A2P6toCq9Da6KfkEzUGCwhGTW9krysruPz3n9QDcaI/txWF7gTOY9ePhxe5e
56eHBCmtK7RZpEgUsWwl+ooPX/5obZjoJzdpBlodHzC6i7pUMbp8cP6ARDM5
e/+ovHGGWZHMIXmsJogCczhu9gggJYOAo+MQpTaOkPYzj99IcK7DVWPzLMj5
sbrkbdVyguqz26SMSntEEDDCaYVwHMe93nsT8S7iPdNIeMvmYCL26oGB7lgZ
PiDQPqkPzL63TeEOJLSam+4QMQRu9yc3qNSkyEKbBx48krFUwozORNg1sI+R
zsOoeXX34agiktk9Un94YWIF4c3SqNnKHSDHiUK0Lajx5SDSRBEGRM1WRfKH
qpBZWPJlypRWr4xVfnapvcrjeGRJjDvcdFSlcnY1pVl92aA33qMd/przWJt+
g/N40sCLB0aG3Y6mm0MZeEr08fA1mdObML0HhFBDMhGGSB21WNhcLBoQTW7c
gnx0ifHhVHq30JwPx8Gwve7sxZw1f3LisULK7JeDmeSOxChka8QH9VmaYGrm
L/77iZEplpq/8MlcV2C67i6RVnszZnxDksgt9ihxR7RK6Rjw9vWRnSaJuGWj
yxKVISNACGdxSRbKE83vtlD8DwPbS4Z1Cxl29rtYptMMKFhJqcas7beGL9+C
SXmeVWSTMiEV40xPI1mONK585PKKf456oX/pcYL4Pe2zshEb6Xj5BpCfZ43N
p2Hxc/9x0zQozIFYokm/l9okqr9c8AfXy5SWJRBRfAog05r0uUkJPtsKPiYO
qVmn8BVB1fFGxfaaLgzk7RP7EQ+GdSHZx3mWlVHyO9GlDdDUrVLF558HTYcB
r/zc17V5G1oNg1R0R+9JkUZkVAfXejXcayC0l8o1HC6Vn1FRpXwESYTh0mji
a1d14I1zGmZZXaQcVx/jnwNmllypea67Jid8W1vGKpQUgvpVLk9dMOGfACqF
0OOxV11ddLSHEKkfDB2i/jbySZJN1A6NFH5rdWwrHmX++mFrV9AiDvF1UZUT
Tcxn1+Vu7hOpF957GagfGhLJd+UxUQMTLodpXAcd8po0qKuaNWPMsuAR3wbW
jtLU8RvvGV3410JEllKNKI2SOodOf1LodklY93teocsPbY6FmFwkIvQkWl2C
zCOJDtO7/lwYfbYKUpxYJmcfrU9MN620YGEfQZe8blvqHo2cNjgi134nYmJy
EfGjB2VYSWvpYsaTZENC5H/lcXpUOkZcmcBvr94+pJoxr7tWvHXHjFtJ0PI9
+9+4CAd4OiCb412sYiyEBA6x1012VqZMqJSg7DjwLHhtsHS1RA0unN0Ze6vl
GZZY9Inv5Q2ePogd8k9bjJGYE7KcoIo4nyXG4bepX3fFeJWeKrgA3gPDNPtE
OPch+F9V5uV7DTjLPCyXGmCN0R+rqWPbYKUPghqxuTI1iLlSFWpLx/HNGT2n
ZewChEQuLsDz3WjVHGB75I1HsZOHppYMKSo/Jtpj0szlF0/iksq4dv6/Lt/f
nogQRw+EJ7Col9PWIfjRUtbRRU/mQEzk1QwGhWwejMd9bUVG23EX2WaHAzER
M4nPwepAiLyEmLuB3s6q9oFlcaZWroag8TdjaQhsOuE8eRQ+8V2O+fgjSW+N
KBW/isDcPyTfdJ0m2OqsxtgYNNdPVfIxAEWxqcVeStlzFk+sAWkSB81nq9no
2RjGAXF9eI1XXBU2UuxRLfJA+a0J4r2YcUm+JsPpFxgPMaPrJeUGD/aM4Ywm
5LJBapXAuNXwlqdSs+FZ0YfxLs1OFa84Ndz7GyA7SquqSUpZvG+DXzqcxb+v
9YEYg/DRv+I+Y0fVCtNklm3KIfiQHgBX70qw9d8HauKt830epnYVlU9Xx8eV
Qgrt+6OxSPxyfJC9uTybTOu+DzAWYtsJRKosVRIkMDlJSanyW8ryOll0ZoSc
wZEY7uh+Ue7ay3vFohFs/LR18ZKAopybDwE2MiJyv/azg7c6SwLsJkYuPJpS
vG8Aoj+xO+Xgi/fl4wm5HZxQSC1/O4K+K1khKHU4lJb0EZko8OxBXS2RTEdX
Kg6FrKOZEAr2y0cfgs/1LbRMa+bnFWDlZria5/GnoyyVT5IgAUXjH/ySKTMw
c9WQRkKab8SSX31StEqxVAdwUL95i1PFsJ2+plVraZpZudoGkoiWp++Klk1a
iC2EguMxmtM4wvZgVFt4uhfMLtp5SO+zrwGNVCUSlwxWNbstyHGPTNHz7Tcv
msc77W97SKHK58hyLo608ZazAKDJwjlnzOd/N5JSA+HFm1DzvwiZskx+RNcE
Qw3iEqsHTm5SZc6zzCsu4zFa+cr1TJXwb0WOwUb1UK4aRjZASb4+AILQTg5b
YtPSD+4bdTWDxFyZs5jpea2ZfcVzHKDZUNRGMnGpxL6B30H0mHluif4n0Fbr
g1vXMtqvsIE3DC8vzvqy4994AM3U+I+bJmPc6N3nX3xNz4ESShjX/rLBePks
O6aEfH+PJRlCHX4YyN3Cp1nB7jeTlmcDEFfWH1ixVYflCNfasMoUbELgjU1B
NbawYgH2Xg0X8Wg4+wuKA0Fx/2GBi4+gRCXew9pQ8XepcOTqdE3f1SVCdbXn
uOk7A5ALDPs8sczdaWa5yEA3I5FunlKEYZCyKjJtK9fvAP1ouFpXr77KCNkV
ePA9uc6mr8g/tfrjS4EPXl3MpKmqLkqeaJ/HJeGDZudLy4qExqxzQhKby9at
2UhbcikG3vAuphP8iMmjybrl5OoP9d0c/ttcNWCqfH4DfAXIfsM26mX/hdNS
7YCa6/E/tKRfya6/VRlEP2nW9Qr9ItVCAJc8JlnHwd3qDyfKZ5Y/q4l6FgNQ
pREBd9nm+f5AEvdCLd8TzOiyLE6tzlajL+fhksOC7mVwAsnihAVg6jawDPY8
2L3ZE+UmDo6w1lDVH/e20PMOeEtge3eQPdowiEQcg88H718MEXNdwscKtMjj
1cZivZa+dnchxWS/FHBzozCL4VlP8yy6T4PTnhAUCVJN+aeNJHmfyjBh3TMm
np1LUgyktGVHUw7ylOtFSwK/43o5ejbP8xTxPQTBF3ntrjONsjGu1rTT5yRr
gSF6SNvcIamEAcKNsfr176fC5XBD7r4WgDXNtvCkOGhpMuRFwspcbENaOziO
LJ+73sQ5z/TGrNIm04ML57Cm5vIZKGglyn0pG5iKkbLqCeeOj7WYGw2CRzen
0MzYGoANqzl/MnvUBPTZSIpIZbYafE6OM8maPW5lOVEuDk9fN1bZrAiFNacc
M80U2iS7Ee5hGDxREKcYLr2nYcdKx4FcWAY2TjmfdQvMuSjbpsSyEloPMNPG
FGhZBTjebbYnhif/YEURzrWwXLDrhpfL0b2aS8pTnV6I7T8LN4zlR7vcHqkL
4wgzv9s2+r7Cjf3f1RRpVaEjR0s3K2GTOKsx9bFXPRbe2WuWSCjUHhpQfEB4
N5tqVDxzKW9qsBxtcuXUFKjsUZfN8ClOD5/M725UksnmgNUENilcrLLZEg+r
JS/somVzi4OICYSdna7WQMTL27Lr9FDeLWjQqrOgUzUIHiarBOMe1xxgziow
s9NQWZyXM5skwt+WahXekjdI2KY54K4nQLPUUktdFkdeXKI0STIt2QFOJMPV
01zUrYcJCzPDM1i2zGj6cTWXVvhfindy+r9UyoYIEbaw6z5lp3+sqcsjGiQj
o8sXTpeODSJUozbE65nmspbKYUF8cSIH12KvGHlf6JjkgM0z59V9OeCzfI9s
SIFyN3fVw0dZ6U2sr/4dMVUdcPxW1N1DXZrPwYQfn1YQ2wZGDfDvCtifW+yT
W8VKCNUu4kbk7sQqx+vNVWr8IlHYvOFtq3mDR6uKxyfMtZQTFExlx5hstaeP
EY9SU5CFRODXisUbBzpHP8GxABLTVFHz8pJN/+xuk1r5bBidT7eeEE+9MmF6
yoVsMBu5UisRBkgyE60p6AAO+/ZMZtTg7t1+8qzSlQlbcqzVW17otJJC/HtX
IznPuu6etCpxPo/uvm/Zev0kHINkjFjyAKDhJHr0v/CT9RCZBmrI4jF42Scr
enUVqfMT6v8rixhIRRkE9xzng6CGuGa4z4K+6sJjQnNI36cjPr8HmYo8vwW1
1v60sq/C1mtAmwa6bUbZ8tdi8EHXxp8gi8w1uNSTtNR7w0SwAi/t7G5wbEaC
OdcdPhB4Xq+i3SXXxHh0Ipab8cothLQexthOd4PWsQRxpJhp/IghcnWRGLJd
JOg0VabZ8YtZVNQoAcswHGNFdo3dG3Zl2s+gXhlOSgETatAiGgWCXOtztzQI
8DmpIFAyzc+CqnS8aZorG2ma4BKCImZKQuOvoJtlCxoK3byGsE7zCVEeHKeb
wJW2Y0nSC0WbPWXBbZaYg4bKWvMb+SQrZ5ZOZlRu6fM5VD9I0ltcKlls7Ei+
q2SVAZI0H7Y5fl0AgH1J+z8eyrTMwdESVPbdySYOlr4t0Wwl4KLEjWvBqinT
VncRrKaY8OInKzfOil4lE5tPKpJvpkhxjakajGQ3mGSG/47otDtVKIQcF4lD
ItJUs+sT71I0RnHivQKITGIBgmGa1CClQEi46ZJ1hSdJynb3V8j/c5NC24Yh
ZFcBJzLOvwWUbT6KRoQlpXO3ywIsL0kGAGjeu7KvCkI9eSqgy7DMQWWP+Axd
HOyLeYlorMhey42WuOrU+BZhqmXNCMQF7/AJ0/h3VeT88NtmFapJe+UTfd+j
mMI69MrsqmGtOovJAnVPAJ14YjIJNKMYJDClhWnIlGyt2rcMpc65mc5LXJVF
61fqLARcaomoPFU7/K3R6+0i/aoz2BSDM2QRiY1139jASofkpnTnBB+JYobj
fVpPz4Wg/Da7bKUonhthZ1LGH20BheskSsckHidu1gEZuIaCsg6bPX8xczdj
Mei9KPGduu3AW5EMKEV5a25rWeDAKP5kn2FaU/8N5gYpH/uU5W7wf2SomK58
pqgjKBTEVT13kPPMhkqAKt2Wxs8ABnKEyr1zXS0uUO/TUTXHpKFb1RmmwLOz
vE66tqgYLL3sciLr4pOtO+ub/IX9fToz5rBWiOOMWd3Pb3YmSt1sbf80xOZh
j+kszxElFWulH2R+H56ZYez76ABhOEjg/BHelzZagm6WowY+E4xOYbk11yuk
As7iOG/FRj+dmsWQG8QuMrd/K8oh6YWbSDCx/FMmg/F7V+wdP7B9IdJogaIX
ZsWYjvDiqK8Zjq7nU9bqPXgciCXl9g0HjkJO0S9DNzLbQl8Ekr8Rvw1YZxoB
JFXSfmRJSTxSps2TW93sITdvOvkAMC+n5RvmMxupvppxJ5h4utfNnYBoHNOM
pze8fwqBoWZy2o0AHCjn3KH3AtzVd4qM7sutyhLTdaCQdG3ZRsldMswexRiP
wGV4RBFF6UPJF+Iz/xk1vGDPoWFsHatz5DtwkkhRC8fkzzdExcrumRFtn7R9
ge51SzEjKARLSeCuINUw/slTLTS1tqfMgm4LLYmGk7CfTd7T4Y1pZmvHPzrH
gL3lAahzrUgq58WE/duuoBOX2dzNJJXRuszo32eN1nkafK8+RrojnAp9J0zL
BeoS6jaFO/TaeF0WXO9j9fJemLyLju3PkZolW9S1Va0mkRI0WThvnKsTcaGo
HQ7AodEHn3CB/Pzd/ivJMUp15Uab2Fw8KJhZhA/LXV7Fx7+80wzfs0+eUo3J
oiDkmfBmRrif/aV2XtVxi3bGfszFlFE0O/0sUzgMCeCOfLyIZH5mrZM0wO8j
W8VkYc5DZYR9LC1juLgc4zExmHwDsXJbf9cIlQKt1R7e8V37fgSLq6kleQff
1qssvbWmqLCr7i49oFi1fo5+NewEgIF5X1leKEL2zvnQwG8o4U+hHIH3Mjib
7w/c3ipQ97QzwIjeXIIHHk6wS8ow7fKpGoIArw7vZJRNUHsRKGARfgROzLON
AD5B86xQ5Nk0yCp7EYAI5RUenyhEAHInLHhPUyIRPl4Cm7HSTfp9HF472cVG
AisqKVGPQPMumD+zODC3fuCiba6rUrMnoCdR9aJv2oHLZzkw5y3GGFdVX0ke
+FMwtsZTL50EQhOjuY821n/lpWetXJ8XaUscaWEetnoThUY0YzxSC9GBnzcD
4m+lytj+q+Z1dDZ9EiYNaOqz6623qIiDgWVKyYwdMcacjo3eEnTtakSAAN8V
yssZwQRv/BreksxL5eNhs2E0Uozhk8abjryabIpxuYsRa+pkoT0yw7z4X2Pg
xjLqtMrQ2KCel48N6Oqu6wMLwuHKBDOxzX90LWqzNmcIpGRV/rQXkq5V1lps
Ggs65Njw5qCff14VfCWtIU6lvOJgcSDxac6hrA6ddId8CuzJYVtbdQ6mkZOB
C8gPO5fP6+qwrSFMpIuIk8OaN1P5n8T3KNLnZQmHiCQM+rLXiRngTL2DyZ6d
3WOAqfMA1bivPDM84P+YcwQIZa8i0w0g4zgnCxNctYDcpQJ368RNuszuXH/c
xkJvAkmjBNN98PRY8JhA9romEeQNQgyksKYhdvs9cgk5puCfZQWA0DwMK3im
K/7XHlLN3V6WgiuBLH9ysNDGRKmUyytJVMfFDIdNdmY/O2Vamr8VD//2nUvB
VN4/KSlwI3Clh1cplr9LPAZEb8T0Njyrll0cgWnU96RqpsNZajkDj9gsVMcA
tArqSoepw8RNMTKjcaTvPlM36ze+VeXM604a9V75M06nP71PWW/ejiNpqvvF
balnaT8QrB5mvQlUSoacRENCYGb8Mha4yL6SILnYh5Yk/f00or/8C+CtU4Px
+dDXdI46i6dDBCFv2elm0tdpLWvJSkMbpqza1Z+RVpFXHQLqhhEoikzVNBQC
9xTXIU0DsKpAPwqjIMk3FEHWu7OGU/3mPxjaxOy0bxsJYjGLFal4mBoz/z2V
U/BA6Va6BZVJeIvdfAwY6IZmZKhIdvNU9YoRzDDTN49m9Fbt/kslfLzo3Dm5
ARouogM72NVyXf+CgybTLatSTaY51dTZkrlI88unFlK1HEmSUZnfziTtn9SN
3uncNYV/GMv9U1EYeAEyGtEtzU+0QJn81CKoIWlrVhGLfofUo4Mq7k33oUkc
G0JjJMRDGN1Mu0T0R6q0qHKFwpTcL4ou0u1SBHQxDotjqfl1gbxFOwFEvDZl
thoZbeAEZ5djepuj5+GpPD/IKgxXq5y4/JKaT4W3L8ygknxkLOEi72gQrB1i
qESoGfkdFmTf2Xtjs2O9btV17R42EJi1ky+YBp6wKbu0gpJkmf1Ou1y86rgI
lCpQ13KpWrryPwIs2SK1YmI9Ju494Cn4fZdqWmfOwoxBPTvLPwCcSapO9ATJ
ZVWugP7rbTWYy9vgdxgnalRoozOdK5WH+/9EjfMHOFJ28KRFHYeP70+8GGHv
MZEzuCtAtGt2JxduElG35/4arjUuCeMkZLdegpU6ytN/4RDdcGaG5Ci9Az6e
fqDxliweDCk4UAvr7O4WYUW4kkyGwv2OwEnXPeP2MpXBqsXyo47C59dYaain
fzdhPqI1loH6RGI/UVm50WRqLvWcqI5lMe+fQdER8NKGdKQcIDdu2HtUu/Kn
Zik3OTw5WKwroPw7YGdYwzr4/OBVHphdcc/Gf+BKexqlJ3Yujxl4s/TV2YXa
PkcuDvf3Lz0hh1logrOviXsRNv94+9EuySINFXi4HjmPsBBXe4oG69f9eI21
IC3LRGr3LQXkcUkRSY176qbug8OPteNPMpUp3ee2nQI+Xb6mEFg0RrhtsZdS
kQA91jLQuCMj3Ie8bBbW9tXuTlNQms0qtfV7a4gNyqWHZfKc8bJ5ymLLGekO
+LUj+4jGm/PQgfqLitt2p/14z8jgi/jRpsgBbcze5f69YExDfeqaoiGVjW3L
UuPJCrO4eQggm8uBPU3Te9Sk1jKytvoMt6WkO1V2zJzmlVyYaNbVaUuCtIe0
7n6DEqvpJQ3BM8tW/Ai/FxSQm2hDLlYo8TvRcGlH/W5NGcwLYX+PGe5K4wd0
H710Oh57XhNOjToTBAIVkb/fb20TxveF67v/qd8X5TsUkOiv72maosnzpjkp
1BW0jMuCp4gjXV77KpIH/KpoIvlEGEx2QufSzBKI+gvHEGf7Zd63PxHbNqES
MKLh2Bq6eRCGF4kpDh+ZE8Wc/L2Few+5XVoJxyxoLXF81SqDDgmBfdewHfOo
nggW7cOApcnu9nWpAQTphODYkmCDzrAloCc0JaZQkDRDgTOgeF1RrayAWFiw
KlL/ub3SC6ERSNob8AkIcbUCqhkU8of64RFOqnWtU8aHj2ahF15JVP+zMbig
lxiCSNXEY7bQsfvbfrNvMcfFx0sRa8frMBTWf3+HpMpS4pBr+ffgegpb+yAW
N2y3xDcfVUPDjoBv3qwF2I6MUgQbaILwwDhVgtjzib96c83/lulj0LV1MKUV
o//qvaZnmsUThhmpTYlmBVKoGMIfpeSVrR6p+zXkgRbu4s1EwLllUt7d1CuY
epYfY2cmaZLuX3+X/sJK/4GKhVL8S2HyqXMqe70x8kXaorCNXQ861xKGYRCx
sQaA9SEnzL7NpizV6FtymDKfib3AjKRDvREsOUrdVy8K4IMf2zNerm56eRmA
EXwssaRFIFmLML6G/xVbJNdEC1oHh/xk0ztCpMkww+kbXA4JFLdjL+CT9sJz
tZTNpFT9CjaOZxLlqMeRUvupcE60bMMCQck3/S3dz4BRpfsFrO6phSUeMM1a
TU9/ubbGZAR0DVAk6pMLwTw0vVETZL3N6gLZbxBGi2/v8SDa2lqgEBQy1G2U
G/hNLO/uB9l2bfrSJPlPn9uYIEaNRtTQcoGJG3wkFXo1wVHZs8+IEiyyiXfl
zZGspyOZA86lOM5VkjMX2Q2ceudu1kBYbedMNw5dTsrKvXZnpUPhiKujfnGP
E5//tYRKcGBsQsYEYJNswMj5bcKTcHmWoJfgMQhCu1mUuXxz8nvzkK7AJ8hG
9m4vefeiZdLMj/L0yvlKDHyrfc3PpJjSQ1fmKpg24bHcfG4YntsKnFu24JYr
XWOwmBA9AIIR624aYlOQHhK3P8Xnopz8zABuwlFgBRfX4MqmKsN6QDQrnsvq
r9EZLDhjtnocbwu7dG5Rb7NLT+OZ6ol47v0ALNCASl/DdeLam4YExlkBCSJE
WVuGmtqrHsFK7Ji0G98mbdSWyPPMfLXToNtJ0TQvRLGZvhyVfYjEwzC9L2hO
0DnRsoi02jkccbfhSZc1VYo9+hy4RJWyiPpnAcQfVRuhQZo0UBgc+lltUbez
+1wT944CDPJDIus+L0CsQNMGCwAXHHdfH9l95CUthXOohukwejCp0zErxNeI
1ChGpB/eh3cFsknQ0R5b3/lji90PW9hdqG4LVvTxmFgR7ORTSvIfQ5vJvRP1
DyJwZz1jeYrcyGI6FnXwjOnpFL6t0GTb+EtnT/GAT/5Oywsl58JMODgEj/w4
187svL70ZQtU/BOFtHUe8DWhYoPyXyo3o93F7GigaaAJNpFeXmUOl/xuOSci
y8SaksQfamzTZtPqZN+dOfjd1/i8jZlCIIcP+ox3f587px79u+HKn8ue0M6F
MeQw4hgZOIaDrGUqQPrSbS2Vrpc5qCFtws7xE3ci+Tr6JXnb+gNXFoHFqY0S
6ioYk76WRdNe+mQOX5EySCZ9+xTV+mlkmPwxWQYGv+N3vbzqXGXJBqYeU/AS
NMjWnMba5TNeIDpwaE+2ZTqtNfJatucwWCQYHCsQJ+JfyCeStkZKFEjHR7ue
mJ8w5hC42lOpU5qPmxu7j0u4KlwCAPRm+e1uY3f+Rp9UbKPa1mF+qXHVw/ML
FrUShMEEBMuKXLaVatLigFTWus+foFtxu5PexpK3JPWCuV3WVD8FjUuKJfaQ
vyolMnKBNjG/pf+GDxisJcF7xifF+pjpXEtAInNv0bNFnbLTxTJhmfznc2BT
mMckLkJiOIyTWelGe50O9CbeKhApGSZ6JcNYpiJu9ERz3TGnwSQTn8Zyib3J
1crljZDuGTwGEak3OVliAlddbQfX86G7BMZ9qOYvA+/9izXsCbqCCrO4yhcK
XW/RAFmC4b/QEN1pjvf/Ndn6yshcFzL44s+SN5SH8RkEiY8jIbvrYxwc7xT8
7hFUTYLNqaR19gZvEteBRTh2lG/zJ4R0oA3sksGJhEVZQGzGeF/RtdwB/aek
pheRZwCvBnNpelmNUEtqJpzCw4NKBIU8jrJWof/9/8QcTJ9eZgJBuZ8ErMB8
y0j8Mw+dyx5GnswyKdRhK1IkSyg9COup48T9vDJDyVvTsOlrjpTCZjvdQ3zi
4inBI8aiMKYgrNDWWhqGMNlVHZyZmExkoZI0qo3qBU4WvFfFpC+Zp9WVcsNH
6jh3eEKEcx93YCtoZ8lnv45uYTtPKss5gfekEuOq5jWhPvN6m+KpMsIkho/8
IOYu7EQxYUbLZ1oiy/B0CuziAOfiVFQgpgzE8eZw9rs/UCqszoLa4gCYnk2h
RpaTBCTTUH5T53tpUXjT6TYkpxE4us2V1AAh9eXKyYSew9vBBJFLvhc9/ErI
IPdcrWPNRtSic7RdyNNDb2JpCI7DnUmDZ3Vv6lTyrQ1q1yvrZjbcMZz5/w7q
pFIAk7FvIlffPtxe7LYNr1wgBbcyjgeCU8BUsVZGr7bbQx48ZyP0nwcyyaVj
bsLDc60curq9AlJ9hkbNJp8iifgseSw8RloEwYcq42Mvm7Baj8r+Qbp/ueBb
7oTg2jzQJ6V3E6lA5fD25ft3rpomXApVxaHsM0VofhMINYbqiEasbssB6Xzg
COdZ8DTOC36PNBwYbORl48JtXLqDHUqUVk0S+Xu9yvvXLnVrmTruJh3cnOV9
ftgUxrLP8wa/pEsVLS4+X/MfPDDtCmA/1BB/ft1ZrYqR7GmTZkx7YlBFiIgr
osDNChl9PXDoMjUdZmkK/DCU80T/nvKTM5Ai1JqP+2ThPmHkFE9n7lIRyeq4
ZMOgYPU6Awh+56hNeSHJXjrdmu6D5jV/ek1GPCMw039Cp7CNvpdW2+93chTj
eNFM/WJ2+GvAx/fAyqp1B7olvTIGsPP2798KjSYiEv3BgSNFZT1ZIkmP6/+y
g17CPZ1OYjHb8YSScwUMggofdMezZqRQ34toICun6wlqZEyxH9P9q2vgSYMX
alfIE8xDMFZxJXTKpMgHua6jcLirVSbRXx4YEvlW8nJjNr2bKiroy8Z80K8Z
2+utamraPpuDUwkDTfplUO2lFy/+kbiqZCLwjcz0YQvf0DplPjdglL+ynS2s
OfVMeo+cnBqymj+7iAPRQMkTMa+g/AtfAvK4hl4K3dw/qRC+W8K0sfMjojXr
a90uj8LtqEMumm+b/Wq5hqgasI3cSymmR1RVQqbb8sYwflytyKpYfd/MBsbb
vdSx7V/qRP7rSMv6QhoRnR4IGWJFicA8xS5fHBGJ3Ihb2VaPP7OG9LhvGmpB
71d9309KFzy9XLR5dhFNJEz2/lj3ITGyUl9WiRhiNQB/uD+VThJW/5eXGsvC
YKeBjdx9Lpu+qxp3AiW0n049f0BGjr6IO0tMVPoYe7zcl+OWrK/LRAkaTFpA
Se2s/78bZLe+RD/WYfgcJRxoTq/jnAXATGOF3YXrCXhAF58BIGf4doe8u7j6
H2yog9VAk6cJ6kwPt2d63Puu0uoBoFR4+OusSE5muWzs1nZQtlSQhfrX+Fom
y4g3Y5sjIjs397Br19LJttct9iXJHLV5az4OcT+GRVnjBXlm5iuQHMxOhwCj
FNN1dxx/qdsLmQOPSQ5NuBihPINPfNvu6XlJ/oRBAwcKb6Pj5WenahRTIYIO
rl1aHqQYanCvOo4hcbg1Wmb0B+jPOJD7T8W/ldh3y0OOavbUWdVP5DZqCRGM
AmQ9WtdRDafILheQDN3M1LKI816f5D/wTnWZZm+2Qt+p7TRjWz8olGIDsPQt
AyWoSlcVxVHJDZLZKuZXa1prC2twirwDib8Z7QJ6clF68EDq2xyuNItVJfqM
SMkri+ZaULkDbYP4+MShvslK/p9pptPP8UWC4ex0xss42KuxvqqFDvgpGDw3
+cKpUwrj9G1EIdmLNzTFf4ln0/V5EIcHacLuksgm0xeDAc2XBEdkaXneV84e
WMotrEejLjMmL9Lib9bdG/55vYZhne9JhV21kVSkF/IPnCfxuT2nY19K+Htz
3SUzX02qZEmmidyi8Gab/ajgXNtgJNjc5KZdx7M7goCpWyyTDbFOrEqBV+Sa
OrFdDpS4svB9C5j+M92ybIsNmAe1Z9X16ElK1C05k0v0gZLh1MwYu7nF5faj
TDpnBM9OUvnkhLxNMMXxxnW1vZixj806L6Q08Vs0P0NjHSooIyYzemO6os0R
5MIeqhizS8TNlQwSQfiGvzLHzbtw5B4Gim26WnHkDvl2J6zMzzdnw48CPuUI
kIbSAP+MyEn6fStmYNXf3lzxoWayoFrTLPXlPEXA5hl1RsTo2jOAeDnxAB6U
DVuLGaXHRFrQgwwC/qTKIpZ2giK53y0nFohJOaK//SdYzVW0aCJ7TOQginyV
k8GGYWBwXR14fPj34iQnH8d29C5/Ok+bD40ZPVe7BSpSOo2LSiSSDjLSbYL+
I3Am5SDxNs4vUBE2F8wqItS+jyjvvT+OxIzRjipWJi9eFo8m6etoltlUkjmh
HbZVkmTsd+EqXg7d+RzBTM1A5gEdQ1V9WeEJHqZ7C0TydpNRqNLRXit8MQ3V
vJG1Pvu9H3qvQvO5isyA33OD/h96wdAukWRuOX/2NYllLV9OzsyPd1jLnio4
iZxATwor7L+eZiRFUp2Yljf1pHuv+ixjyp8fjimq27lcRBVfTVq4dC3so2iB
sctSoJXXuC1zedjWFagC9mVW+x7CN9b9W8n/AtPImEcWHcyJpkuJwKfk5tuj
LftvcuHVdnruRKtVIpcEOtsQQKwqMqezHa/1ohPAQVCPmDViopWaVX+VL6YB
QOlnCKM8XOAP3g1zr/vsdHgd2DPcrisrPpWXggqtvFBxwpRR+kUIk8oGoCO6
QK9wTcRBpHUlEMtfoZuyPg+sBS5gWFc9G+Pe13evU3jZmVwr4QTdIMCpaB+8
E2VW+1tMvlbMsEoWn/21S5MybvAxL3/HvVw6dluRdpNRnxnBEYPRPeUzp4VU
/HiEpVA2OCuQiPQSWTZSjyE8WyubxVkAUdfdkCW+77yJbbg6J/O0xKDIlCj/
Lwl/cgLoB3UiSWFEzbZhSaeKEgtEHytRzJZWeST2QQe5mTBQLYTJFAdHLmqH
Kdp4FgkmyslxiUkLGrrXr/npVtrUyv/sUE/IzFUBAjtd25JxQd3WuGA5qlWW
E/Gl5YJNTTUw8azgB0s2c+5N1UcPT7LbYbYWy5t8c1vlP9S8nl4aXJtHLH2z
fmGF7S8o+qiAdf4DQSVIpYLD5ZJOQs5jyqY14GTnPzEuvIOQ84lXW4jqHEle
53MhBC59lfm11y16Rpq5zNW0xOvi0H/8vlUdVG4apJWRG3Pe3iw6fAerrapk
JUMKF7ZrkCAfGFK459+kbxY+Z21Ax9eZC6Q1q/Zc4gRU21f6nOMILyWxyEvP
o7FdMPcP51lMgnD182B0QgN3kyY+Eq8KJGkBUOkxB5xO6pRkATmE1YI+Bs3b
AIRoK01XOFwREwMNZ5sWSdX+mfhLpB1EELEII7xuA1rmtd34+1jjaRnSA4sD
CTe7HGKmIoh6O/MeYOWuG+03BwoaEVuNiVsyZqFFyG3znr5UHgulWfqeyRIw
6XOyk49LOYN848XSItupn6XHspM69jj3eoMdtj/J8XfohGb8j6zTSYuyPePx
cDWQ137/fkAlxE3S8U5wNin0+olp0UQURrFL1SgaBMmXC/UDp4MukJAEko73
gGVfXuelBRq/Y4h0vYtjKB60FSM08cK3y0exgYnErJvw4oCGFHC/1Jr2bBgc
FmUNrPScic+2DiwIjN53XlJoAqfddMc0yDt5RzFo2TH+qXURGqY1dMbE3dwV
OjoZEkuwsR693mG1y1XJtwV9efT2rPzqpaU0cKEamfd+x3QuaVqTy5i1mLPS
JgXhu3Uvxx37JhdhG5thYZseCvHRGf+DQgI22moSjDHmawoE5WPUifdzDK9q
GCUZoiqTiKw8pHZb+YIu+e/i6LTT74EFRKLcLzDWYk/zSwIgzApb6FMH6wDz
/SZtinvI99Gj30TuGTjlRrfU2rIdtbwTV5KtrFooe1mtZcRrS99AY4sheStx
hswNSoR8FzTHZlbLioJiJ47yMKvdaL3oEycPcpUiY/fvKXCyI1b794vCXbaW
EIrlmPaG5fuU7O4H2uxfV+GZV9aqd5gWO5NasUsTg1JOGtPtZ0PAo+v8QFZu
DHw1MFYZiYDlSy+7lhaeEH4lm/rZpR1FLmtjCWdBbQ0gL6jGJoTgQUlFDiPT
PF+GCwmMEjS2rNsde+du/WeMerMzlZeppM1khQ9dNzTqTxCaO1p82LdWtGwk
Zk1FsG2v2VIC7V3/JGzKMJ1UFABF/6NW8asx+VPEmhYks8h/aIZm4i+eK+vq
1+PnvXZi6S9LLrXCYpnTFfAQ4iKk5ys17BsmES2kFae2DuHW0+F6gpPXnWdR
9y4ErIkSHulACWBES/y34BF17EDjtGPPTKsbBVkx16kWwEJv8EymbHZn/i9Q
BsTa025aZz9q+Hw9C704LlSmTTRPz9sv7AJUEAlJP+o8MtbFPwj7/dy9JGtl
Gg9hmhvXtOBDBrxrNAgdf2p5J0n+FFK3GI8LtnbJF7hjvOnqtJEAu0UEBQqY
D+6UI+3CZ34SsPtctU1H8Auv9n7medlitzmibnIQ9WpNuU1IZr2HYvobK/wV
bWFMFGjifcsOvLUvRTB+6+BVPwX+2b2zNg1C/ZZDvh45LrhsFSyRQiKhaCj3
VWmYhzBX0s5eWLBL9+euM+672NbqYT1Sao5bZGVO7dvx1MysrCYRJo16/HrP
n63Bt764EQIVgUsZqwlcsPHucVCXOyb9veP7WWYPHXdl81CQdAcZT4Q/2j/F
EJ3cXGopBn9ogq/huWTirzbeFvpoxRAVyTlIZxwAjpsN1xPw6UntQkRCby9E
TR4bLFEJIZpwjHKsTZqBqXddup0s2UgaY08R6zKAParsbQfFzXRDJkifSapV
VTLuqEa4IDb0w8x/dCP9wL3eIK1c07jgVj3pfkAAq2qLRlKn0x/E5SAILvil
wPI3oqua8gTZbihP/HQrsCo3Bgl00g+hSF2GIKR0ydmWVse/7il4hHU83i02
PflYTzha3xe3KHKf/WQyxWqe/4PL9no6cHMNmDvP+05I9d4yQIZQBMK1UsqL
IOCjhUmOboJTQs6azyZYXU83pu+6nnDf9po473SEWmWN8jgSHav+6qi79RbZ
Kdy5uq5ZUN0ZnkFauCtiP+MRm5M2jrOPmHAYnoD0pI8EYDw07EnN/hSMe9eE
AYzYG0UIASmnNBtrDLkYdQuwrb6Sy9IiqxkikRu2ToXPJOXPOad9MsLZq+VL
lWrzPGBnbrMCGRdNBDn57LULsorTyXLVuZNgY+P0x+Rd7rd/fOdENXMNe2o4
NQwlknMdXsvQlRarKf6DV7y5bh90W2lWIA6pQ9Sz2sjreVnw2dUFh0cT8/sc
L301fEiVmkiqUbKLY0FrdBi0g6wbc6ti0EZ6kWCG4iL6mRNZDdWUEh01xofE
BbST4RUEwVaxXk++kDO01MGmiWvjDrealk2fLPZSBCRtDiE0m/HQyK2epFZu
Cyq22z/VUxEjfGIQV/5HT6zdTZHgMl0/odWxtIwRhyzmAY+sM5GjVnf3fKLG
KpEc0ZID5dolAh2w3rowUhSZtSFoA+4QtQULN4AoXq9nMSI7e7tvxsB3ivta
EPQYyNAq+dc5yJsIJ1J9Asm2apIN+4RkyH7Tt2NVZvU6RWIIP2yXL667pmUV
ZQmHj7y8KG7N6zYa+D2isEHJdixbZ7hvNQ6ZPhiRkN0JS/C5daGJNIwjPi37
Hf6XP+tw9TVN51Q9hyi/vgje/f6Ev2sxl4wPtd+xYTqUr2fuXwrB9T1dmZUv
Exx61+ZRilCmAKqO7VvVJaRe5NdfU3yIjbgb3nUOf6Q1uswLK5t8F9nEEVjx
IvZ3c2uv2XK5C6SU7RDMElAhaQEYTNo94JADrJ8WdrygeId7G/ckm9fZy5aR
1axuDaczRygw8CizKxbkJgqPl9kTQZ34eHHH44oFHUcCzPZGZcRnCQa0MsPZ
YjgRvvHpNKUNclOPLcVZsXH6Sww9uE+WPK0hQXQVgFQeD5WODyVPMPt2m0e+
vu0iCdmIEEI5JRuzLFuexES+mrBhxc6vupAXkQFLGurFGH9mQdWb3XGuZE9o
HzTk5BnLItWtycralON9TwC/SJ6DAny7GRr9AowXGPpqjKfGzJT+E7zHXQUl
XAXVWE7XeWAW7WsdYY86RqY6sXHG9Rqs4V7rKbS0SVsipLE3voyUeqSYuDbJ
o5TrJxcClzwBPr1G9kYaWjP2F4GFvQzqH2pCAG3AA77h1D6eQRDsjL6UYvDG
V6lCkbMrddy/0Gvv+WPIqw6FffqRnNHDUB+qwp2bIE50Rj1kWQegucj5gkA+
QmRrfP+5JLOBaZ2sOesn8KVa6FeTVuG4cAKRZmZhLccz4ALbRYtXMNSasLM1
A6YqX1S6Tce0ZT184zRpF8DMHdC+Fb2gxiQKeYwEpoCR/J8nDcoznKkJp+nQ
Dfp6LQPt4M/VsUwgjt6tH0uxxwbT49JUBudzN9GXDcmgxbh20xZwAjdnzH17
l4lKt98OuHx5TIs5hfoWih3nzJRj3lY2PAAlocwd3HuOuwt/ZsA9ZOGxaer7
c4sza5OB3wO3UaMaVkHCa0ao1YWeD+ULmnzawK7PEiyuW6wcEWVgouasnGCb
vjMVOjRQmNwau5hcUaXyTgSTSY7Z7GKsh4uMJ53gFOHeXmt0ZLHLizogFMpI
+gxFFDHU/qSBSZZeEPlaCXuI8JXa62JsOzLJwx3hs9WwXewPotG3Ieq1LnTC
i/ZUnDhZEf7egumpReq+ta0++UYkmLrFJI27Hww1hjlpbr2zUu0LmO3jqGLH
janh5KqNVjDKewHsqODrBuHsgl4d/oSb+kxzWhnZ2lYs7BWZogc1o7gI3wmd
C1grNhj7lw171u2Zh3aXkeN5lYSA3DNDoxt51XCkPYhtR0HvuULHdzeh0v0u
AF+0XiKkn6e2GpWg/XnFNuuUUeFGIfVOkvJfGA0niBfQafc0mN+ASVR+xgzd
3DCfapcylf6hECnkU9tccSVqg9Dj3POcKOmGo+M29YJjcRKJWXpi0gaQmjOK
xEaTTEPhMHjkUle23eAO+ZdiSceJeEQ1DOF4mUyw0DhMvkDKO4M4fkMLapnr
ElBN4MAFXpaPHJcgF0iLMMh6c30CQG3BPiy/aaDdV0GF8CYwmctPl+dPdcZI
W+FTjE13GxXsA2cOwGSdGLio7Rs+Ab/YjDARsDXNohJSuEO2VbdRgLOLEWg5
n/r0BtouD8TP7yyx6lf/WdWtlRdFcJdVvrA28pPP2cASf4NAkIIiMhTCIqzT
nUr1aJ1UlWUSRIhS944SJztvnX7MFpl7a0yiZlaPNZRnFiPMNEyeQQjc8WxZ
lCYe6sxNqmjfaKEUofAH7LDTrinvXmVQ636m7KQfASznP/Npigt9UE6JozGj
2pQTYHKlEp1XzUI1wAMgB90fxZ4hU7RnND/4FTt2WXgEHR6DYHgiWz0m071r
hfmGXxMR7QyJOakm+jzj+0UZki7Lbdv+YovbrDH9K0hWlAnmU3HL0P9kf1vF
c7Z2J2CykZqDrRERfBI/HYuhqIU3e3ecZgMF7OAna6QUZN7lm2d+P0MDxB8Z
78vYvqQ+wIvxvSDPydjr186kgxrC9k51OdrXP3nNtigFvpCRLBKB6ZjQY4QK
CQ3hQtd0ZYFFUFEU0kkFeCEo4F8jy763xfHVMeseKYKOH4Vc19o5Th9s0GZE
uRReZZ7Hxbbe2KTCuCVuM4JprEftq5Du5SpbnsmmfLpyRj46lGbyssM3QM5u
dVzhLrijqpdG9y96MYgHRZ2Xl7A4szlwxiZ3jVYLovyYFTt8K30JoMhnsLyv
kICJDDCxaOQjeUOIqF0LbP/vkPakjnr99BoqlZnhO4CkdYZCDo6ZYKQSU/pS
MgRe+fos5P3zvL/vUA/8/iQDyhqzDWteFRS0pywaUZ7du5bvPogexVFRd33P
HMswQ0OIxSZeOu1R4DzC9uhiiinX7Dms0vxAJwsFMazN2md78CX+1iOkO+Xg
fU+cRxUqgsFvuKGQQmGqdEUkigm2Hjsd/ED5IetYQuKuJjqF2t8jUjLJULpL
GkMla9VYDn6iMW4fJvRGAP818fWnuG07/tlZh8UxYp4Ru/9bmBt/PPCvuFet
GX3ef2thTkaRbJ264SN16dK/k7fq4kilWDUuMNW+Xy6I+qQk559B6bfGUI1B
qUsOueOyoACjnArswijvlvlcN7TIBivwNTVFT0re5rwgLHE1HyxpYkwy3VE+
DZ3PWbS9+oQae0XR3OJF7qBs6xw0xX4h3rYl/mSUi+4yORQtbI8N9LTuCtAq
OG2XsGky+i5gCzdbjBWT1HryKk7HxjrVZHqf7aPiawYgWmYswNVXKBbn8TjF
uYZPkZOVSKf4PhAjXrXRoux0855wMxUjiCVXYQ8ZyvaNlnvlO8fchFuGTBUr
gd5oXBvn6kEp2MSa+WGkVKzN1o8WhtULpBJxeywAv3dH3UbPNEZb/9EvAAfc
IWwZcvGpnp7HayhhUkqHMRYs7fIQtd5XZO/+35LUnrEgHanhJ7mpjJprMzQ/
zATtXJDwDvdl0/hCKRF9LTGaGFwICZ8BPpJTkDlKNczFs/2buEldftCl7/bo
8bCal+oJRWXyHPLaeAGK2iNxEG/+Y+k1FaHdPu/QMZy5WhKq0CNBxM7xmHg1
LxSkneE9F8iX4HupilrgrMJDMwJRGIEjQDzGcNqNxlUPnM8duwhEN0naMoSp
UywAu5sH8AqrPqeQ7NxBo4dripn76JrUyQNiMnPLKOasCxRow6/OhabRK87G
hq6bI3g9DdTN2RD8N7Y1R2c7vTyp3ZgIfbnKk5LJE5glq9SrPesaLQPZLdV8
sCox3EGcyCRW4degFSTybMwLBLdwrK3cVKBEGVNl464c9EX1gaX2+uAxVMcx
EvuLw8JSHqbieYe67YacvgWuYP7LpZYhnI145b4r/yVIDZAGbGBM+Y0kTT8E
cVdQugtkdr6rK4vMwyXbVKDxQSVl6h/rXpx1iKX+0EyY71B/PFgZZlqBTr6l
zziHdDyo7DHI/Rf1Vrii4BM8xt5S8CxXWitAougohmhRO3JD0CGPO+4Sy3K3
0+N42feh4f2nN/f+knN92lAp8UDz21wH8IuiWTL0HvfYieZiEEzb/rd3OZje
nOvvWAj9TzLhkF72PXy3fNFGDRHip5TqUY3Y04pKkt6dRB5YLvk5TShRQle8
BKGe8ctxuHqJYaLSiFbWFpa4mQV9TfuvOMy5CY2Hmrd/Y+bk9StC6E5RqODZ
5v6gQaDrHQ92FeuvHSpL4tn6hMSMRTxIfp2nxnO/3oit6aIQBIrRl6VSm3gD
w3XUNxCpcP5GNIdVmpVRuyuek8YJb7H9L2L6lqnEktvwtMKkj4vxMMKXWdiM
wuB8w46qdogBfBXt5ScHLgOluYAzxMPjLJOPmSeszw6GnytNhHOfHQRqmv9S
vmZbYxuIvPAjXCtCQ04YbCcoTRTfgBmr2Ec4hKjcwoGHqtKdYOxqZzlTKgsW
kxP+VLnHofifUfmcwD68geYuz7pyQ3znt6YOr1+u4I/JZvL1KWS7pyksCi/X
UKkQuWszKlCbWNVFfJZTgjgFcYlU6Cct20ZMbgUazBeasCBbNk81stUNpDMH
vciZySNJyGVAKqysF2pbgllPOhc5fkEPeny9YzcovtKb8AilEniIViVUJbjI
9FT6lxph4S2kq8OsI44Lgh3bm4JTIV5DTD5yb5sOQ5DQZBF24hZDr/39f13L
pJsZDn0GG3/wyWkMohyxfF1t6ozez8Kbt6Bo4o/Sz4Lf7gsAPNcTgvPJmgLD
3QciGJ8628slqzikaKqPe08sQhsxNRJF6JFY20UUYKgsA/ZbtkGLLkXhiPmT
HCqbcTkDqdoFp52EF9R/glFycCOFPD5yhbCclqGC4dVCZwryxQvMQnqKU2gz
qkSNOZTB6qyjco78kr7kWLWdfbctjlADbOIQXSvagIkuEpRMOcpM3X5knGMz
UDHxRRHGHsY/9MTXnnA+99GFlmUbN2xPIdhEB4m3/zn+Q42QVJyh5sckm1c4
yMFv45hLmPFVtjFBRuruD/Am9UOTysfJ422ZWyKrk8539FXOcHfA+qf0lm+m
5B19kQIktMEHM4VzJM8Xr0AvEVbvbeD9DnI06rKv6X5Wmhn3KXjdKTNdLItF
1DGI0TMVMNocnfDSxS4kVNPsruv48gyIoVkME70QbVskc34wqSR0YoiFwMY7
OTeXrNSZDzEn2NaMxe+Tl7c6UBN7LQjTl2JRwfngq1oQEDS2wGsa3KP/bK7z
z/LyQ9vis8ceoOtvgTT9lDMcwixUcX/U2ZpDoiVpqO/oP4xpNaCNa9duiVGs
N4QE8jvdGADTUrPfPxBp1mSkEQIQ2rrrlsL9J9DCbB0GtQvlHLatLygVRBYj
Iop1LDxxENSjOVKujs2sF0TFaDm0EULWf4EUYV3HOGa4WNP90uEnuK4nsVEU
s3Yrt1dmWORcbfUAyy7Sv/8SwkZBrlspCi9iCYt/jsryoTnzenwUh3sGurch
2r2VBxQk1yFrN9owPV+GNNFpKp9wJu7TyHzqb19Ygkpa47kGrSlVElx+o5y6
Q4aUvfvQXmjHzLilDcV/rc8JoY7rB+eQeeN1Jrn8XOvG3juAfDIHVmiSKi6s
XrTyhI/GhSX4YKzOV69pmaCzT74lGJJ4tmNA1nFSM+ciQ7BK7iHz5jESlrr4
tTE0U//mKwFr6SsRpAubh1DEEL4yjjOHhwe56nP8UgVUEnhBlAa+uq/6u8D0
aYQLLmJ2yHHHQc5MkbZjCJP1yT09UhkxrAXqz39zvQ5/u/1IXx7Og6EjSpOm
aBMsCN2wQW0b6ip4Dc1XudGFaaGyMSxvgT1aVVeB4JdCWPPolMFKKc/INfBM
DGH4uJ1F9GOL21CDaeg6csDHxgc3gfDIPPLjiMCRaTI2Aw7GmC/yhpDzRIFf
kUz/pUQaGYmf85N9tcng28vhUdQalBg1MDQWcPQ0mS9nUR9EFZe749KRM7bT
HAGNg0rcRtUL4rq9MCXmVE2pFcHXAHIrGw0vf1we94XSD8xmPj31WgXlZJJ2
6nqSPyKvbEhSzTE71wRMFONRdYGUNpHAHH8WC2kZS7fmwavkuCHjGvsteFEI
mWkhi6NLVXblGovjkWdYvMoq4KVyAGVxHTUnarNNC4wHpMysT2+Ka9oOIM4l
T0gTDoZ1qofdzBpHDroMiz/pJ+N42ndaBeCiDVXEfWYst5M+ooE0/KnGGa0f
pjR7l2JmsAFRcytCOJjlFPxZzY9fogW+8FJCSJcZUCWFP1R2lta/zEd7leVL
QnxZDQQEmGxG3UW4o10bc2ZF4qtDW7wqyOm+01M4RDtMmiaosOx0x1TGvD5g
Oi9irEffVwXyaQF1ZRbbm72VAJ8rqRVXFvNJC7uxlgVIx0WceG9dyErABOp0
Jxevm6yTUPBLfYToEFiftsunXUNcuoHLQIW9FSrZ9z4tJqYYwLrq0zZKuYV2
4qBJD9cEibLylh048TTVFQLqge7m2MV0zkynJMuLGLoyoRHkqO0EFgw5TxOC
tPkmsCH/bfwp8o4W7Z9tmhBT5SKjL/24tyshQ83jpTm819DjWYJrSpM0TnFZ
wmN+i+XRM822Fl9+QJ0cf8AnbxrtV10EKnHCDMcX7toXBIhjnTA5jOpAqZEl
5dgCz15tJjXdQszFHFeuPSH3pNyQlabsIQpWinH+jcstEKCGTSS/gqxG9DXv
htAZ2mijneNmxQqXE8DErN8MKoIe+rBzq4DeZdMDk/wZ5HAIoXmbj8rEIZoT
EGaxNEFrJsVCPY/4amh2OyYj6OFRkTSPY3F8CGK2agEZRXk2Ip++E+NJwLQK
ZYyjdPG3T9xTKuovEx6gsAt5Qg//TR5AkrtK4N5n1Pr9d0/dkYOYgmjx42be
lyUeok5Cr+7Ks4A1MhkhjYyPoEJEAOiI/d44VicE4PytB8jBjsFUTo7y5ITS
KrWWwtZi0CAHIvPK25G3IQoOsS0ztRtrbsP0FTwD6JuLlL3s2vvEfZcW7KN0
kjlkpE1PBMfPe4ObXoQX111cJ2ah7z/ukGR1UMhQKW7m4BhZ6Bn7SqK4FfU/
LG5vchd7xpVUj5cc12FWcsNYdk+Yfg4x9HKbyleLL9fLKNSfSLgB5srSAdR1
lGM5Vao7aQ8RNWsXl91asDi7sDmaX+d3VBJf8dhb64KF/SEmSsLLs/zcKgLK
xEdf27D1cND9il567ZDupWFj3P5pij8qvcITJySSSEjjA4UP+lFF7uggG11p
pXBlttMqx+WiVE8slrmOoRguh/p+eKunkZo1vpM9t3pmzsSvj5ivW0ZNJm9w
mHDoq3oSd6kD9tPFUj/j9fbB4jHp0S/aNi/+kEV58xuYbeWhWzO2S63RVrc1
bocrDdqAOeOF6gZ/Rsg69nnqvSoUEsCACI0jz01ra8fV9dV+2gSaRkYZvqTm
GybW7Rxq+hpqB+v/xCndNc2f2kKGdKN3yh3Nw4Z7hKnEjR1M2hvVV+nNCp02
STsJ7xjJBtdImLKPFj8BgURr+2EgWX5eEPYi1f+kM5PZhf+ohP8zz8RbNib1
rPbQLE7h+/mkMZsr2pmeb3iVTHjLfnYUBYEH0fMFejkCOoppGenybcnTbrd2
gMiQSkrD5J10/vOz7E7p6Fw2vIsDaKoKdp8zwmuk0Iq44t3PgIHPKuylxndU
EKVp06qmsVuHx0D0C8hJhEfp1ItOfdhazU99xos1dy85VhQSC77JOL3donjC
pzwk8sLDGfSW4AY1VbyblmYKuhA4mRwMCh61Y7wUcskJ2DpjIqRKhcnoe5DZ
ZC0MdVeDZ3zXx9xMRTiHxQ7jZ9s8KTBeqMJwTjIbLAsw0J9sN3QP6kY0nRqe
JkGsu2sB8f8d9hpdhdDgMjpDyg3PTvf7CF856lyYQLha/F2AC8rCKj5CTi4a
7id3eb9G6dkocP41rKA0H/sKzp0kitBvInChHoF47Es5vzMr6mq0MVX4gH73
YvrmHX7sYGOL6xvP7H6g4vVelzHttqxmf9yP0AxkTrGSV9T1YRo4N2vh3OC4
mSObjMbu9Drkmu1FvuPmzTlA13pDA4A0wHGeywnEr9MNyRtFTtFTBFZndFWM
VApyuwbKX9P4Uqxsw+f0M7WMdRdHa0DpIbzUqjplvFNMVnfgbrhdgg6CISjP
AsO4diNkZ+BNKe8K/NaK23Eki3sbYbqnX5QW3OYHsNhnyLvddUps+yGB1T26
FT0pwPk+9CZV7GVg6q6CemmtynZ6QR+nvwCAPME7gNfDC7VZu2WOjjGy6Rla
kCyDOgsuWN7qCbDc128VRHzl/D8L/MHXEzn3YfdUvQ0cHiyJzlokd6QS0uW3
iGD4O1m5fu2Ahu262DJ08P7tNToUJY+P7b650qJv+Na3IeVLbSbhZ5pad0Jv
ewDw418GHUMCUjqIN5xvTE+VJZ8tojxwf5CRCeHD5ScTOwq/TGGS2Ba+/uYp
jAjszm0d8b9a1Ko7kZ/KrA+gItWjHlI4pDSNt1WS8BK64mh89xPtp0mKJAhy
KsoLEc396YUeRB6NhY+ADoQvkDyyVCiVmLxftMpi0OON1zQcrSfE6s8Hcc+i
7O+XAoGdH+bGUJMlpaVjmqN/VWSXedFU/+WlTnQcbsRTv8PG5Z1pf7DsmbZv
s6g0nYHofev9qd+Epx0IHwZKPV/rZz+yYzBabC7F7DCCVnoR4Z6mTToF/rBK
xu5dA7yovyUkSS59mzqT9WN0g5D+6ZEhqcqUNbKGzJfc5wbkAIYEeP2Fjkbq
Fj9m7+pFIdylWvPfxs5OHOOaOi+o4qO3icS84peheNPXJA68jqcTAa7J0kA/
6R2suCal9COT1nAZQIEvEzjLUdeSBieNBVUMFTrJKjKIhn/LZSajfj1+JoIr
RfTiFrp71wB1mukA097Jzb4MIdHEaS8Gj5MyS6T/DWdwvkUMpi9jeI3XROm4
NG9mPART64CUbmz6sUxt/cSYINLzLhZ+HTOSysBG5s8iWHidEc05iJGtYauV
TvEvtTmWCsje3/+rYRE1d+UB1UzmNNczE0AmuiTQbiCCSMWiKsWnM3UlLY+E
be9f7lXXT2dpxozuL0m12JZZtJMYhtRJdflooPEApTwozVV6irUrodqCjcDB
0u6dLXZZGNL7Osl85GC2XPxnwH+c5NGBQ5zvPajJqRvssVIOdEBrXnKoykXH
7o6LuhWrHyvFoO+Z2DbOpp8C+WFCQuZSwujQ5vashTFed3wrDnHvNwyoxQ3/
YlgOM1TiGDiMkP5JXlDqUSBIawRBVB3Im5xu9GFNRNPyFdDx1FCYNkkW6yxw
RqRQv/jrCygCTgWdqkqzX3LIZHkrrTKvjJV4iPSjzSD2r24PSA1DAzbLXeyW
GKege/gYMIZe2htJotRZQyq6OxQ5zaEtcRr3JULzuHXmmqACAXJXqbBJSob4
jGKFIPkTqsLZDxdNWpLzOf9nyKbbGsOS6mljtT+3UTvsPVMsmkV2i91SNjBn
HVA1q8l/F1fL8Lt2r5Xqz7+f0VeUCLe+ErSMoF7HmlHaKWmUijc753RjnFoi
yoPV9N1SzNexJs73JOGu+9/FgkSTAMghS7/xYBz6/GIgL6qXoz76nJy1/u2t
zr7agiy91GMMgybxUq0LGG5+FkuLxRGsA6t5z/62vkIBDnh1OMGJvPXPI/OB
eaB/CYXhGMQwBbfpOm5It03oijJrvpEdF3aiNIP5ocwYQw7W87BQo/pV8AWi
Az9nK9enE+dGeUhi6/mXeT579FZxqMsRvqI7LqycdzRSX2zp3VKXohM5OBWr
bNKDLr7WULqXwPGL8ytf+6e+oNZuIl+alT3RzW0vgSZscgG4vqXgPj0451OI
Hulxrh31Qf6cItpmdRd9cJkY/rjvtkmhxbCKVIKlKi464QDv2UgrvO5JOsLC
mrOJY2Vlbb67exdmCdbrwE371kq12Q75gjvICeCGvtXNgj0ClO7Yl1QDL1Tv
/teoItJFreQh5YJp83fuznwxrQP1dejDl7bA1v9AYVsD1IcoOOsxslSdIZ41
wDIeHWOIuPTNzEL0SIpAbZRzb9lUQ61pD4wcGQyFMIUgfdHpkWeyXQjKZgN7
SbWk+iuNBTYvjoPAAMk/rCheETbg5B0YzFAdGRhNwAs9mcbOKdOmE+gnKfol
az3ABFg8zfUzvucs9jrnFQr8ERorM7vD/z4wsjLoatvAH7DyGFuvJcGl4uep
JvaRcPvBiQX4ylYVH5akXlppD0Fp8dLHH9H92Utyg/RuFg1SYOcHDIUPYhDx
XcNTTqgfonbGpeL7OmDglbzlFQPX9yBtXFD/p75lF8vzno/KCtafe75BsxND
oZKKJYlfm6kz39ZRhylMD4fDauDhuqAtp6tr7ZfU3gqaJq/lZC1RGjPn9haa
Rc/DCIXF4toki8czuuknl7JzAhqdOnUgSQQY+u4FLIM6Z3KDJq6I8tjiYjxe
iPa+Q0KieYgZhn7HMoU64BUgI6HJaaajQam7ONxeBc4MACJnD1kj8x42GRXK
efwRo2DIkfQVJcngCPSrMcDPixuwI2ptTIRlq0Rvgi4gD8F3rjmJfJYQLK9W
eA8jtGdgdrwXE2edATX4G74D4cS1eyvAefcrFvhe0YpFn7Mbw6ZSTDsgEFbM
nnIJuYzztlaXDs9fqeQ5n7TVkuRbMgj0CXL35vtOu6LMIDd34Jf95CNN3XNJ
JM1ZLnMoCVC0a6d8pwR3Xo3KgZoL6I7euLU8i8BmeFhWbb4QRogGdRmOsrQb
U3Bu6ckWAJUOqr8CZx98ewpTnMXink7xSLiQhpp9gOE2Cf2N7WuPkgc7TD70
Ofs9x5D+eiEd14132mKuRCu+RLEsSg3UVzUg5NZyOtBATABnjZSQc5cx7IvF
v7yjKPmt8pEkvEAk4MWJ4BgHBtEDylCEMHJCu92L/vQpbk7udk7jwIbJ9X4I
y16wQZ9ELvvxeiE2oHih1UjkERu9JKM188AMM3mmXolxQkhfHUF0L9f88wXD
J3GMqi0JPkkGE78TSrzCKLnarq4ZhU+X/PujUSM0Z0PDjEsMZWcAeWcGytg1
7zkPB+Nei9c4c7fLhzYOAndpG0+ZJ+AbW11NXKxUO7Ib5c9epk6NYWy6dMAa
VDi+EF26JewhsaU4cjye3ifYYRYKpbj+kZ171W6V6y/CEHCSz8GcQMveAEQW
1b/4YhPWbSBAcIanmtSVHkVqhiQT0ryThi6Zucmcorku2onqD3myvxpsTxZR
qw9Fd8YvNp4rocYqnUFUzMYTS5J5DSMv65rZ9/sUvUUF5D9ZfDQ/NdY7/lrL
O7CMYv4/Wbn0Z2f3MOf4W58d/KmjjPLpOVIeAWxkSsNwPEJ3LK2rmEebdJps
4PeKIiElH0njrGpTAqTguf/2UBKNYRuS9pgGc3fHwaq1gk+S7/ibdPBUYKNp
FZOOFREspWjYJTwc6SHwubPYHI0MRgN37m0B9gIItLOVNJDckcHvQpQgCtt4
AKBZ8rO9Xn7NDMX6nzoaA+GKZLBDJQA9k9lxEbhoM/XienMHZE4algj/y9lP
BkaQ8JqbG9ueI8hc8tLjqPKyESTwBN28dK5Fhhb1G5+BL3J21xV+LQzw2wlg
Ec9KFcgHOgXzSuGO1pso545fank1Mds5t8QKPJoj3ljp6aJ6sLU3KtFkwHXc
DY0D/cO5Z8NTBmCsNaqTcWJPMB0vQmepcj5GXKS4/+Cqwlrym43ZWc7L+AGg
3VduTJl+gOcQ3rNcVSpX6bPSWIgf4vWgOAh23G9l269uoNf8gfuW8ekmyhZq
ZS87PJTTWx6MvdgmAHKXe1g5NcQeWp6dZBUD5SDV2INMPtgjKsU8heoeiK1y
ke/9KiCCIkNgWbr6Sr6p0Two2DLjaKNv3TLv/NpXX0xzTpNWgjVAJAaQKBbF
yLnPBcqDvu4SN2/LjTeWzWcXoiAhDrF9X+kh2whbsDgFH3dpn5WK90v7tx9y
TjFcI6eHGYENtVlhMclAJ902H/mfphm9zw19Ij6v2WCufXFigIr0YLhFS9qO
vKn//mHDngnJNE6Z53Y0aXNNowsTtZS8Dq3IpYrHv8+CGgEp/LK52rBMoauH
xGkiZZIqGP/yg90S8MdxCB/2GVUowoAhmBGEpHeVMobdrlaOa02Tn00KJhMg
KnGr3tq2M64YSmB7TT/Jc1OBNu1hQCVYs1is841cJ2Jwb/x7UIfJFjgkXOrX
IjqlyFFCnyJHjbb2Tlfcmm2JhFnjbNcN9Ca4nhwkd1wut1KYPrnQF9hUtAYb
ZraZcbQWya0yc2fe1H0vE4cZoely6/FNsjjFMiK2ZRsCa3J56HmvA/SsoX3b
Pzs+AM2WZRg0QAUod/heDzvSP+JMMV82t7OswjII9nDfYo9/7KExdXQUyivM
uMaa1OCx27QwIQ/CAAO1tH3nEkbeMv8aVPOP5xSLn9e2KakUNY6fvC+3yL6+
4IphKFGKqnC8TPj+YoYh9vGLwFHjryokLZaMXLA8t+pQaXYw7C+I40vF7aDO
T9JRBuhWeheY0IjX80YcPe+fMOdZ2WtBQrIo5Gdk5qtxCGwMWD6wXjjRG1CI
wQPbB0oeknDRVwhMePz6YM+i3d+RJL7XLdxXSM1cPXeENYd4OUtzynJBJHaM
SAo6e6azfCUGxvcPPBJAwknT+s/EdJeItWNNkymfdK1qwlnpjJlwjWT5s7Ro
cWzVbbOW6GDT/4ZvoRfTcldGYWppVCvT3Aav5bRrf+lRnhnn7mb+z1m6A1CQ
cAQRyClZN5efuBLtl6aGjYSZ0NujXNdWp9u52KA73YAz2rLH133hdZvUOQG8
bADieJOV8x37K6JM/S0eLD0ydFVAb69mDwW9a7//zeHCUY3T2aLkpWQxvIVv
3aEWILIUz3+GvsHCjY5uVma3PFixfhUyKM18WSI95E2O3TYhj8Bq+H5RKCzv
Fc2Xxto9GacwgTRRY4jX+vQzHK0LXHND/Agp8tLD+XfdDimhLMsrQ2MTUOPV
cqmNyHmpLuI5/eoP2DT923U5JkfKofyOLNUIiFbAm0LxMAPoiN7cJBPwBLsc
8P2CVKcQT0MeDV8bh05sw5wjaAbMWzMdk4EIkw/E+UUvnD+PV1JqLWNylzCV
Ql0QUx7VxTaAnYAVfA3Eipq/Qb8P4Ryhl2WAVbF1xhIlqMnLqwqjNfgxEI0p
6su+7IR/gWK3f0D2511UsEoHvytuGnOcON2oqs8dibPKH90u4APECAiesusV
Y+BrPRNDkfHbeyoSYGyiajRxGvrpyYW422JfLmUKO8sqIo4riCSFF1gEf0ho
UkMqwmJoePj4HhIJG+bAxwIRJO2PoovDOGBhJgfaUQWXYciFqBWVMR/n1Vva
FRjvviD+DivpfUY9cIdOksdnlGLh9JizPJSkelQFIAnQZAP8nxU5yWRfjZ6F
nS+adpeu8wt0feMJJZddej+fCU6UpNvb6By+KlW5hpZvwPyn3wBq183nshF4
/8ZDySchSLMDscso2u3/1HrfNMkFRVgIMlQVT+SYNZ7yKF987422rJKKpCYH
yzcmJ8NSgHKzaL0rV1AYEbxuqIMRjyeEoSOAgKA4EYQQ7c1ykVkHlsj942sm
t6Fbfh0P+bw2uvcgiybYmOAazKqNVDHYsfNuOTLKhF+BNsfFRMHTWhTKpmKN
b0L/lZF9ElwqAyHiqL3Uor5f+o4H1DGjMegzGG2kT3FIFhOPl9OB4Vir6DQs
JYL/LCVeJ+MD/PgUSZO1TsmnPWkdkwETIiCmxcTaISDRbXT3xfxCXb/sA0rx
TXrr9D6OVydf6Ke4T4oQLLjtPRXdFHs7HjA6ifUXxfjQyr5cJ/CcFPVIkmt+
DaExQUywxGveNASYD7a/ZH19xlNLhbEQUCayiCHWKE25q2O5F91MmOUlUhOe
ch6LV7Sxn1qiaGj9oMRjK/lZokuct84NrfsMax6VBmYdK2kaHX3aoQ8m4yS/
N0gLINTB4+qktCkOx5IZjEZEOqX4UZDTHc8MGAjBTMtQYW38N3DslL9hDDAt
l9g2xrYEzMWg1vcnwixMjjNnwjLqVkJkwfmFDOEZ6N17LeboXuTxbXgebzb2
CHiawwOTsKEO4tp92i+f9+w1CaUmgeEm1qPxz+s/K7yAFYGpS92IKWkDPFTy
DpYi6o+7zW5uxRrmOhmjnu4d67TSjUF5TvkcGULlzDM1txnovJb5WQrMGOaK
sIatM9koQ3F4SPSzbCLXUsr8whp/o987GzyGmZJnem15rvf+xXdgzd43KxHb
hZhJZrlwYGt2fIPEBCIdRgqrUAuJG/TJEDgPpt8FbUzOKY7gxmatwI5JJwVK
+HF+Aq11PaAEs1dDlPqVoXjesYLsJh2M0g/ra8qmLkTY0vYws4Y8ftQRFyta
zY3UaZF1cHKr8gvJH/81qI2d6dzQpMg/WNBJtrs6OYkdkdQWSTX6ByfJw23v
efgyMso4juNgpP6QAURh+jnuJmByLPOJdd8oz1TLN6Weg2cAd0rOFZkh6MYU
2no9+D7C4jXwePA564tvzZblds8BvK5n6hJay8figktoAUV1iiiyRHGRvdIe
jeKwGhitNE+XcOnkKxlC96ikrqyQKTPuod2ZS8K7fbFhXGjUn1bDr/h1ogPn
cCUraztSxLCoQslL2yNSWMn1cEARvgZU+JlicULkhRKqKFiB8RM7uEsWpghE
KjpQh7QQF5oHupNc3B3dOW4kGCqyaZlcuUguITB8z/bzq9AjD9NAH+EBEHMp
Dc3SPg+pC7D1LiGczj+NgYgN2WGxgoylakLxGta0ViPQ1YASQP5L8ozFY/Bm
eq5vsbCUNcGpVobXLuHbIqEZwLP7uYbMmI+1Pk55SuT4nQ1G2sKWiAOn8/ow
pB2q+fJDwUOVWsI66D6HVA7IbQ3izutcO9VzEtV5taH5sbsXmBAfoOwgF0Gr
zyVQPvm4AByXlCD1tw+lVQqiBABeBs5ie4F95tIejZz6WN8QIVI6vimQ20o9
bf29kP9eWM3AwUluJXTLQECvb51lt48OTxZIZjy2ExX5pwd+q9k1sGHh3AoI
ti79V9FZZ0faJj0WXeDfS364/M98XthUe9L29csmYSF+f3SHY/qgHiJN42LT
zNe+snnycXDtaa/ooa1LNdGLK9N8hUahS+2v0DTFAN+uscZqseon7PLH6wvQ
LzmwY3ckxSSLgprXRv891QNAI69lv5bTk9zRTSneOVSaARJ0P2sJKxW5S3Po
GJ5JIUm/jxDMfYE0+t0o4JY0/gKA30yRFHmJxM8A/Nf7aej8dJ1xTFFCICGB
ARg1+zD+okJmrGIH0M6Q0pViMBh4GXnKmtS7/7Vg/riMlIjjzwd51FQCu9Hk
YBHNcOc8L3tyPp8euqPXtEIk+edoINQbL+62xJDLjTB3BiV2wy3NMrdVW90A
ZKb1DrjH6U5a8MGKvVRU/ug5jPhnL55OmMFMA+i0yuEaPYgsb1OEQHM6v/Lq
h0Wy9DsR1qDh8pz7amdxQi+kgzIHitMBD1Mo1itLu/95ct8lAySadzthXgt6
vLw2v/o8z4wMqmnR371w9LcKUEMsVRI+meHryGUTEniqH+jmxiPA+LyrPupz
dwMFohpVo8cyTZONcKpREZMC08a4j0At2FAC1LlZBRphV5kixrA1P40EQB6E
Sph9KdHM1UT5NfOnPGE7Atl3Ezcm3+BupOdu5nFg8IDA1BxeqNAPY3nFq12u
HJJhiXiI5B/irwVX7tPSI6M3+hKnB2kAYTNqt96utIjiMZd17reBLJd9dohe
/yMiLVKzDaBXQry3jsVIBcAAM8VsfXtMYxaZseM0IyuBd7T0GcbvRjbqpZcJ
eGQWL0x/saY6mSwjLm93kReXjkamwbpMm7Qf9UvuGC+KS03rN9jz7wS15ZqR
FyufrjygvCxSIunY90Ruu8wmLafJXabpNkXoNfqCxYojFWhrvARomugQ5VyO
xM/G/LJuazMs28tVBhk3JKolrJNJY1rE6vhDoiAmFD1grHN23ra0z+CQ6DTR
bDmKPFsEEk29zFe3Y7OAmvpNxxJ5cT4ZXD+l6rBlMEABQwUXvxsrukUVStgZ
tCo+8J2cDb48lIo9DEz9UdvwxZmaGM+jQF9XEJpUroBslRoGTxNmTcvk3+11
vvc2CD0nRoQaTnUgYdJQTkoq32pD+g8viLyMdllOIlRjY5q14dV1xg9r2gdv
Q+RLNnM8BUJRa5vgW/PGBtq+PtFCFhBNQmG4+DhUolA+3wm4ziIEPbKqfNpF
w6ojdPp3vGgl51pJlFrJWuHGnl+Fecx1naMV0hzPhkV37BdXVPxm9r7AaH2x
gLjQkGNHlU7KIe3z0Up7Sk7pOKjUWGAApu2GmHT4Cw7VKh1Lrdrzlzu3m8sx
xLE7EgOentzj/sGfmqDkzi91zjyk7CF+wypDdxRbvaWhH3tPsoSVD4rXyNW1
ZZluTTc7VQvYaBBPnwgkLzOGgkVQMj814un15E5mqJ1WYINyPzasKT3oQdBq
o3l7nAqmbMPKnW780TQosadhtt95wKO0JU/Zt1j1gMFbtl2waGsg20w0iIfT
c5OIax7UVmtQEDukQVtm3EbRbD/J0LrxVoZfQ9SS3jA+Hz+Yck2ioDpjymj2
1Dbrip7rnSi/x9vzxfwjMBQvYtTlzdg7VVMPmseC5BLXjYv+zuDqzad17/KU
88Gule1h6nDNOIICjmK95QSoyNzkLiORnuLqhiTd2cPNx1pqR6y02+v3ByFw
Fr7JQHdMXK6cErp1bBQBSwSkogryCFsD4ckSrMdNZ8zeGbdmTgqnPbT9i0qs
hfFF9PWORzCB7w4ojCTw+vJ1IkeT9fmMS1STditQsUAgTU9HKsoMu0cktqNU
tTbVN0oe3fBT3LMQkUzp2Pa5ITlnshVWbJI4BKU7bkTyObKKC4b6BWrDBO1i
Ftkm00YRAIwgDWN/6gH3Wn3WAAdltn8qhYVt6Axos6j8+hdOZ47dYKYenQzx
8teTNOjVKGWcwQxohUSP3F2+37t/36C/MfRmwTXrIFuZGWswZ471AycuNdsD
FPKmMVZzjRxzWLmKUaT0fCg3dH6igDULnA0Y0435GiMGDuo12ds5HXRNB1M5
dZWTgCJfcKhm+5P5MGkY0MGduIXdzE0vIzuTo3TeBdmdVJz1+piE5WEdMGcy
vo6+ThP2Bj6bABntfV7Sylcq6teHyD3E6iuFvQdoozTW0d1y1IDBfTZDh4JF
RZDE2Y9oH91CJ9YkKuFYZTVGwembMbJU2TIWWnJx9JQrI39KQF2MK8EnGBtY
sLvoHhajg7deHhsprF1qr+FnzIAVREpyES0XZaNypJZFGHipACerZQFbMeo3
F9G9KvMLOcNihUfW+8P4es5DKIDRNuPF/lkySn9W94fRD912Idr0ta+aXjvv
sUOon97nJtGt3gp/MIU3W051bmofpntvROHhHZZqA1gk+5O5JE1XQY3g7pwc
OL1x4HjFFN5vwESPe1MiySymI0mGMg8bS1U2AF2wcTyVyVW+2XDtf/jj3eg+
Pnzbwvq5ksmOQ1jEwh5uMuVLJ6uweMsiY5acP9sZTlyaZsyi8XLJZx9OxmKh
BG8eQQ/fyGVVv/8NGgbwnIipTOp5+wDrkWodXUzSBgfdfT9b4zwciLac5TyU
m+jYfTplgF7lOgW0+2YJFF+G4cFwrb1sxY/1fTt/qse6pdm7Npstj981Df4u
+M8EPsFs7LAFdSfIdb7b/tXEa3a3vP9z1snMrUnj2t6WNzboCo9jEJirZ8JC
nI45Ozjsq7+p84EVmivasOqiCzPrQOmGRGrswElyGRe1PF04tKv7d/5jStEl
LbVPYou8We9hizZTYBgs6wMQ4AZT7FV2vPEzTtQEZ0ky7Eflc7SNz0sbXHUp
Pwx+nlobYIC0691FjOjwUd8h9/at6cCLIAcZQaJ+p4zm3cH9xcBx956NgY96
kYGHD0e8Yy8LNM6mTbCruKkg0waz1NE7iWIaLv0MibRGkTqU4vWqYFDX5Cwh
D4GOJ+sYHyeJVAAehmkw4FlNiEiXzKrxZwLPiNK2WtGcM2y2UOe3+7hAVCtQ
4eZUqN44Jn+jVdUSUOS210wlqbA+1LyPDvj+5sBB6vFmtddc8gHXqqJMVKWs
4MgtyW4chyg4kMiCaOihq2X0ccU/IvRqrKFc8Zw5Vw+RkVpha7XTCNPa/qJu
m/+nRyB0+TomYjUXH+R39m5I1AJJV3pzsHA+LQcjaKimjhag+sNs9C7lAlyD
RuGfNyQSgZJMXdDW/EnBcj4kjAS3UuhkySYkwy+KWaN8At+r69azA75cismT
g7x8R2lz9mgQJUAi5F44+DfeB3fKoKAs0MOFk0gNs2cNWmbJTGMmnrjAhHJF
KT5mELKdOQC8PRE9Q+Z/sRfbv9GzS925ptEsWetnitcsW17lTj4EBxCzqOaK
h7RZp0fp2CnTiAuhozPiEcgId2heB4ROp7Q8EGrWBljqMXAVjMQP8DnEXUog
EMw6oQbIX4FtKqo4Hhx/VMrkYuXrf1g9IoCnlQRAdqF8xcTP9Bc/2DGenmCU
RWigJsWvK1Kpk+BSl8F0xH0gbU6kXzMe8AxlMdjRHcROASPfdnW8JsAf794Q
5BaJ2seijxVtFxjwW3lTSxRJC+b6WRExTqGp9JKZWvJhWjv+ixMuDH0nqNsj
vVvmyueIIU3Kjxo1KXY1pFkqpoA8OG8gZnma66WKiKQ5ZK0Zbc8pQBhcesv1
J867OsclaQvn1UAg8IIAnhuRniM8dsQXuG+sUdaY1JsYHp8ynMPqpGw2/cF3
9B//wmelG6ZaUaYuBT0kbGV/mDz+kFygtCrACRt3W7BHgfj7h3iBFhHeHOlz
HMyOVlR/NKNbo747WT/GaxI+JeYrqmstyHOaXwdVN+s8XH8eUSE2rNvm+5XK
7+2zJWPl9ma+oQTeLzDY4LWpjSHWyPh77j3shvg5pMHST0rgEyG5zX3TGTkx
YQ17OgKdboMrop+lagQCnZ0wvzOm0O9wOuzgof93TLKPJYg453c54pGBTIEn
DHhfAzHPAyBCOS2EafVq+OWnZGva5hbfYTw6VKAKE7sfArsDeoEE8yl5EsYJ
F5eAKbcB+zpW1cqCqWJU6AchvTkg0uUpzPzU8JxZpxA/96CESQUZHYfd6Jmy
qjJqJy8jKD9lLwTlnNrwgo/xBEi1/Nobt8Ba6WN6ldlHVigON4oWlCRcbBJi
YdigtBtGCSJCY0yM12RnFyTTLksGEmntSwDx37jiFX/hTKEZmpTqS8+E4AQw
B89D0QvAwOUp8AKTvXRvGQCbvni37hfEBtsEiy4ZUgxbMKCg9Qd5QtBLEj7+
tlwswW3TuDBzB7YA9QjdJpTTIBh2xx/iU2NGMkO2doAxFocQCcMb87DDdgiq
F0hlBzXXCOM+IJ89/mUKylUWcXjeEb4UjMVN0V1hvlD9lqX5WrgI6l+8V9GI
lQVXlqPoTW9LF5sqE7dxDlynQLwD164HPdb1KiaYAa8Xwg+gjzDQwYJf45sQ
NOaS542sT4jWpyMaHOVya2NA1jmQQYvRQsIZ2YFWqzFrMuOKeObyCAIGiFuI
2YDDeKE3obILyvI/ziOL6nntYYhXwUIEbslwEEPrkyxlUfgCUL1nUeki6hcn
5XTrLim62OFTwwP/lKLqoZ3fDMkkBRo7y4ldB5v//72Ahyj8jfwjCst9iGVo
wpk/zJwgR581cnFprmdmK23F8L/XgVrc23iEcG+ll8BF3DDWGMi1cB6lFnV2
+Gh9HAxlZT71ax1oHkF3iBTn0yzla6jZEWIf3ENFybWrFEiZuXmBm+UpTIHs
mZ504fElKHxZ8AzvzV7F8nC4g+feUMrxJtf3qNrwQj5v9TQ1lb7ZKgRu7Xam
ydrcsWXtZSkx682YTsTpvkeL4wRymA6mZ+I/NLVCY6E1Ddr5/P30+tN/yEDL
Xhxl/qYIqUbM8VDcB6pX4QpNUM+qUAV47RuiZ2StNcnvaUgDKlg7sCiLPhU0
ly5gu9+CC6UA3rWGtZQgOrFYbcn+IeVtASKHPLePJL+FSiDgo5ha864nenx6
+Q1Hihyx8YFeK9Ik5ZK/y5mDdlSAlk7ffOjS27Cd9BoYqfvFirc4PsMXZ/st
Lwmf2jC1eK0sXMRyI3KVpnw6HmF2HkK9mytiivTXgs9VFW96yByu/ErDcCEh
NTTwLoPMm1lXDwNJoeNK33qyz8SD2v3Kiw/Yli7JoyyCu9W0ZYEX8l05f3iG
FpRozX4MAqhdxeYRt9UhcLkTDWexN2yuSljS4cqHgOT7PTZOCr1xzPAaMHyY
J2Pkp1+EU6PjYI5GDurx4abnPvrP9hRV1mX6WVpYASY4XLEBZjDQ0D/oRsec
1eW8fbcf/xZaXLY6w4koh0mpDQZaXyA21azgx7V0eYKtHsqH4XlBoz8ELIhx
4bRBr7ujL73GuqDrsi+d4C+pQn6CGWw3EQ57bWaQNEJcjJJthNoHUr8FjRKw
dN0lc4PXkTJfEQ59MalcXhKkvbEu0S4AZFyimWxD9LCvG1/fY1aM8i/tw1sv
eNAtXgk5pTgJ0y68PNPdJL9dFYIV3sXFET9DPsbqBkOleOK2Zk36RFvljMza
JWsMdJXGsPYETvAQrBLF59R1QSCHgtqIjCaMoRNHT2iONE483LA6gtmGnUsX
u9yTP5StPvos9H+tnlx6dl/L65t6+jjSFKAYarC0DbKCXEqfxO/FujFAWGbj
asr+YsO1bRMTlZx03TSaHFA6vOb17j/LbApy0zCO/zD2u7l4Vrss/+IE5CiA
Vh69NyP+T7vCXJeiFJH3gbkB+JZpbvEDO/eGh3dzucOzTSfmnwlUt6xSR67F
AJQdXKTSR4GHIp4ga3irthrcBNf88KGAdupq/5NEKNHbQm8NkYZZdCEQ19l1
ZKCkLbc3XK7VQyfpSov+tHcmRrBILJ7dMAppS6jWjNxjMAAdYzQNudNmceO7
zOsfS78eJ8sxglAoR36xdIZ/NEzDyLY5RebEJGy9A0WuSWs1jYSVe5DdcFZ2
YabTLlDg4vFgxDPE5yDv5FKb6306G2mIzvqjmFS2550tgxboQP3Fd4gw3+87
S7c/IyAu2XOy9UFT2E2svITw0dL7Ba7B+yS9fk68AmjcCpSscEcO769uIKpH
AXf5iIvXqsSCMQsDQ+jbh341WsS+wQ9rnqcy0W6jCOVir+WypjohKDzM3Jq/
uI9rmgCjONLHytiuJoPR6X2NUGdasmOMjznK4+sE8WbrVaRyqKhAUQoDTNqZ
O8myGGvYpx2DSZ52OSNsGlfg+iYtdx9m/ZbnOWW/CCVc5VUysJalPOI05PQY
L8sO5Wlapv9vMYhyzelB2Xe3lcAtIc2Bi5ONML9Pzb660ykM+6z5eoBPRw54
BCouK29kqo8KWjBTQb3lW0fyg05WnV9sZ/NBrcU9ezO11amaPgFRsJrQFFtj
jD8EH7pKnAJtyd9icpd02qPek5deaGZVDRcTSOHmmvrrldln7rKJTz3T9GI0
YFfTOhIvmFDTw7fhGnXsBxWNdNJ0JYOpVmNkZlmAq63y895FwcFey4OXUlmi
bL2O5FHXaQKGzQ7qroOifpTDMreBDDBOs6gYJnO7sIKZQDTtFGlSN+qjU3mw
Sb4XrN5BYSRdJOabgAvYwukzviKi5BPLNP2JZksc6WUkE6nNfSp6o8Qre0B2
VP0G2EDzxlFZl+dwg2FioG2o2MfJhAiNvKFvoET1/v6J36XbS4g65vvaCAuE
9rYRJF2PRbvdbwND3u/N/bdOflHV7g3qO1uL6psg/UY1crezcj0sD/PGyvYD
7XOW0WOq/e6jSN76CyzntW8sFHjN40elVXc2a/yE1qOvP7I/xryiSPi7uDIB
42UbDaD8ILLx6MyXV7c9GIImoNCTVanTBaSAj9HTHJbPRnrocW9VGfkMrRbV
FZXzcIVE82O23VIxgwHoCRKauNO9x5WLvhu9JxSmB8sejWSOizKE4kF58Nkx
XW4QMzAEC/+7O9h2m/ObqAqVjMab7Sk3RmQUpmDPkvyd+SJwb3m8NaeKfV2R
Y4hVsq5vOyaidUSh6EPL3DtddR3zyUHk6GLSxrGk1nOag8MNuGgLTXTCU4HP
hGKkm1iOkMYRbFnW9sTv7kYUMSjUEao6fJJu5r3KgCD8qWQrSkPrx0D7UKWH
lhXsPIfVc7q5uMc9hF65T0Onni8h1iiwLLywXxhxOabYbKpGck5So3GKSTDM
f1Wvd89C6Rwf0jTYex8VF+MX7BAxpO6pepHTg4flDpeh/Lm+fyc/ArI+6krp
dvAuCxgfnO25yisoYWU1sCksmeEQIZPpsvfL+OxzyK+ry+Qh/+WG1Rswk/Wr
n/1JgXUd8q60DJc4fBBsdpJzzEFVeLrGNU0NrpkNbgYZudwUxY2If+DCouBt
oilvLrr66LN50BxP60fHWM+5L52iqTUqcL5P3f5FEaUbLibZoNSBCBSL3eAP
R/CQ8hS/bMsAEKp+pQyN6PJt72+oGRMR5CuzqY6LgFBiPC1z2jLJsuInTjsU
vlS1DdM9JvfFeo6kH83ktLudqwQ6O9RmTdYgDU5VSLGcRZk5T1W7IRTXNsCI
ik2oB/+tFVuuWcDtL8dCjbam6JlRsnctiDVVNHxNQLg6h/dBYYcDW1I9EP4L
BJhbfEsvRcxGum9k/Lm8kj1h9Y2m1VRk47MrJUZx609t7nttYMxbt9+XofOL
0dZ5q8RSmkS3DTzyGqIk8j2OJD9Ss6XvWkN8muna8RS+EkbM6icIhg6jD0ZP
5ySHoREJZdBEwbGTs7YdhH5iuCQW+jJN1caGLePNQB/bPYquCKgoB046D6Gd
6dW1mQJBD/gyzXt8zY8a50vdRyE+6qHfcBqfOla4UWNDjjliUhJfi0OlxK/5
KZmbUCbPNA3vQLgWUoWerGp/RX91yREaY/Ob3qbNGnBvYSVkvZ4XC/WbX1+H
BBio0AjQSAjXCrrMhYUzwu3ySKVW0JQGI8nEsfFpnoZMAy3U6KtMdrgUgIM2
BsjQqL2/TdJ7RI5CFWZ/tRQX46LK4innPNCPfO7aXttgQdUTRmzAgmBLziuz
g9ZsBD17Jh6SyM/yqIqISgJ2mVcQMJCcf3TNtMlbzHlT8h3QYvduiQKY5yFr
l1HNoO1ECwO8cmtnweG/T2dF10OD2eZngdEIIx4h/fkDZnO6zZ0pIbA+1tSu
8UnczjgHB6QUB1ODyMSOXfJ5HhxCMmkNvLeVBPizeMX67t9VqkBidM/Ig/aT
IrWUp7LtSJM4AVmLgUpaml86hpBNk4wqhp5b72ZRJgq/vyD9zF/JSceWhs6c
/7Rh4oEThx/9bnp0ROapW8fyqmBIwpuw1K6ODzDSjzzM5xJXQQwVO0nkBFTX
BUnBN5sPZsgwx87NZwE+0gXso+gWEoT6DtrS7lWzRy3jLfw/XjU372bdTXu9
mLnlddb/Pvq3+E3wFiDfqgcatgF9K/nvON1aEtcxWKZjhVLooZBLivB++ik/
AMAVDFdt0+y9gvW2tjCQbWnFQSSj9P05vsifUhgICcENjJOaxH+gFp+l166v
mGczlY4iySsb+Cw52PkPYIpptDTlBfGCAiDetPTz6nj/lzp5vsh5izR0bTjh
BSi552KjPVyL7M47JftvF5sWop0scwMNjxKF4X9o+oEygTyl5s7Gt3xT38A2
GldIgvoV58xseD7Q7y1OthxE3zAIzC5TO1FmJkJOgdceLrYu9zgkVmjuqQOW
nNY4+tjjHfp0Xjlz/GRhaYct+/dHQ88LF8CmuRidUCpkMbUhfAJs1wgBCewM
2gtmAmPepTrDyAKDYSBgrSpNXYgh32YRwn+4uC40KfrNW391bgSGesnJt7F6
x0iJSUbVFiip8OCuooUUvbmhon+lS8Vkg+RMdz3OpLr6/OBlQ7eLt3kC80Rj
gDjI327xMReWG8J/iZq81iRjLHW+TNVGTro9Z4FQWByuPP7VDCPhHGAHkUom
M8DjKMqX03PstRtx4HmMPk20mtqzOc8qI8kwCYFEix2HWii6YBDBFmBq5KXw
3y9a4TnYz3FrSZKyEXAhYNDs8qIKxvHLIj48wv7NKqB7lmKwYITzeCYrTIjk
HxRIDxXQKmBAZ1EcCscIpxrGYmjwCZ5vT9TPF1c5IVPNOfkMSn2uHHW24ATi
OIN4+T2rAx1ILs/4IQU/a5EyQrlBHiPpXjIwiNq2sY34bxMjY8DV40oCPl6w
sVXIY8fIcayY7hePycQB030eS5EcCqedqruGk4cjpoQySOUIIwBGnWr81TpP
75+ek12FRbTbDPErtpE5cRQ42FFFdW2qFK7ZDoFzqunNXq2FrvMsNYGnosCG
5+qA6pk4szwgGSnEXE4qJkzw4E/W9kg37QGSWRtFjjxv/QH9Ik5qaWXQD0Wu
L/ZioFIn6W/f78PgPd0wdRA5mHnaHF5pqQNQGeym8wPGw9oPfIXYTcEY29nF
SrDBKUgh8girL84DH4po/nXq3T89cg7hq6sw7kz9AHU6FTTopAILn+9DsTzs
riHQ7T6WeNwk7wv9pxiziAyWSAxK/ySK2J2rtwnKwVmkMGAojoEkMzBK3Mi/
Gqe5Xw7fEQllDMPWMCFbu+LivmRJAZYyCbvKm4SPMiXoeT/temEqbGjsSL3X
2oS3KYuxH+7VOrfTQO8aWYaUa1Q1webVosWvxycCRJSqJq1jf5IQKd63VIOQ
9RmYYl8Lhd2cDa9RR70kC0Cz/GDbSbw5HcXqqtw8xUMUUOs0E82Sx3moA1L3
ZakRvOvOe4TEFAVHfYifTov9X/8ESqTNNHDIeclbrU/2I0OLxvZYLxjdElvW
h8YpMS7SLPdtlMMXHnl7Q5DIuP6hUh2XklWq/8SpkWCgNyCFO4c09D6pppfm
zsIfUI8mFa9Nlrfs9VPhSxqR4m5mcoURGXGFTlbfy3pE8aiBb10GND+088rd
w0knhhi7O0aQdomoPYx2K+riFfpfBNfVl2HxlO5FxNLOForr7NxgUvXgEy+5
n+ozKDxKXvHVeD8+Xm54Vp2phZe9zzCQOOYQrRW67V/DzdKpOUwdI6j0+L9r
Zh1Ciys2rUiG0i36UwQlynVP+ATi6rw2Mmk3EawY4IKvPFWnxFEafWVT8ubS
woHotJqR+VVHfi1kXYF2+HtnGe8BXURWL4C1b80Dy2nCbce/Lg8UVKMvlvnv
u0z1DXpSUOYhTKaAyNti7QvR9u+eenzNBdHE5Rv1KQzqGxK4+p3lE8zP1+70
Vl3qtt2BYII3xKRR5CBcFumpceZc8S7KVNGjeOWAJdfj/7Ywq8mccJI9JCWz
oBUURchhmADPM5c3yD+kTuMr4yLg1z0ddGamrKHwqkBtSGx976Dt9hiWCk0H
9E/IX5OY42xhmaJftywUiPKiog2V/Zocm3wqi2LMYtcEgCUhxqlCbRa4ZH1k
QCoEKga851Ghe9ER4SetMmE6F8YfgZvRXo7oYSOTlG8PPuc1rAftdXZTA8Rj
2Nr6EafLB4aZmOh8pO9JC2VH2+YUAAdq2o49OJAnCcY8zlMrUJTRPOftrAlL
XcZEjUNrG+APXc0DnqaHt7O2E8p3yKpyNxD26lUFXkkhYzcrMgEgojOWrpsf
FGT+UBG75KKwNF1WJe4N+JTdjssNKsf7V1Yqt7LwNeUkBnNv+MFAgoa+O2yo
ucxS+1hkjF9LOHT9/swvZ7pgnfYbFB//rcJIJWKV7ycK16bWKol8fHJvmfqs
ZwhWCGVg5ipX5E5sZgCrC/H0FJ+ipDlcxFZTfb81aRcMnrTNHGzYvjGHaG0Z
hMb45dCCHgHpc8h+fXtlzmbAvVfrp4MM7b67LtGQBZ+RkYRWpQygiJHGUAk1
OuqbckajzcqwDUzX8I7DRKqwXaJLrlt6SqwPzeS63nFlRDV/PmKKwQNnhevl
jZVhNYBF/HtbbVA/VuVDoYZ8MQDl/kpO0w+6uruHWwoliJTneoFJVTjawA1Q
RwZ/4e4iO49ltYNwiJezirXKJD6cjjnb5bvcHd3+Pa8RxCneFNJ+wq9aBV9V
MfXU3HpiVphbsGrep/+18ICaYm8erAvqhVEZlXhk+XYcSpooaBQBOWZMSg+B
dKix0OuCrafkc8QmcnEoUHWRY2LTqJ8hCTXq55vtb5X///eJPH4A6+PwDMUU
3KJ3/sKcvYCNo8kuyzkiT9cx8q8mo7KMiT/ug5M2/d4vn+c848wL9rog697x
6N/W3WpNeaOof/3S2BXI89GxT0kHcnghbjO+kDK9PRoSXz8MzqSoPX4lXfc0
EJxzhyuxQ+c6Cpy2f9B8RoqTHkEi37UaAgK+TmzF4wwV1FoszxCi7rxks8VD
ak7GVYMcybvmICJrj1QnQzIthwKQhNTkQMf6ySjJD/qXNW6VpFbMeYWc+RSF
dWIuAo2qQgsJmVo734rSwryT1tVt6QYug5IClyhIUWOrCfOCZEknJZd/ZfuK
XdUIb66mcl24ugtqLKIvQ3PhhpXfH5XeyCjmO7uZlFsW1j0WMlJxSEIc5ohf
2X6d7XGbKHAdTv39uVlaSd689/U0I37gBpZc63INHd3Qneb2uHREM1derytA
iaBesyfjkQimkTJ7ZD5wU5M65WiANfGWeBGg3UAb1B7wu8NuwgoL2BksSroL
/Lra7Qpm0OsUKz3FKke9R8vrkOgRdW4fYbpAfw18E8Goc/xsK5OztDJcQRkG
mtwqF9k1r/Q3etNI5Y1JoLhfXUswLbqPHPMHvlIy0aEEhPW/rFwWIVK/yFFq
WGL7gfyRS6dtTiY0WgxjhO3XbsgoR0zGxBe1RRfYyJhBgkCFbPwyX4RvJZJs
wuMPJKmpxezJSQHSxVBb5FajzTN3Y7jueQgJ0O1zuvPSBQ2XOf7ZiFVSkkR5
qSSdXgsyh4UzGO1l//QVXdIO2Q8jMKVXF9KBJ5rgAJBW2/G5JZHJUafqXewU
SM6omF+bI5lwtkMm4A3tC91LWUnMNOEYKJY4uFoUAiD9Kw9SrmgbKzqrDWaO
epVz507jAdWVahVG8PuTWkCM9pdWTlColmQRZCZ4+ljoYyNneUyoavnfmRbA
0yCFxHGTwHKPABOwJ0UoBWrG253ehDSoebcDgTYRN2xTqdy9EmoAk8HZ2P5C
C8QdliEv6dSA+5yZerOT5cYmWW8UZSOfGrD7pykc9t1cw876s6M8H1NxGbC5
cJW2uL1qRTy6RPu1hrBbR3ZC44wniRWkTcjU94ZQEMZnxoincFnVdzn//CYh
WHP7DABl2N68R7dlWT+gSXGu8N8Jj+ErbN6gjG8lzFpJAD7QAw6q1GP5/VVQ
a+crOUL0wsa9Yqr7bvkNnMnOVt69iq9KnrDZVuXD+NwKzMKTWUYbFrZeaNmC
I/9VF9zSKTo9hYQJd/WaooVLbpm0NeNQWQ0fPmp7b6+9+QuvxR+Lsgnefydf
Uwzb7/XtLpEDZNJzEE7W0KzaAV1FcrbqwiJ1gYnFJXUnh219sl62reIVefCZ
nyPksHaoSRF64dj5KbQPk7IodDG7+cum74tzoL7WCiTFxRXjvxuciZoWvWII
BIQWmpIoPXKqERcMzZkVCREH1yZG6AmXdOCmHnrIvRZSviqJwYcm57L9h6XZ
wVVO8D/0Nfue8nzHt6gm7s1E5QozrwJDRsYY8XWW3c7wlqGELX0renB9IJHe
vKRBFI6wtDilHctswEyAfwefzFoPbEcg0RWo2wNS1CVMkCyuLz0Pl2ZSKxq9
n9v7+/peto/L7kUowbcnPtXUflPvTHubFiclHbLu6Rl43DM/RBkRuppsVzkD
U+dVlEBUAVfAK2X9aA4IiKDx01QUe1u5ko5bWOvpi57jqtNoJjurN9VWWhGW
Fo/4bYL4qAQ9SYlzuzxpY+2MczvLFRtTEiqo1Yfv2kk6P71/doK22VhOP538
53aDRamZkKZogCHIVuPmEFPwRGUdoID4gPmn3ebUKHFyiCPFSQ7TdnCD44W1
Q+6mGdhF/fXRg3dD7I3lADw/wy4ioQkrciCmCist9ajTXxTx8zuWm9jbsKpH
SVpGLceNPIBwyQpFsWm+vZIeJOzfies+NxjxC0yy4S4O1B+xfosOPq7oP8++
XlIWfP3+b0JQnJlEv/nfbmJ7Vy67LAhOuhhN8lwhaymULpQIep209POPqcJc
Vic+DrT50PcTQ9smoRWK5xmW5220sRAyPNDqpH2t5fvdldjKSCQuAxcDqB3s
3WdIUeSTBDwzSIIpv9bjmsAuosu6mxcWlSRSKshh2ohdD1qs2XlfD0MzKw3U
nrDSLNUGD5KjcZit+mPBYQRsws4v5mUwbu27NQHagsKCKBWlWiOctBhsZfzc
PiqPBqx+ZKzkmeOHvf5Be6R3SYhV1KL9d/DJ66WR34HEL+eitfMemjkzH30x
Trj3vi1dLfqOICgz8qQa1yTE95o6u6M4cPbjUj7lwTWxqNU4uELbsb/Ab2Px
SgKpkgwW0bqbph5Z+jF9ABxi9WyKDhIyEEWGYW0KjQUlw56h3UWzJEwO/InA
2RUKLXZx8Z1TXkSi1Tve7iLKkv+1LoKWuU7liJxbggbFu7m9LyRkBo7+9ghF
X2ZbYbwde8D4EEsO05prXmI7bDJJwLrauYtdKjND4hQT6688BHmT3cMrIru1
Qzb5uSZS0icRC61/ZsQCKMo2snECxyayglXcb1T3eur6yE6xOWUamt0U2deo
lph00xZEJ97tH6iULtGiv6kR85eLqBC64R9iXjqD3Jc8H9gVzrN/jJRsfjZB
GYQfavGJf6xj1B2TKQ8zxws9la9UKiG9Q1cIk1cC5ZyzEh4IwRpDJ8uMMZdH
2TqTAo+jpp3r2EtfOS9X/dCXt6pdqUmmfbMTyMqtES/F++XN/JhO8NitJYnc
WDeix8YBFLXX6Yva8AOGaL9L/i+UWLFxtkDQKBa7y8hgR5E3p+ALn8iNlsT4
DbTPJRKH63fsCfhx2lSEzeCz4rxnZT6nyxnyWJ6I0BFBCLPJtreIF1iAlJHZ
NaWHDOA2lIXygNThE+01nqtUBYYersyvVPerxVfF8jnAK6DReVryK0xjz/0r
QqtI8W7iADzKM6lsgB6is7ToRuFelKuKPkfZTqYYdfqXtF+MhwItPAMX8C/b
sOD2pYvPN/JAP1iD+BQp1JYwy3q6oAVDyau5a4Rrwm675B/g9sj/DBVAk28V
s8iVY92wOHBuhZ1/oLhkO0hyjEivMdGcDpLQhOQ4ihYr2J7pNTtEp07wy+6K
VhxT0j3od8muwP0lXw6OBJx9bgW3O+iu2snKVwg/KbCCrILovwCAQ6yYB+9Y
ursHwiQEYIzaa6Qc5S7C+G8AY+1zVA1tHbI1V6rONvfnlzOfKUIznlMQc/Q5
rmYlCkdinlci25K1RFQWhoGHMM+vI6DriqKcQXO1NIs+ur/vhb6pJHL3lY5u
6xnBSDKF6CIre0zSsf9bnKGu2KaRLCJ6L9UwlibkSV0oM9ZD/OrlQtvgZH2e
zwmPQvWeNAJidW6OoMtqpP1ZV9Ou9vsRAkklEW4zQcHO2M9g2FoA7Do83+Xw
s0VuOWz5fbMcApfS0SJjWGzqZ08BU+AwCdkK0dD48Z/c3WpDQXL5H4CO4W07
g8+dzHXGZSF7ZJIWouRZew/3l/SymK+X9+XHX1aBnk5R3OkxnBJ4doTa8K9t
4kihF1SOqjNx5/H2lbdSUiA4z88w/1LW4/1HMrdWRq6HBx7QbiD5pphL5gLj
CKDvxAV9n47mTtm7dZvP1H3i10DgUTRZPaIhGdIvel5kkq14T3IknMiqr120
BeRLC//h7a/VcQHUw6xeekX0cUSodlRXgF8fjdn90fCLpRSEVa1HsKlAnxIy
yeZkRRU3DXd2O/jivUzntbo/Pvfxq4ck9B5Az/SeGP9vBlu9BUCKTsZ5TWjB
hyE5iJro7SVMs7NGa7hCECWwYY4v9G08CuZwYEJYFODrw5qi4hLgRHpzXJVq
q3eHs4N2PzjY3KiX617kNC2ATE5Yil82+cnEwIpW7RxsGkkJGksvlnSLsh+o
IKbIPkgArBbisXIGLj1gxgQgl4+rCNA4/vI98yraJ606/xESKHwHzUMf0uRg
TxdIucxjUxjy4gH82rZAteSf8Flw/f17YtBffJqUs3Lz74NTs3WVj/q0WFFS
XYTSgt19GCGHQ1qlcM8JoCRL52OMT4kizsRkMhbBBWV9nt5JAaoh22GE6BnU
r/VtOLcEtBvjFSsBqBv/4HOoiCw1r68qOE5VSo0Hr9fF5Uhl2KCzvK+VkbkB
Eed51meW5dvJdjE+kp7/iuuHTVJNViFutt2h4mIwEaATFqZx0DFRDpiR+EsJ
MAsoFKQGykz5JyIqW06mhcHNk42JPLVr3Uq4EnQIUHZH4v2/NQmyktkgGeRc
KLWJPai9VfnLfWpG0Z5mqRtleiwLbsLMxdjPEh6ABKEKY3UVw9KSHTI8rlFm
6rqr2VMGzlRVorjQW2uVhPQ4oflBm20HUIFZWHRyAy9DKfS8DxckP8pLL7H2
12HkYh00JDjkx2DF9rG2BUVG8tsJ8a/LlOLGh39+PfUDYVTnoAQNDJ8WuiaO
RwgXTHjgE1wAVKqfIZpguEwHYwBf7BR9wgLq4fpWW9wcjf0evU1OSLRH9L4r
qcP72Y9zqlCJbNJEYmXa1d6kEZqFbmyFDBrCnriTApuv1YTqtoCMJSgBm+LW
b8++gH417x62kUacdh2oOAh8t4VZ91/v+U9VwAHD4GivmoDdoLz4MG+EqPsf
KZdL0KngBvqSnIAVBMsFhEkCjVGj7Fd5CtWuRthQSuBqePkqUFffXJbfGdxb
fprNoabdtza53iv2GEsPDiYJafbsWDkJUa40T9rWEufZYPgNLXAo6+Mjzb5k
R51A5HdDLuGPps4/qv5i7Qa7eFaxjf+VWoedCgIynfR2ClpuYIVXFOjmKyyt
7Pw75BmoRkUZXKKcHzgvWi805d7IYP/5nO5rusA7dN5n96aZRt9KxOOObWFe
nPO19XqQOziCJObkMomnM+bntvb23yL/SfbylLcpeQrUJ0Ejnbu9IccwA18x
FuLE1+r1X/QPBCQjuYg6IxCv3UjAXV0POpwnVMDUTHj7Kw804ZMy8RR04Khg
KXsWLLhyWc9/DhI706UN0rPlNsdFNKPFGY9A2tS1lCTWBwsj9Rlo4Iu+953Z
h9IDzCKdYyWFX3yvR+o7OkVAE/VNRBmNL+8bVgYwVSobUmtFGLW3LdGFzFF6
YMMChN5xUdAGfPM3qh1a06Pvda55oaXlCuc9Q0M0RyUxmWxO9LImzatXfJoT
q266EjjMtiFkGEGa5NedJApOaBv9OgpEU/nP9pUxJbrzN7aHzGSalLMe520P
FZVDhA2MhATpA5/Ah38DYZGmPo14fmVD8+lYmBuNQ7TXx8Otu2D5WevUxuVc
A9uJWnptQ+AlCHCSdjVXSMWyxn4vk95W2CbE3MdGZlp/rerY5IzF8fp94XT0
VRxpDyTYPBMHpYy/fX09vqLoYVBKUiRnxdxh6DtHlUpOBdn0MNz2n68/Wbm6
eQM0AABJILU3qGpuSO1cz9WRqDXLSbgztnXGq4L7GAjIIUgOf70gbKByhMui
f7OIzaxlKrPJBbCgwYGHpog81ejaB5lEFMUsc9XW7XVpv6GYYeJMhnvz5UIi
/r6YYOWfJY5ah1WSRUpoRI1jRxa0HZLyEKRSGNVd5lhaNcGLmnoJ8XQd9AMN
bHpWwiWnSQHVl4YKYXUO0FJBhXXnll4gJeiwX8nQqnqB6tKuAv/ggHiSwE+M
AgDMnFiOvPmIioHENdFqF3x8fk9jT+YxYm6RG+O2wkwP5EL5jjYAi8uUfji0
X1RR4ijaArdccBeFy1e1W+d53n8W11ZsTpOSwJr9cmn1u1S9EhvJn6u/XR5U
1+66Q1z8LEi/ZSfsq42cYl91k+m4vjBLm29u7MN4wJCDcwqxpHc7YazfRDhS
1J6AkWuQVJltT+4iaUhUrHn4aByXBWlj4MMj7QVopHta9KR2/Ddc0i/TaccL
6jDG5Y4TuDgfAvejf6Dl52Q+8gTYPi/lxhjKrrq7lGsmYplOINwDsKZL+QRp
y7itkymASHpI3gEGPb9mFk0bIew5huMS+6qU1t+CcEnIYiBwbBXmIK6ehjKt
cpxWeH7PgBCh8bY6gmbftiu0JGJreVWUn7IEDzbad8UVSTBx6ULtxnGOvBxk
iY1vqh7PQcTagvxeqK7oksIbyTEcCaqktLpvIzE7kST2qaGfe6XzikoZkRPj
X40XLCyoIcdMQZXyc9CpcRgC+gdcb/35H26fK+0kCB366BnwSxGphmiKbNCL
ilSmkcS0pnvPBkdQQsvPCRNW+AApx7Anyl43m8WBOFRz2H6gB8VasqVwPvGu
dESU0vf+45jqEatmtk4g+M6h5pr86pvYJF+zwF4Ibz1LH8CVwK3WnKD04Bq4
hURnmhK1BuwHhcTkKVwnggN57y24JPzjv1XYrWKKYWM8LdRa/k+tRQQYei0c
0Z9cw7ktGKK+GXbeUGztElNhWg1xDxCN53aC2yVuyFQZ7bDZrsr6qBUfJ/wX
gJt5bG9IL2kVgwRUUu3YuoMVb5/Y26ACdAJx3wOhfs9R/9dhsu4Axd9lfz80
NdVs1F5sy/T9Cd66qSaH/1kDoVXYXaIuDQXJAUZYTnKMJpwmIKzNqZNy0nDD
5/KinU3KaZ3V4JveyQKnDpT4R/CRIvQSQAuCvWUJfTT/TliUydFeH+SuhSdp
Sq1+Q19LIKl5T1Lk+8+PxMef4gn0Ok3hq5Tpf/HVHJTYUbm37FlXOZ3fZNOC
OfVO6XUR37C5lgq3nzP7vhAT1/YXD5tmRf6xbiFpVc9UN8oYxOaticPob5zo
tgJanHva6/0zwULp6HmWagcdhdKlFm0hNfpQgpMdfPivLodc78tdmk3zWXxx
gIjbLn2RH8fn8cyKyheWA4G9BAapMZEVIhjSjBp16X+1C/LhPNBSy0twsg+t
sJMBJPwIrciPYflff5fzgtykCgRI13fV3sIytzAboaGm4hb/FBB+TKoDnaAw
KM2trtE693CYUGMujLeTNQMdvGD9V+mnWsYO/v9XMMvPc1bNG4qX0plDCvdJ
1MDz9kCxdS2HgEcQ+hhC0M1bVWNDufmhQByU3fbEdaT3yoIXr5lcEtzM8Os+
iT0wGhMGPYDaeWTvNB9u+lRSHjRIBTmyG00T1NYOIH/mdQO3sw05siW4UdCn
99N3cBIIwbMjPQuqvDHle0TQRnO5wkXLFdG3kJ0jEqE1VYcFRRgvl1/JWgzw
V/7nz44YyRXWaTxlMjZuuduQfyozKLstpUzrVYQE3Rm7J2+UpCe2Nu0fX5of
g2A+4qhP4XKBsKzUcTRggtsNaIXZ4RJnBEuCm8fi3Q98RYOKTWTXmY5maKhF
yk93MiIu32ZTQdRo1iJ07JP9EHDoUL+ByWB17RRKE0kr4fgRqadErzQld1DS
Fpk/LmsJ8YQ+R3BhVAHE8vav8jsiNPLEO24D8nKax7vXQMJ6GvCNOOdH1fBU
0EGKKaYuXQy9k8XuujfKaUMCWx4mYwpH87FvylU7LTvSB+H2m5/1t2Z/qWCH
EsZugNLvjDxRX/AWMrBKJZA8GyNQOwqkM6bVzd7/lcPaqe5xEikRp35asghl
rl4cafSL4z28gbk+TNgGt/h3usJh6L54Ue0HkPJi6F2EnoBJoJmCig9jiQi5
GCELbmANmvpQis2llP7kH2gdxvYsWx41HklN/q5/qWSuGZp2wEvesO48wttC
VsSpM9lTk/LoZoSMoM2wC0e2vxshJMZGyK7dDFZjIQ/yCQruiCebZVkJxJ8Z
Vq5wCLU9SoYOH+wHm3rxJOSrKcY5SF3ZaS7IUj/xmkNylRwKaZLFI+IcCEGQ
n2sFsYTPsg3XrJrhDwF1lO3rZrjLjl7M9Jcloo8uRMnvnLAuyDFBHt9fDTAI
STmdOX6UdTyH/IXlpzQ2RXjz+3YC9zGToZntst4O9wQJ5UWcp0YkqKnO/8UA
0yCWAAMN4ZtZLVsmSiRq5gb+BHZRSwck4W0clnAoZ8lOODUOeaHRyEsF4tEf
S8IlLq1qy2AShtto1G0kJ+jryWrudx+plIvyIGqlk8RJq4gadXjTysf4JNz7
/dWE7Y9FRy292wQ77d+SbqnbQnJYL8hkujB55hZjdWID3Uf6humoWO/wS84Y
TVkEPdN2COdHPqZusI5meYn81avIpen2TccVA08UvP6JrJJfilZZvl2E9gSu
zSfatUbGXlG/t6qJvBwtFrBmeKU6ZX+qmVZ23A9z+7xB90WM42oH1d9ZKLpW
kGrWPpRVCdnDO1pTh3xMzVFRYz3Om6/+KxEb8IBjaW9zu3MwaG7EETcgDbf9
Ovx6w4RWSORcaMdpLS1yb2Ihwu6mFKR8uIzBJvDqhVnGjwYxjctD7rl6xXVy
w/JZ1jlu+pB4cUeuzlEdOId1bfkAnpcdbi7/7hFhuPKGag4v7styHXPf35Qc
kjAUQWv+4X8jck3NFOs4JwCrnDQvMmcCNdl2RGz7Sq/wzXb4fp4HeTsDuzoY
3PUFeu08gq0dBtECCQOfQIs+6OMdfAdZ58VZZUryLRSqbR1utCj08Rg6+c37
sd7nZe6jSaXqVBwto+Kftup0rw8R5aBz2SM/Rc/gM2wg2XqrmkX7Y37O0xEs
mYyZz1f7s3xcodwhb7CsXV3+U5WShYZ5is4yWl2nWuTuaLHT/L3kNN0iSzaa
onXBW6fEbcFStMmrH9hdOx/3Suf3pHGml3qOk6d8gqCeBM/bFRYuCLo7/PKd
aQlDUymVvoVSSOro9EBfjrLHZP5MUO5GNp9pJpurLP2GFLZnBb1KFPsThmPz
Qw4Jir/SwnyLacTUvVjEevRcM2Xtf6YNL3Pzks7u3juf5uA1R7P5nrs8C7Y9
mUbIHkB/ggK6JbkJj+rwKa32y6Bpi7eGM/oLkJJnp6kzYCJsoNT/mXxLk4pz
CosyEKMNyicC9m4oVQczONwndPvF6fFMcpuqMhM0eo2Ng0iUjt5s48SoCRUH
gzH9m/DAjLUNnqPkzfXRV6YqbBv1v5U8fr4cvlANHcp8lmwM/l+o8mcNwZds
VJB3xSqER3vYY9UiiIFCK8rsacpCr89gQzheetujXPB82naafHjbnczqTzFV
K/SQHujnYnCyrt77CZqOb8bvrBm3dqyD9WzOMwZxvUieVPMZqfX85k0G/oRT
jppqZ82w5b/+2/hy3GznvBJtetXmEEyTVUFcx91/XJQKemMgvgllx69Rlm+N
Xt2/0WEdDt91dMYcuQ+dmEWXmiufAAqDp84YaKEfkLljtkeQ3+9bMPQy4TUo
JH7pE7vb56g5AuGg6tbp84EFmRuTYc4WAiYhbz3UG1Crt/SaReRdNSjtMw88
iHDHr748IlF2bbHwGxE5j1lhonJQQJsVaOKHx35pJqu5kj4tpf3Cureb374m
oFPYkve2C9WZMXPFlm69vKM36SHLPRJQ4SNzPt/hlbXWRLAsR2zOjHCNKp/N
Rwj/5NUolPyF2tca7bgiHSEdTQL4OoLiEiXNKJR0gMLy+xf/qUUCtvrac0OI
3JLHlOhxfZrZ/DVF+w2oY5D99VZ4DTL/PPoPET/6idskHXp49WBtBpp36Yc8
ATMIxMrJ7plXneeHHD1KH2GsH94x1GdQ7bBz4FetkP2Nwzy2z1YukS8L2ZkI
R4iy+yGaOJNZ8xs1URQC0fExUytlWpT+rQTO3RWGC5BVEiegWW8smPSaybpH
EdKTWZkq2JUhVeNzxI8c4p+E1SLE/IczUFyvOK9sz/p4Q1UURMooggVtk7XB
o7+EpXKypbje2IaNpxfxE9snDHWRI8uIXMz3sjN8Lu8BtH4lpO9Wz4tlEw8Z
pQd/5xBvJGLbV5Ok1LZMyJ6cOkYO39sh5e4bGwT+aHRFJtSXlBLSUJGDv8xe
yfP3ECDRFybj92TYqzHyGG+vRZFDypvkad5dnpnJ5SXWA3baNlyjSVjvaOXI
sRCVZrfQuPgsgN6Pc2LltkscU1VFwuW8cko9hagZ0F7iHKE9iuYBVhI+JZ2c
xVBsmF4a49rGyGYPPuRXeT/43vTlisXkyfS6bhH3/dcoz6hAHw6lWyPewzh2
srSUUAEGcuQJpv9uC3bXskULxnyRo8iUEpvDUexkk/TfXfjzTBz+rBSr77CJ
6QtY6RSXSAiozSQI85FsfanOk/A4Q3p5nw1QQesnySFjLT+O0a40TwwBuMbw
o1pPMWrABZ1uEEmyx+9Wjma+DHvDcEcmBH/zFD6kmt7SVbP9EAFh/49rq/4T
mFbrO6S3/ep27o/PuhtxvnR9++Ewc/8s6T8iviuUwyvMTrJjNNvkC/v3bAma
jRr+4aide240eIp9L5x9HNRYQ9rzzgQn3BcOn7GykUsEYW9oa09rs36iOK8O
W0Kao8b9kjqKiqivvOSMfjmm2QbDLKO/9GnzvjorngFampZxthCVZWYzKFXM
pN+4UpEXfU7bOkQiIi8eJHzmyjLhEVS5urEjSnRwTf99PLuDy+/OdxHr86Hw
ilp3xVoPl0FaOaOQ/NjM64RilgLdrfm1QU5zAUJu5IWI8/s7cwv1Mn9h7cXW
duol0I1YhmpQ0D8JSec01DTxv4EkeefS/pLwtqSVuwIXhc5o3G0714KiBVAv
p0QKQUnutQMmh5D64WnD9tWU+v09TMgojRqUpB3Se3RdB7EhdDZk8uKlqG28
yxQfgDwpoygmIrUwlTD7dM28LNqvuMMPTwG5tOG50haK6B7jCob8j5WiQ0RI
Jrr0msiFxyjpqk0NsHiRogQUAOpnIsK/8r5KEuzZROoXsYBYWMbiF6OLqkAg
f8694aOnOexNWe05piMBMY4WBdCJoVP1HRNBUV2EI74GQA9EbarSrIH1f1Kw
KcD0VStdBKhHql00Q1HpN47FWP5P5tBYxJJeVCgrszNKJH1ap+7BNB4E/9jh
VEC+/hfflIwbUtb1O3xvZG3MUsiyd5IaFmEIyBe5a2G1JseexcxdjY6sViAw
39NVBoXMzPG+yMyG7qK4Ib61KRNuUzb2cH9X6GqSqbS+3OVoqYq8FusrSsDW
F6j4gLHEw1r2ONfUO2/8EoP77TiTlAd5N0OdM2qqR6/wevU/6vtlVnJX6XHV
G1svUgJNUX6D/ypMzLLp0VBkzROp3b4eGUj8yuVIOBffpUVoRTsmZZfn9Izo
3zgjCZyNhYcnYYbBlcJ91BpTT1kiYHpApftdZ58GtD/hdyApzgPVapnHnPzA
jRSyTBqUIXEa5mhqHLEVK7VO+m8OKnM636AEMO5ES4fLcUFhciRpFXyr4JpW
f1d5tDknqSRY1dUazqMNKifIALLeLM8Z/+PiXMvU3SDBcxhIeKHzZwxJfXsa
l8/eeikHC7VsXrNMxj+V7Gk333Ig7qsQdvCbSKnmdufbxE7Nzu+i/yVLrJ4/
oFS5TllaA3aX3sCCOUugY/NFOom3EXHS4rKDyNNdqZZy8TWBh3GkAdNi6gpG
dsXcqolMHOWAFeoXgnHv88trfoUH5WcAI/ByJ39TJjExd0xCv5A8MLqEUKpl
bOuwiP5KOXtiNqfFxa/lDghMaGbmMZIjaYdt2ZIlTGGZ78p62rGFxCt2WF/N
kHENxNAz0Qw4//NkQpFkoKlGjuUI0dH5A9io9KW4PNfBNRk/LIsEO6chK7kL
QvVKiIPaxY2lDH4RJuFKD1fMGSdGt1VGQu3Gx0B4G8Uiu4/i/D9fM/fVOsxe
aLV00Yf0aC7MW0zml5q6m08NoaA0OLyJKjZqeT1lSd77hA4glFZU6o6jKPkf
53MS5FcIWh0ayMkpSVkPx/L4G3mlq4ccF1jW4eENAEqYiAashqV9soBCk5MP
a+0jZrNLlaCAcc2k9wqegNlooYFL/Qh+givMOAx/uELK7tBlzGlQxLTNKAmK
XjaM3vOUklMTc0XElKBdnhHB2Rko/jgs48QekZYOGBgOTxPoAeKZih7aDT/u
/lJcwZubcbwEOVCG+FlcPNRmXZ90VD67Lm9Ypi4i/Ocaki9HzHDvbVvBtxHz
UKvMrDVNNMcn+p+POkvSwXG2ZR6id0bNQZMolGf1dlyMpZ0tG38hRiuvMvRL
uHIlfktHqwAm5ABiNDHWzpt2TiVeo1cS157mAcu3Y7wtZNyi/45kYLZOmzv5
4Oc0TEypVw0KyXXXr/Ay3G23DJR/lDSZeWjd8yfc15oAqRKzbEj/GGUlRdpy
Rsm1iCOC2pxmOnmR3787bCCohOGRdB0mhD0AISviiWvwzpvsG4K1gDXdscDp
ps4OEsoRqEOOE3OHqlskfmh3WLLMp12uP8f9eTtDtqvX5D/bA0HFCSqN2fQ1
BHzcDoWLoDrxiHLtXI6CzitztfNIJ0x8lLo++KHy+ORuzIGTjEtGg1VUiYvB
B+AeFN9FVpRljGt1rYbv5XfwfVyazpQrliP48+S22S+i5UFRPze6dwFENXoI
f3sEJKzk1R//pg9TUOx7miMaASKIWiGB38b/1oRVl5dzLGSTArT7RxsitojM
ObKvE63rO1516iBNGHUdE1hn/cXSZ2vU57eyl6t8Orws7ZDnM3j1BTbE8M8V
GBTnI7PmN7o83dt8sTuKmglkkDIGfZuB7ZF5RbVY2jc0qTBvxr9rK46LQmAU
AStby9iL+RYKdjdarUM/cHhc2TjQPyF/rVNssrHr3FT/4/9GDDceX79uhRyW
Km58Pm/MuOIpc5V0FmJQBxLbJpgllQV2pY2xlMquopOjIFZozF45LRfPmtAB
16M3imDO+mcZvnM4VEMBqfgljanTgTclznokQv1Y4RAwFWotqA4x7dm4m3BH
lr31k/48JpGSiPWV8d/ny63wR34ceUi63HLazKwWFoSYjGYY9eSjAZvEZvGA
B8X4dhurYfGtDVxKfpny0wjirWclXfQ2mR5+uYwbHZcDDESQDdMmc/FUvDI/
YHyJvPcb0PUIDhZQKV8L7nvK/PxLODM4ETSsy+PZlXIK6k3OTBRULSQVpInr
7+NJuT922pZAjERB9L88GBmaEzG1IdNC3H7NHyp1QVsc+t47BZKm84Rp52Uf
UTiXdqXRjzSVjnky5OIQ6zSq0r3NPF0zB11K1g/SaEqk+/jJsq5Fke6f3p7H
z59UeczCBsAMnJsApcveL68Wd6ZsTqsZYPOewuTcftXehNdmBvO1OgT5SSkV
univCbBDd5XgeEYz1OwD9V+qGcoUPN7y4EqChrnPH4oBOP9EfaCwDzcQScR3
6zacEuiYSuWr/KGaZ2zegvhHmcVxkIs1DjtVNSS5ovC8Erw3Enuy6Oy6c1dk
D7+hU4PNAv37pKbgseD59JrXfMNDcC40FEIqbKntcey8amT9JuNk4T981ANa
gMWwhzj37E5cngXeiB6LkwcxCki8q3uJSjIa4WuAtSIVzAhJ8mKTncQmV25u
XVdrObYugQofDtURLQel/wAocg83QZ7mwtBfQ2pwqToDM8nrPW1SHBteysYp
E9cbV9HVi3Rp4wJKV95SZgYDYSe1+p5d982zDUJIhR0sp2lqkUoGv7+Z5W7t
21/k9Qu8WkYCo6zSogn7H4NzRnynW7HBUh+IUo6OX8TvyJwD36GTbW8XqHa7
v7QD35mqXUA9zOo5/uOQ2xIObvle/z2bjFtAVUn279r4akJT+8OxBrgpxyou
r43sa1tAeP3XPb60YAl1+L0nn6A7ruCXqJ2gEv6KrXB/21+aiHllEfBp/Q8R
04YKYaKHZjPUYCz/L3o61G8qFmBjgw9rRdDKZDcyKiWRF1f+Fc5rpUBJGSB+
4DQcjX+1qinTVPsXU6AQb5ffzZQ71D0kvMAT2KRCR+hxuK0/qX6TsqJCwodG
NZsJr9jcTupNBlY6SUwQkMOOI5w2iMeXWfjHwjJJZnB3T/S++LZqQ4pva+In
QZLuwseyWC7D/C6CO2kqvO35BnsNNYmKUv002h74Aw5q4S8QkVX78BooGuyU
E8tns6GMvH4WDCJwydi7VhhoCaSAQHr+P0dNzhB/upCyXtpY+/ISTjdRTBPx
N7BauCoyX1sekDf3AYDbW8ySFSswzgEg6JXUQJDSdG/dj2Zh9mrN7oJfF+eU
5DM6QVk4ZdE4BbLQRIxkdlcnzVpKyfvohJEqEy8r1GG3aK6/ZcPV6mltTFAv
D5uiPQjOJCT+rbcwkHBSJc3gjnkrkr3jqWOyp5Db52UM96FjaHsfSVV3A5pT
E5U65MO6hLX0DDjFksJOabedse7bh0ILN5YmJN4AqVhQcfoDGYdTAIbM7KRA
mc7iig8lhFhNrVSbd/BNxU65UT5LQ1FOLS7fBBpNNxeL4Y0jCNt2t+U8Yh4N
dKBbPwATS0wB5sdw/0BhpTvjVNJyhzEs0pzOmQpWmafrAqsP48cq6iGucahw
g645m+Kbb//m03oy8bSN/DNfmtiqMJlNMQ0M/DQllxVbqLQsJE8GypbvOUAQ
bhT48bR5cJyHxgZleb2FX5teRF0s5MvhgFHcFhlZSu/eMt3V5TWe0yD7i4A5
8rDGYUHbLeZzSYdB6Ck9VnoFNMUWQSZWXz1bIkY/ohF8CNkrkV1U1aKVo8h0
f7um6DViLBW4FEqjiaERpAeZqwQMGgnwqFjJy/Imy9bJyeyluNySVZLDOaeR
l8c9aCLYGw4e9nbHH7ZzEFk9LL69SNiF8XyMlhBbQ9V28n18O3xnVdKw+Iqr
OyhfXOTjiFreCGQ7vp3+pBX2fFS0zdlCxn5m5RTvtvwDuQ52pPAdeWObQioL
kuNW0bkgD2p+zEBTfKpxDBFwD8htMLz8VGRRqCymK6i2LuPyXBz165WMtrCs
107TIJSG8eC2wnWlnyKhHtnv2xXpwef91AhQLP7wZw8Dyra6i801pAu9vfC3
19zRllG1Szb4yn+qjwn3gueDzNeaHjSNzObywxHwRtavn0U+zsWamp3PdBdW
/rOmsdD1KcMcnAMAl+dQw6ZFKqWcjU9vv3QQywa2AejBt7YimMLBkm28fv8z
35X6eogIQo0In2yPz3mYO521ErDyFaWIgbV1+BoEgy3BvuXu5JvZN+1vJl5P
EVIsybNsqZaYnIm9XV49VbJoD8gUXZwpc/jr5LlnQL7DXLomzrHUilpyB9Sw
x+Z/xzKofZOEmV7chsyxbsrGi7owIrrX9zT8uj3ZYnh4zL/AyVMUpaDOoXNL
KP8DdGEdMPhUrB+Sb5Q1JPdYYcQ1/tBUUAV7ijIkSMVSUES2g/1XIMSQ6F49
ysY3Kj5IaQ25NT+Rj3TUFAdIKU+T4hRplQ4vQzc/XX4dbxzud4y9z2SH7X1N
2Wbk2un791cXFO60IimYvcFvO//LrybPH94lG5v8qHfXdHfuL2odEoAEXR0N
VC3ZGPcNbmK5G23GPY3dFr53JDZoJT1tNzqqATvcUyiUCGmWj8zZ0yv3AMkj
yYDdUPu4dJ9B6M/mFUM0fbiUuWYxMzbv/Y3xs0TFc7JpGHbshljdg+RFpEdL
9dtxKJyVbEm7R4XEm/WK+X0to0BurvC03nJkxA+J9t6d7HJJ8j/DfZdRZt7Y
+M23HZa5+IfaEbZFvNl1SZau3G1tQ/cfmwLuvmfyRfuIWhkxrdYM0TZMNN/M
5aT8E3aqSbb59oDTuhWAzPzqkh4XgELvZbd7GPhsYZYfriMrDFpl2lt392fp
Mqu7bI/CjSc5WkNlqG2qKu2oiBt+fkjmqAKRmM5YZIhAALUp2g3n6XvXw2a7
OOIzcMbt+9OnhRiln1unZned7TAnbdVqr8uJTdu/wInL/3kKNfbWtv9NFs9b
bfq7na9AQ4x0zMtUu+TUp+DaFL5cG6tZ3TadnjFcRpVDrRIHjvt6pLdL4N3G
HgTyEngwj1JujwbKM2UY2h/7wrUKdM1AbFho0jWmVuoqsrDPH7c7+p/e/g0F
1nC0m1SsKh1RSN11t3WWhIZ+4UTRtD0f7mLHMjMu+k3TqZhSlNQp4FgaFj29
OEx5TB6ybG8vVrtu/UERu+RX3HLbylT0nYQrxc9ejYnOxIxhNMEdjoMv4Yz3
3hY02OMT6XRpMODpuwujr7EmgeyOz9JsrDywYYC2cDApSkxuuIpbw7LaJYPF
7vDtkx6NNG05fpa27bJkANOPh7QaqieGmJSgSzA33aPfUjdLSX+vNiNRFPf5
PzZr/f6nyw6TgOfIJRKId0iyVOkxghSHjyGa1iYDok1GePIN00VUxn1t4rg9
7nuNZ9Kp83ItsKJkaxuC+020GTOF9KfWMa62Sqb/FlcDsmYncAdkzhbsn+FB
o/v74Rp5xAIi+SWDUaw8fa2JU2MGid5n+cpCoeVjVCbfcbT8sZ2TeFuXq7JN
g71U72oYE7M/pDXg7zM+gt6/de0lU6U7Uk2ydGsXtTLFyX1O5Ac81+4Df5GX
3m0b4Or08j5JFhjdoQdKvqYdRf49PfsO3QfCG7uTCKp2WQCTdJFfwdV7+B2d
vGMVDRSoxPOLtx0a8u/o0tc+6J+BaHKMxV1/NXacSpStft6bW8HtylwT36S1
6ZQjRElFAN2vxZ8wRHVAGo+pbJy9iSTWMmjVIrnfcuMuJuSiyoCq0ioHdTrz
25KJVOkYlqHv1TTlbaKJDhFx7XJ0744z70+sButXaqn4hG/Yc/hCbZpE5IZh
SFgYyrBjnXY6Qv7vPT3Ra80HJ3CPUDDxYwB7uimE3ONugs3Yo0LdX1Qe8WIa
evywCl8xCUHd2yZ0/8qlY+Y3s5Slttp+R84IhIm7mmtVHbt6eXRL7J95q1wM
/+7Ed/8YWkdc8PjfAZPi6Myj2NAxvNlES4VAJELZULuVG5eU2pmiHZNrO9C3
PKaJVMbV8shcfoRu0QUJvPVpziQzNirpBM9otw0xXiZTJSmxxixEzABfL6bo
9hWZYAjmuxQ0HdVq1s68YPL7ejvTVgIV2EpOX0cjMY9x+hqGkz4lpMFsGEJ6
TlRiM0cTKEJzp+FnGakHrwlwBWPkUyhf+xUEQLSFNrL4V8wCQ/x9WD3Qz8PD
+WvXtJT96bNR4g8b1JB+MrsDI6+jQxuSHx8lbc3DBYbrrsIxFKS9KgJTVc5e
T6p2d1rfp1iR/wm2engNmWyBL0jgk2pr6UVNbHdz3p1XuhEAj4Tg3qbCh44H
c/95YnocFOWl7EI8jNybM28yA9uHRgP/mZPzLYcDaSx8Ma3p+O2gIAJJLm1x
RMoufOltWJUPgbzvOT7D0xtx9sPfCi48fe6r1O/wHXuenNY2w7AyAIc1Pa3N
fj5emOlHChIYl0H65bRr18ZnaZZ51RygoHx6Ro2d7ZiCDOd+MHcwaLBBv2j/
egNxHIUGcc+o3JAmVG6lFlQ3b18haG/BCtZ54RLbTKzzyfwHisK6HlaIGUoT
ZKJN+b02suNo12CW8q0FW6DHyzr0eBNdB3To1FY3VlR0HqJkiT69MU1lik43
o+WdBIf5pQUxT3kgZbIZnLudOCSdSSMGs6Oc8HiQAj2iS2vcvCQkfsQWEWvy
/ydOJxl/o1kpa/eqmcJJYBClVFMYvT2s17jYG6WxKQNjQ5oZFwMo2i2xUsi0
btbFfphtSiD6JClezPRg/AL1Q5n7W697RP7YrfRfMcsEg4pld3kX85dFsdX5
MOqw+7dHTVDWwancxgMrMx7RX+ZWOEnFx8fmjtET0u4pHmsuX7EmNo8jBaK8
Vykl5uOaDnFWXYWkKEYQpl0i6zmy4WVeNggGVU5Q5JBvFAOpu1INUIzcmAC7
MQW5Azq6MXs/320/hZrPtGBs99QwqCnkwEmfvLhGufNHwABdWyLXut6pjXuv
LmY3kuDGjSkOLcnzpOl8F0Ekf0ewTrwjUScor/WpCvx9qJ19WiRsWgryekUv
TCmtj9g4c/nBHaK2pm8ym15zIwafT3MMLWD/ilrToiFSD28RfjS3RoBzvMGK
4xDn374cQbe1ZN8hWUB4Nchl7geeWb0OP9udJYJoDWinZjwceLpx0K6jJ05P
KShjlX9pkqXHkzkziTXAfib8vy6XHJVg4UAh6fqye+pZaSNfWkp2Vdlr4+sm
ooD4kGS6WgKFhfz8BN8J9y4clqKc40lSxYyY6riotSrgZIkVxDLrKQ8LnBoy
rW0I4T7BnuNvdJwvy79ZhHWOZkQ2r23k+DLVf3M9vISbsjZ9nmNoIRnTDaBg
b+mzj8lN8kvUKHSpeGnfm2jh3GF+UIHPAv24bVxZVLRZhsl8Qc+LtyHESbJE
cX/vVq03S0ZvttYTNmPv4ubXRJXnNdHIXylKxZk9Owje2LCG0hj4ob7X3h5j
gkA8ykTI800+Q++jYjhnwH5ORrI7mdj/FEcHZH8uFI5JZJquyFnAM9TWZGgY
aj0noen+IX6qRVXON1Kd5gnxTdiwVmw6zLLoNvJVzqQC7lcMQY/MCWmr6DBw
8pUSzWIXTUfEbliNJZ69aYj5j7x3S45gAiG1+I3YyIs3lLeiwo05C9fg855A
kRq7gdpWV8bX22YkVSy+j0YEanpFu/OLtojA56lA0JSDAO8JsF3BIyy0gc1K
qzD3gkJVD2BvDBQ2ZTdH4TO7f3NIgNPue8TyzGupQOiIVbBeRqrT71m5vxje
2ygmADLbIbGXp+iRkTEIsPopaSjDxOkUOkXwDfwlUzlMi/yA6b3MnWMlAqsv
srcAa68UPbi07JKp+YUFRhziAAftMn3x5Y8IlMlbQGy/w+jsnJ1HkLgDOTR+
Va/z4rpeg3047IuxMlHSt6uUHBgI4lzV610bYn9suNuYd1L8AgzVd5OT9Jv8
Lxd/3HjYZZHDpSN5wOoXHvJRTg5VI6IXKP71MwxfsPJau5FEIs0HjrHiwEcR
RZ4Q8UqRkCF4rqdZiEAAdxxokvUywh4sHRB7zMxlRjFc4r2v0luV5I69d+K5
vImF9k/5Ejt6fMy62V4IC2wS7QFzCVNWBnnDynqfRGsLOKe0aCcwuHKFilqc
nUIku6hqn9S0+HrekPIn5+tZ1Cs+MSToUxrPww1dOKtB/HltWlwXP7MjSzn7
k9d7nF0GvSwhDMMnqLq4IaZRVM5/vtidzEDYEuWZFINot3jP9ccxLkIpLuNu
4TsX2G2KXH2+wSf5zZglTtKtTe57bA1+inyvExjuEovG9W+rkXEi5JyR+FUv
t/sESzpcF/zGAIuIXC926SAHQosS1VB8eLSa4aPj40YlIFq9NYrofIiTIXRf
B6z1OR9h2Cs8nsM64/x5HPo0DKa7e/wCNkufCGIZUc45E/KRDrokqjV1SMgS
LJOQVO1/AmYbOVnTOMTATBYLyZ05weHw4f8p9yKpodwZNawE+cZVSIjgocfi
JXbXt3oFPvlCrL4orUsePqBdOj0orW2/JcFwxfX3Qk3FxXGtnpiVD/mJKQp8
XyzBltJ6FlGVd3LAfJier5UAKwgSPeOM8GzrLbxE/rn1dxXJFa6iCW4YzCTG
DEUJnNuQkMj0WLWH5COQuAFsMqC5HyH/+fJogLD2p/8rp6csKSpcsI27PfK3
3ZPH0wma8eE+cjcTY6xgY8dvS70O7xiAxSfHIBVOpcla2BEAswiixo8TbSRt
eKtZ+RKbJCfPXpxuabFvlyu4aYrMxUevAMzn8j1og3WDc1IkIeEt/MuaohIN
/x4pxERxehkJjmY6DMfNvAvrFT8NGoCQ2xNtvulArd7bW2rvtfwf5y55/avK
v2A7qmKtCCDXLYiduZjs5c5AnIIDXmPIN2XvyaaR5LsR+MDd+O9iXVg508kf
vZv96s122bofOjGDBctmLVddO1FBW69MhedfSRGAygLZgJYmEwkCVUAYH3ve
7fkGTLsHX94Pon/m2e4UGZjiFIErtq4GmFZQa5w4+3mvPvE13PbdinhsH7Wm
5JeRk/OUZ2FfxVyqjYk2+pXDLVFqK2Uy9eFnbgAJlRHZLJJLfILbNt7jjjG7
nKbTIkIy6rX6b5b6ASFZ/A08bLMVvTGd08L+w8DZyTbu0wpf+wVQSizHo8Y2
xczTUGv//kFtEGaGzqRQJppAVXlyM6U/gsmnLCQIcsGC75KlifDUT0ahNopB
+PZyW93TJxYmpI0eYnfEcrsMLxGNll6AAIWrXjuHHmg3W12XCg6NnQUm5+Ww
7zQt/p4rNu6kIYWo4NOh1/Ri5oCUsaoNHhW6KZ/SJXeXkr+davo8kOTODZwQ
N8bLA/J+/F9bTfqy6yOpk46Dox5yIii5qEVcKIDB9loOu30gI1dQTFP2vguO
rOHOpyaL2nvWe4ZIvz+lWKMR8GllVqDih12B4to2fWQaEkNsYoU+i7XHI2d+
0CrCVyt+N3h5j6/rvavuEz+T0aNbg+lhcyuN19DqAa0Ctca6KLmA+wzFbzhw
qKvBgauGIcZB7Yu9lIjTLgwuMxRGWODouor11w0qoZ8iD9K6g8NwJMnA8c/a
ywj3JeuNmj7A2TGi5M+IomZnYVcySXduapXxv5qyf4Zwd3YIWQ6sB5H3qBXt
2rJokhPh927OYV3TrV3hYZYprthwkJ40sJ2JwpvCcm8+cyi051n+3zeTR2GA
lPaptXFe0GnwPCInLhO/8Jt+btUTtHOd020vC8O7JwCvOm2twKAvHlRqhgf4
dIxdaHak4hKW9YtgQvwsYaOmg1nkWd89UNFz7VphTI287WXmFbI8YAxJDiId
ychBbns8AvVLh/ZPFCmmdht+mTrrhFWz2thPNBHhRXOgt2EpeVaIgu7BbFDS
sgVVRn3yHRNRAZ9G+odq/jJQRTbqQ0JMggkgwx4Xnh7udzM5LQrm8I+k22ez
3L1ssZBrEMjPDMhurnqC4CZU+F3mc5+miI2v+Xp7jKLx2BmRjEls+3E+190K
zZ6WtSXEEQYaYW1uPwOBkfU4XZxQuNc1y0kcd+rSvdZx7knTI7aE751O/3h+
OpexdpLFwjGFjUx266urHva4RYW0W4VJXcLlbmGyKMK8sVC8q/sw8JaWeWTC
1RpGwhzyaNX2hqoID3Hc8gMZ4QIljyCzPetXIAy2vK26kair6HPZOyr9mng+
wtrhY9p8eQ7m1FvT2bTgrQWKvQ4zM7vUYvY7uplb9pOcyxcH87uJ9vhEt5y1
5SKHZk/qY+/vhSXElKbIWogHGunt1Z6WLF83XLiqbBkfEx2X/5ptE8sDQBE3
ShGUe0VoFJpaArxf3GtCwHV9AqhK5d2rme5DTFsIqjEfbN8HYHU6oCM7+tMS
KTpJjLZzv5QaWjsXhbjmaZ3WtiFUYroz07qqJ89PLRmksxb3/nyQNvlWLsCG
hQnz2xmxlZsAGd+8V9EXCBTqy5TuneTeJbKojaynSZW01xOLL6PhIw2yZ9Gw
jlu1QoaqTD4LiplQRWgz4cua0T7m7LtzLtqf0y8kXNPCv2oaMCjMeCiHt5oI
6Y+LL8CLOdoodbIiRyRdpzabGvKp7UKShBI0WQjcp4pKxrn/B1VN1CeNwXyM
7tYFqCEuzNFcNda9wup9ihyrVAGm0YbfyuDuFlh+aYVxzKYEpEvGxN1siS3u
kJcZwz7N2Kz3SWfTSe4clq1qVy9+8X0nMzFMips8UpY4ZUbDezeSRXArRWmu
IkHvoC0MLx96z0WDUWJ9Eyvrdi1fzn9n9W5Ac2T7UCUVXmlGs/3G9XhzC5Ia
rBe9LRpgLS1xohZXW8OxU9wgq+pyNHnSZnTFJj06Z7xHB7NK17GDfD3bBc4t
Tp4I0GNTh/CrNq9d55B8MQJOrUvKy17vseaDFBiBwltlJz2te1SFi32hj682
txoZX6INjERO86cL5cS21JPBMfqFWPai8KNQtqORkmC5+0hNmG5HHW572PZ3
1WES+rUkPCWHYu+yk8NiU628hYS6MDLgzTXxLnxIa0y8WIaX4uF5ptINsUCY
PYny2W9oScA7uXcQRURPWQb7ORYZc/M28gIcY4dNe39aahAQ3EmmEKs4ax90
i2hCwqL4WOIBy6ug1IdhSVPtXsxvmRWqtb3MlSP9MN0NWspOVEqNHhj/2aWo
F3A4zYJshZ2Kx2Wnvg+RMXFa2dhQisV3w2lRUDhNC9UNOgtJ3WSACiz7xwUC
YjJRbD6oMY5cfAzmn/xmSSNqPCVjRhTuqy+1B1hG3tTbm/ZGaUcr5Wbbi8hY
m7m/kzwJ1ngbMz+jfBXlE8ZB0eh8oyREwwsVSj3bU3pIYlWV5O8ZTzDltjZU
56ki6WiILu9UuK3ut6qiKDyYtqzkPPOZE/tB8L/f2wBNwUa/xp6+8SeBaG9r
g0rkVy/Q5Jb/vnL4rJTFWXq5y22jmiVLY3+9ccDlaQ8zrVomMDcXposE/aey
NFKKbKokc7dQ592aYBNxoEPcatIlLfjLvBDi9V2o5Mu62LnJv78CfkkaHhNl
KPITxRAE53WMuTKexBiPNu5LOY+2Sg7z6N+ay32k/ftFB/mjbcnvKKwG+g90
7F6mnEx8dRnxfFS2mYJiw3TK3O3rDlzCZFuSmp5XF2k3utaoH0r1eSXgIreD
hg4qHTq6lGJagLz+dyf6a2YtZlTh+0pnuVRq73N91/41IW1K+HDyh+OHH7E7
jx3FLdaWHmX03v8OjI6ljNO7lViZpypMdGSEc+Vyine1/yVEZet97Mu2diD6
vkX693UNdVAUnEb4vTtYQ7epBofR5lVrackjJUUVuZx9mjt0SRaC0kttjPLp
mHBMDT8HYmKOkqlLqwhK9etGGZmssTdfVt2yZV2xrn8BaZgJaDfGZ/AObYaN
f057LL52QwB686nvJlkpuAYhyd4jo/Xc5xQ3mCp15PF4+Gic1eLZ0r0zbQbx
mtcnSFoPhbCbrMfrdJCJCJ8ArJ71pmvQcilWgdtEWXmTrqCHknoCvb0/bRVk
y8gH52Uzg7GRi5+IvFzuS1FrMKVkgYKNfzc2gcj5R6SiRMemPltFgT/Yp+Vc
VtEct2b/8oKgGbSeQid41xtG6yn3xMr0IMXIav0Hb/UNI/t4Ag8qNhVwhfWU
6bf0I5sTdgFV1avXSWENGv4oJxijKu22Mra+F4oOw4sUe5xLGJxJljfQTH5g
Y9g9Mnl/DhCNGF9gBpoLtBR+FP1KqRHThC6s9GJI0zSrrqULUq1k7Y2+ZHk/
4THZATUvWXgbCrsx9L+uj1hR9ip/IoQitaLSN45IiiLoA4T20+UdQhNOrjvs
yGlgL4cs2bf/5HaT8lUyoAm2z7n0bWezJQPXNGgcRq5y8l9x7oA6p5BERXOv
8aDhQMnHnJd5+uQJA2fsh+bjalFN1FdixTo1Dn1ItxffP/UXyG4kxN7Y8XNk
X6ulJ0zkx6KnRN/xaMwwKPWrwrzYFArCvHW2R61FtKMLIWk6uf55uYUFvv0M
Ac2bDbC7Aw11DgX7g9ev8OkKSCeDTRC6LfNZSjix4HudBfDCOUJtcWVJgL3c
7oNswSSy5NCBQ9xlXof7IL/AyvUy/ysXNU5xE9lFq93/UowO/ZH4b3G3Ko3k
dNMg5rZIEusawsmSkRFfzyAIuFLOCP6GACr8bcI433l50T2I6na/lvseBUjS
ieASMdN8U25Dpy2rml3i2d+U5cHB6fjU//+WO/KI9ivdXgaRoBgrcY2sytNU
lPGbwN2L0wmvGrHhEqEAvWWUocoOqe3Hr9ExJGrc4V3bWR+dlEAGeDJyspKp
5HKcceaMKJ3WYvlGNRkmORl8qJ3xSzDf1Qxk62zrzZ8JmqUk6WAYO0kAmZ4O
EredvcFW78QNesWHUPPQMz26T8Rsk63f+syjuyOHwQVMTKyxo6VokvMuv+Zx
JadOFzYnqrZaQWDBvRVa2+m2ebOs9lz9kuHiViAZC9Q/J575YIqXlcCUVZpi
4JzELts5TKxmBJ9VYbO7/3jSh1VzqfXqAHripR0m+IZbZgSLkK+/SNJh/rWd
+EOmNTGtpSpJvJnntuM8JEi+MGcVkGhJ8G6boOBF149+y0aEdEzI3K63E3wk
vuynjcNFf2Fswd9Q2TftKBylFrnBeVVvv8ACz3gt1SrWiH/YoGGqooDVg6xS
fAZYMBeWOa5yW4uWtLHITqSKO53YUye6bIN7azGnCu75kaxmVytNvlUtBC1o
SUOwl7gdhBzSYp9xAvIdDif+vBklEs14bMA5ebcF6mDrWIdImmrXiKrydfYH
TNu2S2Bw53bkiDlL8jJ/RNXpDEsaASH+z/Yu/YaPS7WMBEmv9GgFFuCfSyqz
wFhP9RfxPcznujZkEdAYS8lvmCu9FBjCwxZ15l/Ir+eIKMjpq/LeLXF4mv21
B/AvW8o3nRfYjqBtR86LiKER0P1ZLiIj8HLdlHygVWlywA8sQ6eMei4OHwkF
ZAUj45x39RcczZtWG/mf40LYEQoqexLYxZdpGZHgPF4sOIEcGWuA4T5GY336
VI1PYOMhOOX+VzZZp8AM1HDtuLKgs8IsPJUUukXynqYmflpzdA2NOuB4seqC
2r8HOuepx2pknnjaVY9SkDYUmZCPUwSZd++iZBI1271jnb5OmwLJxlZYUL15
HAyCWiEXVCPPc5onUOSAbFVX8NNvWq4vF4RbP94e17AWvxdy8Ood3uxx7wRp
H1cmbvelCpFOu2dD97eEUE78meTL67cuq4kTs0OAkq6IDvRxuPXDn4lH+ghH
OpIYAu9FWoftLeNVGSi0mGsOJjeQpow4tSQQ1GHOKDKhK7nSx7WZM6hmo5qh
0h18tLcbJ0XvPMdVqHCLq+hIHH1epNG2nWwnfHwwZpSFNWuSrNmtGKqDlOV+
IANvo1rBMFiuzsMoFM/1lTb7/9dk6xcHyYOgq1xyeLTUN/xMJsOaSWjbopPv
LlhFnk8Kht3WAuR5YYLm1/T2GROBdCMUuLmU7tnlQynDK2MjcS2d5bX9pGDG
lCK5lS7bvvi9QlXdESBJMQtiWmug8d5dsc47JU0UjQS3ayqp2LPLAcS349TG
L5oND+L4Za7c+CvuYsOU4svahFrrQtALF27R05vr4OXpAW/XHkvtalnW+mW6
IUX0gGxqZdfg2ll6thzTn7ygKBQpMn2iCBQGap/4TUKrSLy/T4ECvWgt6ngQ
6lQVRWOdEMvTxZFvJ6FhW0Xe/yqAvWtywK7Ep7F6r/xlFosCl7J32dhjaFoB
bY1Ogt7TdpixTi53or2fnls0a0YEjGf5BUHZNpxO46qITAcN1v0Ac9WzLLFq
JAHw5Q48Uf18xofVjECpWLa31rSfqwrccykwpC+9nubxoNFkW9MiQmRf78E0
muTxHCwDEBtvcZJ8ezbeOMeGw3KsFxgdhNOuU9GHcZgMlYCob+kLAhA/r3iU
+3W8/0vetJTcqjMGoiUS98/yn2a2R11jW8wsK96FLEhm08dtESRgKB7C8+eG
KAIfKi0taTiwX4lz16XWx3c6MOkWqEHdzK/J4q+JdyRTX9Q9oXXx6dd0ss4U
ALgRG5NvtfDVf0ZcN42kX0tTpUhG4+Vo3pFfkwfIo4gGz9J27CLpPpH1xliH
5wJwhBQSc9TLjxiZi8mkEHs9qy50uJjQ0vvG6DRFy1JrN3cj/UrYV5uRKNJH
jsxT7Qi4OsJjlN/l9CKMqq3AX7kT/WiQuSD60Cam1xX8bJCjO0cKrP4d3evc
Zr1Loikw4PmeD+NkH97GdAbMw55073hZrkEdhunSpl45cMx1WgnQvo8rjm0a
GeD4ND+QOS5wPSCxdr24WEng8nmthKeb6hnCGGVCAmAErNf0scyqvKQqtiKM
zsxScODFj7HjVhCE4w0xQhX/zhnd0R7jPQo2TcJdFnP4DjEEB/yvMsv6moMV
JJeE+8nmWFE9yM301JLdVNWlTzznHxeJilNML6KMllAQ3yBZGHKCe6+OMEOL
Jic2Pjg1gWgjlV5a7Js0vxF0ndhba7/YPdDPnOb4E85QFmsLgUXARclbt4c2
cmlaWZnTjE5NUhdvGyFUNO4CgWhh8Fs2F4N0LXE21LDg62PEAS9kb00CHIlh
KtEgHH3yMs6WBPhqEFVz0UomfvLGOCPa1OeK2/qtxgeGV3mw0EGIX6xmfls6
snBs94CaxwDI57J/bFedKP8MeoJ2ddDWjIh9tbg+jRrhhITChjOPCP9knEKi
ntKgsvYkO+zTwKI6T3fOiM6zlnShbZto83tUC7CsZHh67hQSEfsdLjj8cC9D
BJOLJgk9ccCtAFq5QAAB1hOD9aXhISNrZIPyho4pWeNrdYXqiaoJbptH4A9R
Zs3sMXaMlwA8rS+BvEbk+QBN/CnkqYi1OLlINz/eLZamG1aIZwRVrXoOvjEs
m9/61ND+9BQ5bzUaQf7T/MoGFBkniRw2EISBHKW8DQgXSLP/n0Wci8gdsZF9
HVZzrjgIumZSvEStWSVKryMyeV2lttTS4b2Dtzsv2LJv1+mxnvkFy+Pb0Ozv
yMZg8prg8RmYsPk7d2/2qau48jM6R+VBbnmBo2DFaZbaTsK7fxzlfhJ+NhkK
jV2fGxKqLeBjBBpCDNyeviRnrsr4MfFZU1axmIRn83Hj6u613Shm1vcUWXkP
T8DpxRdSqBy64STVzsuDQ1g4N7nO4EqgRE2D3hwk2Ud/aDCJnUPHE8hwC86Y
cHcvJBEGoQR7mr/vVMr5Bv6ve2sy7pEPYOgBh25pw48X5234Uj6jNHxFgEjs
DI459ZnOBXt1TZ/8PC++ExIhI7vrOlI5NWP6MaRB10kAn55ZuSLeJJs6M0aR
jMPfFTHZKkUMEqG0q0svy48faQ+qwFhZRm+b565+av71hxFEAMLPztkdN3IR
gppi5Iy5T8HyCCx9WKnFp/bIgLnviVXK4i3CCeWArRjbwpujJPsy3fGbZ1gN
EdpT4jIH6yw/7Fatcrh3e3ewN9Ge8nPd5AkIpClY8yMsZEOvZYVR1vzB8uYh
LJ1rEES6W7Qbzgc9qi/YkZmzSYZVrXcnsQ5FgdD0GeLvRjbtldhPtAd2Vt9i
jMHUESOAAeFFC2lrLzg9VFgjFiDW8Oww9vIGgddxk+ZHe6SpZbgRlcNiWXC3
vCwUFu1ofDNTm5ZL7T1UAdtgGVXl98QlzMFLSxiJJS9eNOf8NCuKhJsAnJDy
j6+Hagc7/OO4nuI0Qy8YIPnow4yN77uvzaxXzKCmFPg1qybitvyjKEF2GhIa
CvXTK3x3XB3nOhsn0ZQzjtknVFdCT1EKMELcm1R8vK3VGRllL9W59IHaQQN8
+2/K/4jJ24wEjbiPgU1kIvOOZdkG5tFOYeh7Ok5tyewkOf4QPY+Er76938BD
ws4EQgPFiMuSZv4PW0zUYu67SZU04bj93acsjyP9xGio2Zql5PCf1MgWeeRD
giztOBxoKHYqbemsz3y2QU01nGnhMEwIygiQwhwp0L4tK17d7nmjXNgBBiXK
1EsbK4yEwk/3p/d/xdLHe1OsbDfsG2yE08W84kZ2lBNDifatBbokNDbnUaKw
2u0Ghrpoelfbnit+oqza8KzBJSl4/gijfsPfUvFq0kprzRrG/XEvImMAftTy
BxFwwJfMDqu7CdB67izz4zPQnc2+lkVtUvItEbW/Ouz4HJvGeH1DdARB8CL/
QyyqdjqmUL6/jZ8oA888D40eHmCvq6W2FwhUTjGWaNgdg/2INrBdKkah7BE5
7jfiyf6P0BoAWQ9d837XLPhMyAlpkSYPLJeI5q2GR1iijxGb6yFlw4atCTLd
kvqtPzXN+hCpuHwIoqq+Asak22jOp/52SL1IoeXKypUwyP9cUyroGj1YU0Qq
TQI35B1JxU813Ot0G19JpIzU1EePpwbh6e3vsqTjC8e3os6mrK2yabeJhlJI
jNVPRiEs0TPyW0Y6zwsFN7vqyg03n3cXMiofFUG+3LEkU425ia6eu2sj8QGg
KEODw1mFIJT8T0TPp61u/MnjS9TiH0KQguGBnj3Vu59C6T3A5mcz/hiIcR+6
++32yeTRFrPqT6CSZ62uo1Tu+3xKg0V5XGXVVhKqr3FmIA0h0Ulzm41ZqpR3
xJjq9QHYkvWb9KUtsVTJMFvgOYgrt5R6vZs01tfF2BnBYrEBnHJRLHbP7022
D9/oUjuSYi/ke5HUJh6xSpEC9q9JIftupuc1fxvDxqcsVW6yyWboNgfAU6em
7+1ZfZmQ5LF5tJLCIan2RtNMx8PnHuBQm5tpEbym2MGQnBe5ZqbF/v/0pbiS
3MaXTBF2O9fyXb0mV0bAmbwJuKeviTuQyqR7b4i53NWGhFUlybORzB9yhJJY
TbEcmxK7DinEYzeKBtfGJu7rXBJ0tuqQdrLmXAQug74e65iekxxivhCKGcyf
TbQHj59mOdXi/9nesTxjWHtGip89Yc4iKV31dbiDfFXbmG2K7lEMmv+m7EiT
l+xJivaBD/5P8S8OZ8IHYAJEixR3RN8JCEsJj29v2M7PXPGuBModkFKv7oQP
H4X5fzruRXNqjnxTTk+W/nfX3OYuSOLDTDoEcUQ41n2MUSJXIitIkRLdrVJz
1Gk8I/memuNTIQj+fli6hO7GAksTeVDik48e1kWLDoyRt5K2c78dwBtw033O
b4Yht7/LIGgfk74RjW+i+9wNubezNMfDzrHty8zW8oP6S4ON1Po/u5eeg/r7
SSc2RLEHmE1qShuj3ZuUijG5u8obvRJStFQrCJHjfFykbdk7YtVj7RcYgFaq
Lb8TFXwUk4MDs/gc1lJORL0GJZjmbC+mk6GL93GkfOGlYVAsZ07DylkOQwtM
rUyw5y3BaohT+HIfgVzRlmqo1SBzzWEREuVmHpji1ObP7auHc7TRX6CJpsNG
qU0kkUXbIQxTAAKV/fee1/nYQm455BibS55dZ4AHRjIGhwNdGF1pKuz0EFsA
xt9/Cg1YclzCw1rGyX0ZDsrXMxJ+Txq1gtMAfj1QACFXksRPkilThJggsn0C
80esO3VZxiY+NNWIYRnQBXXYHlI3w0D3GmaosdMWeCAa8JutOeZvskva3LiD
epqH4H0qjhiKNM2Eq1niehhPwrTzjt7KB7pquBAc6uaYg8j/vCVvkcXKwvv3
uVY0tNpRuKhAy1vqu/BuTo1YvGQSbxKXq3yC4gq/Przj1mn7HtQ1+Bh9sm++
e4xg7wUKONQorgpvyZTSIfFiHKOPzizHVYade8WjcI08M44cvWaqiSnRBi5c
0SdMnqKAFmX0zJN9StGG2cDafGzjdZaYVxMqDeNEhAb6QxLHqW+YlpbptUS7
BOtAjIj++nmSL7MdRCkdlxhjqxNTwWX8G9f8ERMu1V4o+i2lIimlmjxWIYMw
n0YKU2v6uwRnc0f+WxS9WMafntw/fUh/5zt5jTgDs83oquBvzPlUBMZhwphY
8hl5Z3dDIiptUaBBodJHoFZcwIAv9AI2GGTvNTZJKsrrk8/FxzV7LWAeFYvK
U+3v68gzw90J+xNEmPQ3CAF7E9N4xpAKWqGSfqWekJHvrVn191RjePlwpJn5
P4vY+D8rwe9EDgZGEjLG3t+0zFXwYyVHmqNATicvfgOrgJvKcha5F4LInN7R
ankVCfmOTPBmy5/yQXfjhGRbuC5OtXi4MUfu4lmpooRqgKPKTYTyQdzw+TtK
r5qdzLsaerCqghh8VOxZiRUXRmWZ/QJ5fc0xZHx8DMyOjhY/i42qLDcv7BCV
HzZgdcPUBqMbtr3ru6EPcDSOtzT90oGXD00lI3Qr2nTdNu9W37RemwlwKbyC
pfapTQyQaGBG7/w4RKyxaMrU2G+XUPmvcw8z/CySHbT/Xd1UQukfnjH0c/hD
7Txee/yy74Y38DGyINk8or31i0uPsUipwK/CGM3Kv+d5e3BrR2bBgdL3pdoC
J5c3D0odbtRfHhKM2gXCojVTmTYJ3VyIvCaWF6iJCbMHpEqH99TvRXxbh/qY
fL5IvtmkQ4KXlherFoEylurVdVa+7L4kGk/QFdDvNwcTvUzaWrwR99g1JQPZ
SpN9ajRIEqpHwh+0tmsyMg31C3syIeCvmU/eYNokhpoIGnDj3pHLfRVO7fmJ
wMkVQeAA8KyMpW0TBG/phiAxqog/jYSmQ99wI+uLj5xk1ZCYUhdrjtE/SxTE
XZ7Kb6hjhR7mxPlZtG3DWfPdufrBT8YOjujxziRhv1+HTTZdoKZXHiCpRzsq
YJ3lJMzTqMFaagv9yhXAK4WxLGqsOyftdAByL3RF6Pt9tkyx5681Yvj9Zg0u
DHDbO957dQ3ndjReKh9M1Es4K2HTJIJ5gbPaFw+hRhzerMxSa4oscWj8Mgmm
a88Cuxwv5LEl0ysZenJTvLX5pLI4LtkkGaBDuBsbAIBS8LiV635XfhH11X2Z
QV3WK3OU2jTItdtATcnsH18yh1qr0QXss4pCXbbCgnMDYfLR7ydm7hbipQJm
XLWR92/ef6FlgxFs8lysVf0aZ8wGpvNO/JeS+Gt6BSWKt1n4iZwfcACdcXwu
EiNYGnwbXRb6Opj/DoXWVIdFJm0zqrjyehBq4L1X1lo0Zn0aJa9HQFz5OJs1
PhKCBHojhpAJXFJ/LxBVIStsvQn35zVhT+LH5BEflRS7xtVnMkGI3auin1mU
6lddwgD/MtLOiIVjFmr3SZuNKnVhILtt/a40+tL7i/sm2WIw+Vb+7ycD6Bah
C7EfC8lmG2gLGrZV44iTa2ailzv+e+Qr5N0Y1sjtnEK5pyPX18B3OreYvB+m
tat5Wa9nlN/ESJQoDGp66eV2HjqVuHtMSP8lgGR/X8Et42kKuwJftncTuKn2
NmCQqG9HM4kvb0JPh0C3S9VdFdinK7ypSoDjYWdk9L1mF7JDi0UcJAI5Wh6k
xgzZbnMoD5/qp61vrLpEJaDcIZ/B3bDsUBvkshtYnH5PKcuJGtQzKiAOOkLP
d0bGBo8lowLzjjmSs2LZlj75fBhuqhL3o6S9EEAvvDJnjszGiUMC5dGgXG6s
Xlr/7oRpqw8RskRkBcBMi6NLSv4sDVtqaE6G2Cd8t4aER0V6egwdsMWEr98n
tV8/IAlGexvinSX+00c0z1KY7Dc+dD/9vuVMyEa/w/kHg1PpuFltTmT8Z910
iYe8qlXJYkEUwo4ehigvoqcToOHDZji4WWgytqgjpAlgzF41ke0LKuTRiuXB
OJnXdBR6B4Xip9xxwL9dEJvXoSgmFMgApqZx1KL/pPtKn3+YfWRgdRAYcSLh
iv20mFZ2Y/c6WWGKGIBYD/yxiZUunVol8p1bqDlIKWH5kikieQfkuLi0eeGs
mRzBq5ABCZOQckEGQmiaiIXmMtpXJnpV3sgfjfK67A9l4F6DURj05uy6L8T6
SG5Qx9KupEnTQdLJUrzTdp85YQoIEkyeja/SKU3Rmxq68X4ghghTkGFxkQpg
QiAjs7VTs/Ne3pDJKrZQjbvZPp9nF0tp4Y9aCojGzYqXhyCeHsryX8yyW+mq
0Uifol57oAckTaILNhCTAtdRonYBmgh1llsuSwLtnp4UW3VwDoq4ZdiDeHhs
yVPxLQuPFMtjps3hlPrqbkhqN6LesOTYWLEw+IXpyUXv6IgvUImhsJopEDM6
nWr7bqpwZMJ4ZrczALQgjQThGZgvcFCuhPuotBLdIkJyRBO1NInlRAbt5eZC
olM3czMjs85crDYmpA6TBGoam4sMwPeuPZn0wjOiu5jtQKrNK0diL+K2yofR
BhCgtMNwzn8Mod28a6r9GXhCipXNdrHCRVf88d5LKkHqLFwuyra4pDEPBOtq
q8iANKu6G3odxTqOWuw0Kx5sWAFBosEbEEFd8w4+FKEX9KNiGpP+kkIZnSoL
vNOq8+T1R7UwVG3cqv89/JZZqYlSoJeOL8NKLs1bwZxNDWXC5CD78TcVaQAp
IxgLl9p9QPZUzGfNS9MUgMJsjdawrfRl2caFQvCJI8eZdrGDV+WG0/soar3b
fx1i+vc30PDQ8loRNQ9CihRM1FXVvVTVs2Mw1HIJTMTd8N+dC3dAnvI/XzO4
eXBcoBSJQosWofX5MsIUB/2VlwmIQd+OJIYBTAyYlL51Box9kAKWMsP5b2HC
T4sR2zMwDhG5iL+r+4FHsY4xnt1PQqbZkNXlU9I27ZCSBCCF3ghmL+fJ4Dcg
qMO2iMmEnDbM/asX++oMzgWNi+4PCnWISlCPZRve0ZRa/V4GnGinA+AyHdKm
/QqNhHxjMv6w529HcoG+4/JBi/RvXG4CCUNhvEi5ORr4pYQU5GU1MRI4GSln
pJ0NUfh0quaCLwQLtWuN4+GW1HyiHQJ/DE76wlvAPIKAmDRSamoxbasQwmYi
Czve6zflES1VQC2R16gsdWhJKV4lVCkj9BROvVvZtW1G0l+8GzFSL9adpPxD
j/yh/h0V7Aq1mYml0s3TF5xWPmVWWrpiAEmxDsxLr5Xo0sDR0Vpjo/G0FqJh
qto6AH7KICiY/jshld7ERr4lmJBAQ+cmTug7J3S45r3E6U+2HRsAa9twP+xQ
4avv4s7XEKUSaXv5G3BXZ9YCne4BDzEvEhXyNtMMhM1+noe2EvCmc6rPfAAB
anVAvdD1W+jC6d+OoE7iY7j7Nn5rHDMBXy+yHTKSAZGFf5Ocp3YyCxo9LNfQ
RCYXpcYwPGflB/d6KtcB7mjfN7iaUK1sGadQk7rvF/8alNDlFkivlrry0ZX8
2egylt2vpD2Ml5+6hfTS1b4VI/b4PfHWau5mKI8LVs0K74Eci6yWgxDFUM5F
TbIBOGSfaz+0KxzolATsfaHRPUpG+Ua75ajP5KrOZ3QCEKNDkATG6Z0NIiKg
oYS8LbwQxC8gotIW6vr2VJhE21BNryUFJo61K3X/4KlgLMuQF9rcAeqjloqC
MNUyljOyXkjWYtvgB8b1EvKI3CverIJgH1O/lQp/QVGeseYFwmA+9jDujEH+
Pwgm2n86waqVmg5r7ZOPZb8s+JWJ17m0bBx4EdFztLgDjAKbYju9Je134dxe
Z0vYtZFAbr+QFpQ5iWZnnfxjE1HXUUiDUW4gTA8JWGm7t+G2Jus3kM8kAhjT
Do8F1TOw7VYi63n1OdSNIUasWK/LADG5lcVPR3ifPcsVAfADMSmbHULlWKJ5
UWzRRQaaurKTJXCgZnZfKDy418t01ThMI2NfMi81GXdBGzYKD86ASSjJoKKk
IJ5OEE0oNDfTUG0M8rKOWfwZVs+Nuiye6mOJxdIU0445kVc+NKnPXqB7gOoL
3X10678zsiFkrMV5D9MZ0pQCnTC8+jeRbte5+WsCNyBgIz/BI4V8q5BHDvFR
+hjd8pdc7iABbWOW98a6Q8FkUJkV6UITeLBwKMjrrJfRisC6ZQsIeOdcYvb1
/zg9uwWkQGvmAVXGkfZfAl2L8uOMTQChkFddjcTkAxkItwBlCnxrooiwGPg+
dij1EsMJtDJqZu6voYrPyzMKkSOJQ+kIgeOansZy9enxekSbP+gGEM2GdGYy
ypMKzArLRhd2jt/mfJ3AyL2qU4e0t0sgqvv1on0jtHcAi39qeaJpSBF7/03o
I1ozcld0rTLG1d+nsu5RoSYLxHLGJdeaVa/UFhVKVypnrwUyQ8ezsy4OJvRF
5UkFHPMZFS/YSdgVBOPcCa/ninz9yrSYKzG+yIQaGKf29b+qo9PVPHx28lv6
x8GKdeeHM3GACbznLV3/FZop8AuYwZx4/uM0d0GAZNLJLusVmEHXqGa/3VBQ
bh0gCRWK7DlLvjY7tjQ7n/My1ozGVMFqgFkkWMbj/jSGBt0DarCvOJiYBu/9
UfkUtvakPyulNDw3swFQY6cH2bAb4tSLPWUHOOFjCdbcoI+26rmQZRMb2j4z
M2p6Qn7WRXdV+j6GT5qLCSoxVaRZLNCsHtWP+aUIHKDpr9Ku1Z1jdJvRW7qj
VnP4adUAiNRDH/y8BWnyg2k3kGe1Ou+JP2HhrzifQ7HSSaa8e3cYPtgs/PJE
BHzmw7LLE5K0KTIjmcA/FPixgxILOdoosGvGc4DdPtD6qz0lUXu+/ARg4cMl
6Jha6IEPCUPpv4coYo/Le1lzoj+eQCO3ycRGmWwohth4IIZQFxe/VA27tIOS
pPmwvs46QEdTjWp1hdhUZfyJQ+bS14bF5zdd214VGkgw789EWbEnueQvwTFC
E0tuTEMBMaSvUhNHNZZAztAHNkJkSKmxEFmBUi2tNT3qJ04lEnqtdJFkc7Pm
X7FccCmxl/YmJrVBE2qfM6J1YARq4ISJ9kvIuIYxRGsc1pYCXYmKyGxJaP4x
kcELynR7EWJVPIz5JsB9CEcp0sqGcBlTqu15MwDY8AcJjx5pbZGGKSh3FY0x
OF77Rm6h+s9MtGAbmVexkI1vUOEcPY4cScDGtB+m8lyfZBIRWZ4bD2IMNteU
osp5YgoibOG8Se1BctFdV5sbjY7t8ETumy1A2dLeWSvWwBKLkmGJK3rWild8
oTkFzPxtQSW5HM3XjzrQvonVHOdKgjBQCq0FPlDlmmq9YwQoROSm92TextUL
dA1J5rbm8/HpQ8Q89J5K5eq71l1pgPc5buxDU/4+cyP8+hLJD1I4wQvcbp7K
QCvAWHPP94Ndkp5MjFSCtZTjDA2KU5OMmmpPlACmxCTVT1OYYa64INY/N4e8
QVpbFYMld+m7vA28+qtPY26gn1aO6Gc0IaWmtA17IaN2O/EWuc/YJOAD7M2z
6uGjc7SNneZ7oPdTHyEv7j7z5g5r1xH7S6qpXuBImhHJ6QLMqh8NjIgBnFOI
E7dYrYWw/8BQSyhTDnZvURO8p9A0O+Xqy82PxF71F+C7tvp5sfpImatR52yF
MD7Kk4JKNqRejuLsd4WqdFjPo71aNfQQwAdDXVXGkGbYPatmG0n+PRuVplhv
DNH1IqyhkZyaHLgWo/YpeS1kPsKn+uPaZ/S2CrvQBsPY2YaqIAmTe8wZEKm7
3ZftNifqllGi8mqmui7GVkCjLfEPXtcS4wgeO9mOZcnDTmCQWy0/ey8vgOrc
EW/Y7XAo4gzOC4zJSR0WWpxpx+uuga8ZmnVDq3If9u52DOPBN2f5DuuHIkas
puR0L271V47WqmOXi+dfwKXlavuP9mB1gjtxJ1F2uiTbhL7udGRqd5mkMRWt
Ma2gP0ty5Rrg2ptU6t/Hkd7UouimuLNb4MzQqVSm+2PYwjwhyKp/dr1oBVJK
6//9taCNx11gKtFEzanm2ujrtzbi8wKszodW4e3RCCHdQunxW5AXRydoCDpJ
Ho2Mqpo+MSlyYlddRmiLbyHmUcOvWNpI2msE3eqdCIKGgh3FGLoww6I2cNa/
cnTT6x82kiMeeBHjAz8vlmizdP5WCjiBGcdL1dpjLphvnVKm1bIPKo1utNkY
aPqz1njIHqVnxhyDQvQpp3yiXCx4sgKPp47eOhKfdecO9bIO/5LcB2xPp/p0
vuPYhWkOGFgBLhPcvT3EGQTzavfLVxHnWwVFjSHgHNrar8rbpOoXVaBcHnGo
g3FgJ05sLIIV7JKiZZSNV9FAlfhZ+j9iG019zwm6wfq0kIcq027Fs9hNIbxx
FW3veBfa3oWd7gou+XzW8Kymw/PXH+nc6Vcom1unOzg+1+kynEghYFN8F5Wv
NcFczR2i4UboqIgxSz1xuP1Xu9Yp6qrhuyJMetNE/q7Ib3rxTr4Yt/gzHC/8
RakFDAA7U4zAyRxMuB2B3SurNxAC5bXnlcaGLHkkEvsr9nPlVSTu88jlwnWh
/3NKacA67Fm2XQ67yOdR1ClDdqPo+C91rzNX6y+hOHnLVvlmoXaxsZeNzxDE
1HgVyDs4VwoQFS7vjAHUiDMKNTyx3jU1dnwQ3CUWSep0KXcx6rijynogLf3z
wXofr1nPQIRLk1tLcQGB8rk7qMmksfo2/+4ptS7/sBVS1FQyPiZmEBKBKDrs
Wdqwh6jGHZnlW4jaSJdXE8kI8JAAGl+5e9gyDTDKU8CEQP1+wxt9FEki1uAQ
A8nk31hOvGRZswy+Yf1T++P7+Wy19bsaPAJjGFmzj4m7syZw/sKwwM/b+rwr
OZUrMGadFvZxM/PtHiWOXUhi5N2aG3LssqIoNkj8gsq08O/oL+hf3NyCvvDy
1g6Mosiz8hu1qxFL+aLnQQasWljvV0v5GmeHLT2cd3TXJdcVCy2HS6eAT8Bv
szD3RXAMcH8KorWUl13V2eY8sgfzwpkXjoKzC2qcyEJcMxRbtRlGmnraml9k
8MoaJpsGhy70xB6ENkpRh94D2StQ1WcGDWtYjqQK3QiljNuLd9mRB6JeMKnd
Bw6AoMRlrGqXs8vTOqLK/6CnUjDJ/eGBL3iAkyekNyMlCDraKbvslk7qksWg
WM1u13JJOEdQQkcC5WJr/CugTlbuRvOwZ3IWAErK5zSMup95y+MWOvQzNdxb
bkETbdpVao8+JzCgcSFxR9ZUVPkUuwSWWZ1Xf7vhdO3He2SFrtaZKwr/GOIf
mkVPZ+FfPnL3GuJCT6fMfrq6d3BjD9Jo+IA1XSjbnBZecI0Dh5JGKpgfS2a9
bbpW2bLy2bY7yWAqoug5Z7s1ysQsXxJCPbqbcjkWJOKizRhN7bNgKp5WDUGB
dJ0cVWHxse7GQfhV7sF0TdvKW2luNjQaMfGeZMJSuFar7Ozp5VP8jNDFquHU
jY64aOFl7V0iYaH6Hu8Jf9YqKSLS2aM6TsUWsD7lYCgxWdxDlkQ878pEhsw0
ZdNj1H3WT8YOyZS8DV5Q6u3LOepxvIZhjrjtXK/SvJlDGinDvE2ohzfpdyTn
G4XuoSYV/x0YVBnbRiZ5r/l/a++K3dy1jhGc7L3//bPAhDIbAfXWr+EXBIh/
JmY+TrzQmticEy1Eq+jJPbZ6CSz98ou1rSewXJwm6njPTnj5AQU9f6yUPjBc
BQOxYMLwblowbScIX/XW1u7oyknBmiCA9qs5gc1CFfaoQ61+Zk3gqWG5+Glv
QL2RMSKsmk68/StK90gSVVcn+WWJRfZ+qfu8HEx/hR5J/sx9aEu86rGEyk/U
FJ9u+9EKgQl7ifKQRRr4UDJP5hfeBZflDYx6jdMNnbN6zNt6D5J45GCbQwwe
506FdmB2Us6LaeXYP5HYIty6dl+wveXog9y+ce6cSA/bNarhblFtuOtbRb7R
b+mhLPscotA8V5509Paxt0s/1OmDW/aqGYHhNXUN4yxQjbPvujK/aA5p3Q2b
PauPq5BdbG/4HTs4++Ghrx2GsY+l9m9ZyWcsiEe2cz/XbC1nMhV8+AtUYPVP
iYJiJULAaj7X8Yw4g2o/ThZk3QJX7J2qAh9FuWyUWJgH2BU8HFkCDldI/IxF
yxwyD5Bt1Xx/0JPNZj62MQ/V45Iy4Y/T0SV/dT+/WYFgqq5FEXRSgouXujiM
WQaD9KJYLQidL2QUIr452Xlsgk5c6FCQWSBKii0C63vS9O9TDNOhvtDHL9BN
zzqhYxFMBl16PxxR/P8UkPmb2Z5ULZAAKOdURbMQ0tLopjOAkmU+Pl1tdfqI
yNC6J7dnO0NbI7uEvhtTv0NGZr8dIh3/BXYij9cIdDrIz0BSu9K3mmesuMm9
P6qLvk0ZnyVIeISeew5bvcrvkrg0R8VV9OcaE97E0RcveLFZB5T/CbTEV9A2
7DsVclj8wSo8x21GwNofpFjQE73hXzWLYnDVxCVe9cQxTj39Bz8AoVdWGlKd
ODdsQp5DiShBF1goIZyAqbA54G0vgjdJSi69Las7AfiRpDPaAI4q5AfZfNx6
qQq7zc1tb3NQ25Li3mW59xt0Ey/pfpq3Yn2rKS+n1XcBWxmCJpT6H2EK57Jb
J7nRQmx5Q5MxPmpnT3BVJ8zSSAKsq2EZWkX8ns5TLrUHLW7U3EJ1GooiFErs
2kved0UPqu+QRo+8eNukgj335hprLJ8MfZ2vi9Ht1mE7JlTz8SvX7QThSBBf
pNdtfpSXNdvIOrMKFsm8TrXKS6lUC6a7L2msNpYGYzDCCqw1XLMaarL0W4lq
oulj+S94RPRA+QhobOnPAg4OEyFO54numMF6cjpwyuNBQp2tlZ3Hvfn9VlCe
C8aGAFWC3IHG9/GtAj5WgkoW0wtpOh9Y5snQnAGIViPp8AZMtUzw3Cfy9lc7
ipqvTtgqgUXz4+FFTZs5y+uXPyLDBe8JwadvuWSc/bUMhKSVQT/lvF4VAuzF
7ik/RTTEeMm1rN5jEDFRKKEXqZkguHL1qzREvkhhhINX6kYXUrdu2aS1AUky
IJa7lmImG2sWhv2QSjTTql0cUXTSj+BOCoPxdppqgcYwLwNOonG3gTyxgjXb
xoEHzUhwqRrPxgOfpeA5eNcGCoU27a2ouaZD3EbOvkT7CErUjCQqpqK44fi/
cspJzQdR/4GdUnnjc8CQ9FDHaTHcvr9U4Kh1MsaRv7ss4su+cgE4dcOs7tPo
F+mBxBVnDrQEbR8WsjcGPPuhR7APAROmPLthoEymXaNys2JuN98xeLZ2C6Vl
z6HPFxvayivCqAqy3kg043y0+0YFwWcD5nN0Ng6NOLqdUJ0IM7ea35gkzgtH
iRe3LYOv1A4clQ4YfMTWt7mIDccaXB6HqLVUxGVMQKgP4AXXoRqTljg9kzKi
Y3uZrfowNK/ZboQWyX271uDOARL928j1DSMnYgt6ZH5cZb6GnSuBQpFr3TR2
KZPh4pNa09X0NAZJNOcFfuwuxw45ipRSyiDK3mZkG7vhb47fA+/jo5gHFst5
mu1Bmt1ASGHt12dU72OGyos+dTTW2VDYSSynK0uye2d1CQxkgST4fQbfiMqp
XXk+lDmVcuS3J4k+l3zhyzyyczrBQnhpQOR42MhMCFrlmKxEZslIjlWXpZU4
457iaH9XVrwnwb1PKQBsjed8hE/bJyySj8PmJr/bt8MYAJiIxLLz6G0putAG
t7VYI3RsPbTjCCMU/N3Kt/v/KZY/QfHZvdSbeXv3WXTjq99q0FLVauBCRhW3
OT8DL4nYcVWaa2eJqQpZ8Z7sMeFcV2xzbT6BfouDOTEYK3MywTGRf/M/wRV4
L3snuJdTVNA3goQx3RcF8TSTSINnobRiNawrM9B9Rn9YwXRTimdf4JhYi0U4
9V1zP6aBAAaIF485zR68Q89PmyK8ZiAe5E3Wr+weyeqIOTGrJO0mO5XWweij
5q5No8s5W1UCBZy6IPoQ45V1OBwlV1zFkS3yLeAZqeHKE3Cvq3b18Nh6hmXY
zcdXOLxGSYcePF4P94dPff7/HoLJ4UEGXCd0T19ZM9txzhXAKpbGvVqVcfzc
zvK9QvhLaY9orcynuQmdOOhm717U5PuOrk7yyCxfVNIe4oVfxsFSIFdvpfC1
ZQmY1Cz6AhpOJuCP7Om8mrli7i0zNkmMCmU2KOpH3sqtcnxhpYoZMIPvRLxt
TOWRFVYqa6spcxjfEG2dPqanofPbddeQ7uvoS6iRbBZQ/zYn2DHcn3buwDgF
yq858z/Q8P7qAUCl9fZ7vPr+JYb3GKLkoVQvGKAPZym6evfLk8v+JXiUjE8/
pye33nR/JdpA9R5TIWkNcGOQfoyP6jaw3zhFHwzTrxByyrSLPpMvB+xR21Md
Bjd693p7DuNjgAHGXAJlafUaEJxqS6Zaq2dAR0uf7++fRzWNt5ht0KUvSumU
9vg/y+3SYHKd0+ZzokzOfkQHNOm1flArY6SOQu+7giPTHi7VpQckJrXHYcYn
KSuDpzVtjbPhzqH8lxdniaIJNWPg8WF2trWwXwqFHlpkGjmMPwO8nQk3AhNi
2vYVJBWLPG14v/XK4wz6OEnLClBMpXtq4gw4XdbSHpBHCTRrhnugOYrpG7Ox
e6nG735e/nhrZcNrfZ8CAXwWI1dIjkJgpHxAx6dhObJaaG0oyllIP4o/PPVZ
p+AWTazmZARGFf+wcykJ2n0KB50Jbn94YBcW1VpGD9xJOgS2/NHgD+/YUvfJ
ZvK3ZEoG1R19a9qjFs3u3GRLVG2TCbtOIDHjOVaDIEOkHh6+/mZEZ1XlYGCA
LtAF+2fpg7JzjcVCCxAdsx6lr+LNRfDQX+QPsb1hTw7Q1ArqtymSrRWesuaZ
dnjwJU64Hm8ABKuEGPFgR7DVBk8/0NOmQJ0NaATYrkw0UrrIceP4V7vQH9zS
cQLk2UyJkXWD4FQrud+IcqJkaCR43LIXpTxF4Na355Sif84TntHrPSwbKAg3
c8X5IgWU3egv7Qsjg6Ott5GgdgOye2DO8LI1K3KwNkkcDENGatd7Zd5DDc0B
DvgLFoLbb6qm1V/7siTjGWbURNfxJ0XH9EW76BOmsoA0CELzMcQLuJkWAp1L
iTKLl40C1nFq+oY/1lNxLYrDKrsl60OMP2oaoLAZyCVrwnewBgk8Oju8Ybrt
IEDixGuYt3bkFEJ+VPBaQn0vvDjyDSueMaDU33Dz792EwVdF7fYQa/33qf0g
eZiohpgeGiX9YbY9t1MWCxkXvG3vb5HQN6RnD8Rn+aZhzj6w2kZ+nH7WBcOf
ET3AoEUSqP2NM/hlsExLrUylek+8eDjScYyKW0WNpuf1pWTjFMsLlphPbbhp
FyTREw3u317Py6oBo4mMcDbCjDkAKSzBR26sWIlALNLzcWvgMdmeSD84UxYl
quDUFCpRTCYZeDBob+0aen4k5P7xTR90h4Bw1isnbjT8fi9YJY6gWmKWHoqh
eNq+doE0sA8bOT3IOeapfXIZoG0T9ev0l2buYIOeay0qG0QulVS8chUleCTL
j2O7xjaKjpmuD2H2uPwq5P6sCVRxAuhMD/5jX/GKTYh+eH6CxGX223a8RWbD
mx/NRU9UpenOA6BNQtb0wg3jrymqrsxPbgeHwk4GZ7Zb1dRhdHteYDdbamzY
sPjBOUdXHzAP2/0rJ3LrMkhyPRxnl/CnMloDS7CegZ+3/X294vJd+xhComUm
Z0x0TjJUKTiG53HROHnE9egC9HuKZILhtGRWta1EgL9VZUmN7DDuIhl+9xxG
1lz9rjCjY5EC3jUU+qs7XG1ULh0HlVrQpAC7lGfvewTWE6DDxOtpE7yu5VAV
XV8SLWm1pJfG7jE2wlHu0Sw4Q8u+dADQ7EfN8APTgWa9MJbT5fMXwQY/vGNJ
ghKzpuTj4LMtjcxq5hih5hhqJcjgSDe431TLk5f985OqqbQivPOKT0np+V6Y
MtJmB4k1OhB/FWGYLHl5X/SY0y52UZqhC45inoLxmu3ZC/sP3/7rzHjoY6LO
HGCqATyKp01s9KDRGqk2SikRjMOQPqYhuRCgV0nys39p0C6JN7cGwDVIlTgj
OVSJguAg89/5+Jy05LgFIJLcVlFrEkgpD2Qq1uS0gY3ojk4094wIGtRlyXMk
fcdacGrQpRBhm0aR6zRh1u67MSdoIPFNJ7jIH0G6wz24FN/6du+2mA1riZae
LUFTcJgq09a9oeyEewtQzv+xXwLEs/ToOXJ6+og16xdw+rDC7Mx398nLzVhi
3Jtyj0TJaimHNYNiOvNb3Whb/5ICFiTvuvgeZgJlMd+CMWI282ogYlrUeDiW
jkTdC3q4MADfjG+TGuy6TgNgC5Hl/qO/mOK1Ux0e5u6CFmhYO5YpKmuH1TpF
7n1FXZw6tPsC2hOHtFEekFJ9tZmdQhlfxyMvc4V9PQrR0U7C+0PZpPeO+fSa
WQici/hMmaOIRjwQ9FDiBoq1RsT8oFwUtS14eo8lDUT7StH3X1LECHXJWoNK
0dSkIHrWLuD2UsQbs5Y3WDIorEKpTIFzpASvQRF4uOM+iCRiQ7ZgorlIDA2R
i6N6V0TB81KR87DiMt3A2xd4lNyyp9ogg/yJW26QFpXTpzHCPGNRuuMgRBD4
98MY0touwnch3NqvqyaBbZpD7BEM/dv4c8jT2WfgStnPU0hMOIfNjpWZx7bg
raHlY8DRL09PTsU0XQU5RIH1DC6XD0WH0UK54XaK5ot7vo268M2i5R5oRaeG
LN23Iy+Ppp+h945uTLnWxk4ZZn2TYeyH3S2s0Y0C+gY3Yl9FGOquEL6iEa/h
HRWQnntk67XZ70R7XfeChgoC7bZ+Ov+0E+RIv/vJpNS6yCBiYDeajoA3qFuA
jWWH1jhX8uNki71qR59VcuyvcBDuQvH4AkZo5k34/khE0E1ULK3QSQdhYPN0
Qm7jL9unjHfoyG7p3higGLT+3xPFcg7iYVu1I8ftMvF8zDT3CvVCzunzgPp8
sI2+pYkMMekclZDBlCGdJ8OE5cpSUX5umUWQYm20pD3LDwx0BSCuNxjXRkHU
3pRaIFqi1rSGZof2p/Q35jGhA2QxYiho0HyvNw2goOaZFvwtSutHEAGDjpGM
jFltMr7uWCkygvwNBj/YktGW6mg+OQvcCJxqLn9Lafgiu0oz7CNusyzFr+E+
DDPIZpdSOFZhTtW6pYuSYhglN9shF8aufY6vqbKOLe6/kavVl/2fOXzI3ik/
DX0cZaVLoknHiqjsyc1xB7HocChA9mJXhjybBi4kUzARHPsIjKz/ziMMg8ZH
Q3IEMvvLhvi523kD+PerHLRwW0HDAyC+RrxssKjIEOeqnpynWgihhBOXwmmk
Jc4j4Rap8SbPtkbscvBvc1g9wU46g+hwId3OFJ9YVAyaNV1DPGDWGk1sGems
DJ8YmtcATNvDRocQXyrQDSzRt+4QqKl+sS8UtHB/Ben7bMeiuWA3huBfSV3V
pt5evFzUMHoHJWDmuiaDh6g4AVyZd+Cjm+B8Smyu+OvxDgfA/5MVBZ4yb3+P
dI07J9F1OvDLlTFDfuMNAWzZiJXsjsKzEmEqKK30FP4uKJYj/imnX0aLHLQs
vXsUSPX3XPvLGkb+TPRiRQ8d2L0ojYcAbUNMwkcLpLhWnKkirobA56qtdypb
XJZ9zptzGCySB3LMQVpPuQbN+wAi124nNr+xw8Jo5qunewtqi+BIB1VDvgvQ
cJP/KnSCiH2QUnZMIO+1QOZQrw0BHVdj11JHqfmt8V1VS7/lYcPuTwFTwMNf
VnKjPOgqT8iJf0x9LWt4zGZpoDAvs9FPbZrJ8QGBmr0g2Ft3xSfxvvn6iLOv
5e0soIcOZp4+GF2tZIIPU7VKGpXUhufJO86t9opORR/Yf0B380wCEBzpXYwm
2SE17G0goVpSG/TzjTXMJmtjdsmzPCuvn3mRw4gH9FalzWcOubJ9q8PjWdom
ZjVf2jvRLypd9MDVryB0hOPx/IUUH3WFdNxtc3YUBnrFTvroQdqb6ONKHhUY
+Fc8C1x5zoBAzvt8jeRJaiXqbjXLqR3gYbO2VAayGuZTdhrOFpxO45HxPMDb
QgqAccvVQCwJkO/vGQFB4N8Iwd0TY/qwYCWAPDf18+FFd5S9DeRRQlSHln0x
rdxMiSiKFDTyXbG/pDRyFE25Zpy42k4hGTrFCfmhuG+F/9wWAwaz2xAmXy1A
okOoVR0uzvfYSSIs2lkQQXeiOey+heu56LQS6C4VfT19EXdYMZ7iw/sW6qbB
6nKDSMfybKSNs1VsThGI/w3F7nZtiNnsUwasJjTgWqSig0faBr4YOG0kWYk7
+b4Bd5e8iNkOSjSly4F1g/Tcth8SbART90jXAP8oRV7b+q2RoEWjXHiI7DME
xUOxlYZ18naXSw3tNEGs3nLbXKlEQ5ly/GPnXI5Di8BfT50jJdzk9gvExNEa
KU1TO3if4LSEaFDVLk7kXx+U5S4qxVbJ3mww6nvvE9DKQ9dxjB5TRHgwqKXw
fkvoSnd+J8dTrUcL6V/qdooixyV0ZNNW9L+6wDH5j+duYEtaUprUpFlnSh3N
jtyo6AaDvDC/yOOogBxdyivkGyllzQ1PyuAb8AgxPjiBigX70UirboDl4RQM
FAHXn1xx8rATpTsBshCYtFedqdjolh7nwMXi5E+ASrgRGvgn3s9+g9Bcrw1P
ANnaikqIoLMZ64EIJ69ho/gbX3W1q2moRDjS0/RccUKiWSHK4i8iY46zzCtv
u6AwCKkgFGjYUQw+ZT0FViHfRJZPhCL2etBIMsATMzhoGIZ8qtT3VY1nbhQ1
OAknta1/G3TZzOxCypTFcOZ5sqGls9AxNPt3Woub1WTelCau6+98PfWA3S9N
ky7U5NaJD0kat+0+Ypuks8SipuqtNbwbtDe0NJEXo1YdcYjkcJexfaqsQFrm
vPQ8mIqmnXY6sr8qa7o77l+CTsffT8yWFnVl/pV4MFwWa1hyqR+NjuyxGLgD
MFMk0VVJo6ptUQfnP/IVFBZEip7f8jXLtJEjDgkPTSIHkESJkuwYpvOEicLu
P41xAufGYqQT1AdgG8f+Pl1Lwu2KRsU7fXVi7j6sjB9KySvFnFdCHPgQWZMq
9WhftZgNcehMDnQVm+M3om9amz4FyMryU7SED3bSrO+oWvrK8ZUmayGj+dq9
sbC525MfogBHAIb6eBJqn3m5JjJI0tFO65QfaK56yKMrvSVP6IbLNtNFImTh
0Bxmx/q8FUD3QWXB088ZAeYj83aH7T9kAr/hwwgcIBvrZu3Xu/dpVyibiXf8
Xoog51hDD+vttfKL/ONFDMrZQWFX6HpbTBo8W7g11YIiPzl9z/CWdEGAnPsX
mTuSqtZqqeQsAsuO5JrZ1UThwbkNOB7TOdOnlxMeXBkZ5RqEKzItEnJ0lEY/
vT8TXjeFkD6NWF04jlpx1xa2vDKYK8ntW9fDCa8IwQAlXDcgLkRTpFuPGdJB
MR5UCC47CyOLv7XuSRFVCC9tks/FpDnx3JXZqvPkW5jiej8tWJK/n866x3qW
58Zg5XztxF3/96MJYZyXD/DPD2GOaWMazu00IAdr4gNqzaJJ/iGqxlG83TsF
Hven7x2Q1GxTDohsBcuxUW2bRc329xkgTotQCT5XKTAi2KJiKsj7V8ZAJu7Q
GFdeGcxMa8OfamEeYUC//gDuNONCTIuHpO0b8XQmP8pG9iwXoT7q+zBB3HGN
QhxYVPUEkGwj5VSkc02Xl31T7oTJXjAsT2O0PpEYN2dVsuaiA9A92EHrCrqV
YBwUzdhNgNje4fCyrvKR41F+EpCzsNBWKqMC65+3qG/cRrOXCAneADBiyIN+
XK0Cp3h1cc2far23oq3rdnJP+lFuy4wcTXaWiwulQa+v6ty/AghTK/y+1FCY
bwbCm1Si8C4b3fA2ACfaiTnjYX72m7c+7y7Zd8O2ZZvsBb/PHkPooXf53O+y
KeKfGcxHi3UvDbqCjwE9PwrD+d5KIy+LlScUaPK9LBJSrjAyiuNj8vt518Ch
7XxGSWAbrIIZ4JmfTxIODbEM+ZT92E+nW9bkhWqNzbYalETBu66K5RwQmuN9
pVcYgmKDKIS09h0KVBr15pZJFlkpo9T/Jl5ycvMsvXFxJXWJlD6eyHAiAOMZ
moOog2SmOIEmkhLwtG6Exrsc339CTB2jLvD0j85Qe8Wibn+gHUOM5Y+FzuPk
oE3Cvmi5lYvQrFTOvoOefp8Tg8i4g75G0FwTi8jOjHgFzqADnUWi8qrpixLT
dQaWs9QQR54wJQ29DbHA1jIRy6E0ZVYhDT8ydgEGV74AhBiWXAexJjp/heRy
3jEnPfnsmYEGZwZFpv0eJgOEf+UMmGPQ3PGNaSXrpZVWnwWSo8lBp2Qb+qj7
ErAo+zxkINSgNuzVyZfSJolQOTpe8NrimZShXAmvVhE07TLzSeYnc1DVaod0
UtkCqNz+sgkpdi9MegPAszWmGTdKwkcagoZj+ZYVXEI7NWNbs4BfNCNntHvo
VmPDmQPk4So0GaXuolFGdonVQP4906X7nqPi3w3KCNRtjmfsrDiUeSyp28Xg
F6mCztvQJgN27yOmfn7j4Xhs+ZBeYqiNP8EAAM27cn6qTapdkOc09RxhB3Ic
jDqNetOM4cWHqd9rV2E2xuIQR1LdC9nLHEU7ioPmu51/2R2ljdPHWlp6Rx/C
kAsYxj2rK3Fj7momSmEXhgpbpjVx8ArJkuGAP0KY4GNjR8+yP3vDf6E5aXzv
dX6nsWCE/ffkSC/3lYqbMWRMOiHNgqtDgR5avpCgItgCOrUH8BI3esrTYwsZ
HaHSgapU6ovxWRE2qEI7Qt74q3Xk+3sGRlDcIzPR43E5dH0knW45ms2ndS31
sZwaNhBOrrdC+zI7/7DRItkZAp7Ehx05blwG82FMpzkyVF4ePtqeFiKNBEF4
OlEwz2fonyuJvckUOe+z+ZLQbdZP2kYLaEYXxPeZCtKpQA1iTmV9oAMbn8tS
F/Ztne3aEvLUz7yZfH0WQhslJF/qUQcaZ9GZ/vvI/ChrapUtpHhKz0Icbm95
xhtjvhqPUWvGHGPi5yqNIRzVZxf9ut04NAwo7Ex6AgjRS8imVqOZm45eAibS
iHNygooD/rNlWKZ+qmypk9z9lAtHhcN6EcXCL1bHQBj7GdYmF7VWCqfPMcUb
VzhpgEROK4O85LHx9I5a1tY8QRg8NrzTWiz47YnudI0MaIGS0tJDunHiAhj5
OFEKGOb3dSKUQquHV10N0p9bOiCyn/1kZgt9YZg37YTnLrXMZcXydty7sodu
iOxKrnbT0TVVu/Zp8/0UAqf/GDy0Sq2hYI38tTEV/y7lvqujE1pMgVQKD85z
Jt1BOkSWmwvQtrXWaB5+MfNzeUF9g6s7iHb50oQJdyJGNtl6D1nkF5jptMZ5
8KFONvQHDa2TeS0SoGjmHxd/CuH5m+k3U9d+PzFETqRc+6QQPa41tic25qLY
cSF5WBhezhwKiUE9r9c2A7xj9pmEP/KSoZ0V74jUqAsaU9dh61RumnU4+6Z4
8KBL1aay/GFKj9Lfbvgv7Yob4xqgIqVzlne9ihx3f3LrUr/Zk83+h/rTrPiN
x9flqbCFgClcyJRzOac6iSDxXSGKLkfipa5tGf/weXSVX2i5u0Ga5gVXsg7E
AQbaNrL0/wUrau0LF0SvBxWEIrXXLJSrtUkcUw9lTMnh7L99JGH4i34w+jL+
MaRhvl7XJFIChrlgONA9cJ8GzlLIvu/mzL2Wn/NHiu1TaUD5yiDWzHSyYXaQ
A5PZHQA9496YoEa6P5dERgPZavr/CgLNxPn5dkxemWjtcY5JpGcyBiveTaPp
Qg3/hifxq+GoBJeME0+yzz8aHsrMRPFExs4E6xZ+TbKVV8jwxuX0gA8NENrw
U3EZMVaZtQOV7xWduWYhC87hjffHjbs/PnB9YseO2rRvfwfpp+AJZJ+r6su0
p6C5n/95vRTHT5M+IcSNZgqxuf+GCKHeS2Y8RuhLgnEBr4RI30UULqFZrFfH
eTUQj3WgXWiJQ9aNna4EgoWhHzXGGKLBiuq5gVVVXSaWx5dxvFlSYwtvsPbJ
44NrA7q4MB3XjJAzcNBpnogTou5nwjBRmen7/asc6iXO3zWgftvShD2qA0I2
MGdXgGR1OR/qocgpFloJn1QUWxvJVwznAlYtWMfqG/A6O6oH26IzpuD9Q2x+
9OY0VBHZxP+WudPsS52vnvnCvxzaJUb3Md3a3mGVI4OqmfPMOQ67SF0Xjrtj
qGwiFlcVLX70SjjGabzV9VaY90vAMTdV+m8Q93ZI3XHo5UdPNLgPyEvEXHYH
cbEetXCsYb5WBrhYgbCaKn9hHlXU3/PzJ30IfDeIYsHw4r30EZplUM3ssYSB
GDhnU0RyotZcnfi+lDCNfQoqP3On3hsApXbI+hHhWEHAGflZzCRj24GV9k+2
KB9LzPINgY58K566oNLscSA/XTTPMz8cy/U3piBQU3syGvIh7Sd/GemndYeu
ZK2wNGnx0bUqRxWOdpMm4G25zwKxGwldYkwPBD6cJ5vbhwa481PNvOQumIaG
QiiZoRPqIjSj9Pgmm4MueAn/uQ4TWgyTotC9hc3uG9UG75pj3ydiZ0EikDnV
xaELF/g0J/LARI0epiB4ZaMD8VvkGL0Ij9mSCSQOvkGEiRcdtCWZosSdLG/2
q47f46JkWLEFO0c/oG8lFduvIIPlev18/2qSYPcCMNzHXD15Nke4k2d3gshx
ViFr96ItcHyJoilrgIkF6nVMxHJRKO9XOqGzdYNx/KSoNW48e46Fww5LQ36T
zlUwh437qycBTJXGOFALXApqgLZmXFiUGTWhfLN70GfsrczmMfDfZqAlwpHQ
Ghgnt/E2HrXSX1pjdsT5N1J2bjSeX9tRVHfWP04XfgP/ddHjf5Q3opy/dX5T
BMgGeoxL0aBebslv6ft6CQ3j2N2E/fWFK/RMG3k5wQka9ZEvasVRWUhHfahh
3IZNCcRy5PD09jea2jwQwGLzkaQGEtxokAM4rVeG8+wHhElx7IKfxOQSqDLQ
WTmIlgkzb0tQKFY8ptP6CKY+jlRePBfjMpCZUSXjMcgzMQm+C88GRKL+f9mU
e+lB8+Y1cQ0gKtobiIJifSoFj36TdY0u9zV/qgwTldQE2pZ0FFDamlN+gz6c
EtVYs8n5vqMYwkDzgSqDh/87t88kK9qWJarRdsrEvn+J9QsB885z08zmlZg8
FEiSJvcRtUjXVx3uB3f5xM2TN6gRcfgk1PlqXLE1ZUS5CwMm1BmNAQYL8cVS
8QhYi6Iuvg9TPS7iquumq20Axelo8LghjXVeMCcZCucG+3P08PdgE49/b9xJ
iru0RJULArqtuscZ6KIzlN4LVxX3qSJxvw9DyyJ7CfCYCk1+k/9djkHsHKDZ
oTQPumwazEhzB20qtZ1eoNJn4SR93GZwEXckvhvLv5cngTlqznkSUWPLABsc
lYsA9wyTyijTXig4/y4uSbILycgEOLRJgWfcsnPVuTSZp6vjK9JiEa1Ae3tt
xUSQ6WJA6Eba/083cRWdxS84fCNNL6emijVjmC5sXmaEJl3IuT4S+gVpq1Cd
T9Ec0lGdBxek6+rAtYtay48rMN1MIROpPmvuPGJe3FWg2dDhUFa3yAK0dviD
i97GSVl2gmp/hb+ZEU+6ajv8FDwcqarJF+phfXq8DO1Pn2fe4YHSc14YpM8b
dW2+Hf7tfbFKftjCR6l7yFBKutd9r7krnyOrPRT+Ad05UgZuSkVkn+5Mk+SD
zGOY5znxVX3X5zBqlb55vqBOtLdhN8W4q7VkhiBunU2HbVOnCmFOAPyt7efe
aECniKRgwtPTbrQ8XHeZmjK8CSnlysT5EVGfT29OJlinwwVv9D55mNwp7jkb
qwFw2KK0Xd/WViGaVDoVvOy//mXmlmahJKCE7aw3iGg4T58xSDQXkXOt3t3C
2fWXZblYaH9hqKEWpI29FjnMn+pTr2/cR+kS+ckGP2PkRF2hYhxD39wKqWy5
KvBNnyIbImJa4sgz7U9kYpqFMJ0wzyQmgLek+bLCktZqzwx5R68rDyaeuGPU
K9zCFk02kLnw2GVTb259IeoKcrtN8wh/G/kPKylL3E5fYnJrAiURmTB4kFEu
mtD1bJqQPa4gKEyztb617FTOD3JHpx/nnBv+RcktGouzA54VIGqoJ2Vj5TnP
ARpr4qnjZAtC/Zrc6SmfNJeHQegfKNkSKR63X2L58JeuePm3u7oZ2Z4BiTz5
Fr9iOZ+WPS3ERvVC9mvMrf8VwNJO4rSHD4w71sJwIyNtIMj8N60vc4FwhfZe
NOTRQhyPZx1xCTVDN84F251VGLMXwCfnZGrd5Pvz96I/1AX7FSYrx+vBQnP7
GIXhZywHbSaPLoyKPl9ZU+lmDO6b890+Cj5vlF016bicrq3bJ32/vPs9tG00
trXeA4ezRNBUuHe5M/wrOfv8OiQrD6R8+A1ytW0CLudgnYALps2uVCJQzmEu
/31/9/y7iE9fD0ctX9USPGKwOpiUFpR2mcnmHRXNa1N13LxVr75z6cEHZk5D
K1yBXDe7Ezwyq3zl9mh4Rwtqe6X7RtZOXSj4eLKxMFGsCFXFQrm5OtNr0r4s
Q6j10OM/qHjtsssZ5ND8YwbQKW5AwgcQTibOsUNap1Tz1xnv7ZbmWicORYTK
MAnfmb+41v6mgOGuf0Q/o9xH9C37ZsJYavmV2HYw0jPRY8kMPRTjTdh9WOLg
oWspe8OdJJkhnyuIexMj3X3yifhlTX6CCDW8Qng+v57YdUxUpFu2K6Og7JIX
d4Ro56Oh3l3h5EtOPV/dJgsPFpgSNkjyHtrDDNR0KU+pUpe7m8uIWs4QlHE0
k9rAE7LEf96uM9cPiLdpxPBm9/dsZX0Z8L687G8vhrP5wV3pw57N0UJj6xlp
DzyH+epbUbGjQZhqdA4rdtrIaVvNgcuw6DykAFejxf9wp8lxXQip3RRKSs8i
x2Oi9Ca97IgOKffGUB8pV2PvHo+YznuR0E+EOT270+mdqMupiQtWeajyg6Zk
XBA0WnHfUU3TSWBFWY1j8qitjkdPu4NpzcjVY+4356U8MXfcZPG2t0bH/JSU
QE0bmaNty1ajOWza+f3uCKIaK4WMi8N9a9dDpm0NPWQ0E4J8Yz+Uq7MtLdXH
qYcidvp4f3z9sUkx/wqaIUpxIzuOm5h0P2Jj+bd5FYPUAjPITsxjRzVRdDsK
L+RJxKk6qO19AKlQBBVjL3ONf4+mjhaf1IIP7Fac35SwY3Gd8LjYFipun4jD
fdMt94y60TsshFAexcYD9Dvf9hOhp18+nzBxnn3++pMW6WKZBmqlgZqj+lpg
bm2UQ4etwsTH258rcmz7gfq8EG1j5iBmBmyXy4G++afFkQKNu3xcN285LZCf
yZMHbltUM9o9MQInUjT3KhDSTeIya2jXkbYS8wtLoCZQ5W38rP0U3fHnxa/5
HH32ExHwETQmFKeSDgm/DgpzVzWQoXeupHtUD4nMMinRcnWZNmJHnNytDuT0
Y8eWnKJY6usB+bnMtyRL5amMt7hZFUsp4iRzh/CkD0hgym85M5sOdABRHNGh
5bCDEpWZ0DzbdD63XWcNBGIBUwuUSRg2nmpvBaApvGyQzxHi1zHOr3kC2BEr
7q3Ac3keuuYqBSlgF5srQqskz06TwgotVTxJgyIJu7PRdfcc50IVm0KxTplT
VnDdoy6PxQF70kFGrKjr5W1f3lgLS33wWILFnyHuVYi/xB1OJWmuwYt3cQPi
b3stau//8FnDB3ALkuMW7y1DS/y1Z67eAISo2uGlLi9qLLb4BtHCJ5Zvl+eZ
YGNkd0r2OYvRfyNArILctLX9derZ4i7fMetEWoAnGlmloDfKBxLCTj037NUd
ROyBTzL9I5NeHKuuimesNVg4HE7OOCp/BTSGP71Ti0E7kyOBM6RobKrZjvkP
JQlz5JEO4TfKznOAiyBt57VLSUuGN9XmFNHC+ViL2zJL2V7cadNjySDwS/41
JmHPtEs20N25PLsW7EEa2y95UQQChIQ7X/hAq8uRF4SU9EAfPvlZbr6qoG/S
7Ub23dyb5u6jAyqGwconwYG6NwU6uJ6gJQ5IeZWrksfV/kJzZuV2fz5xtM7/
g5Sn99N5Y5Q98z0kTxmSWCUnudwCEfFiAgn564T3yR3+L/mmnqI4WqbiZ7ho
xPQ811ZabEsqf3W2vVK/JY8b5icfZ49RMPrwXY5f4T3Cb83G8Stf1z7Fcz9r
KFMwfcZ1ensEEvTJDn2RzwHoSk9BJ08b4lW8dGJrQnGvpqIiGbPCK9OgdJby
zmxekmiy1obh/9Gg27/7XEiVsoeF/o7pKIsi3/ls9Qu8zSmXpQ2H1jhnk/Sf
Nk1dold8ra9DmYaT93DZkHXVBlW7IuXf7ypW8YOQMf6FWrZYTv5ppW9h/hhe
KhNV+GPi0/uEECDHmgnTBiOaXwsVOyb9bnjuNCG/3jHOcdAcoOZmIazj9VOb
/vojcg3nZDuVEd0ow736sjfgHOXHHUFxQv4LVxsRz2F2s+rdqoisQlaXFWvU
oQhjfv6ow8X7xng9owR+4LRlJeysvTp1z6r+X7Vrw7uSK76W7/PMgskgcTG3
7dFkUNo93FOpj5S3Goqq21F5N6WmseDuzzsjUQiwH2skY1zOUwevZuuvNhpH
wMCLJpGdD69SaXPYj3r6HomUpaULszuEdxZ0eg4iyHAtZzJpdd+SiBN4GFYJ
qTVnRUHO/JBqYkSvK9rjz5DiVoq3phxTdpcLw8hx/FB2vrkzRECwDpLJ3cFE
FDlU/ZmIDRwU2sX1Qy2ckABoWr8EkuaY/7KmmMwSBxMR2CHGShEEDi7q8Yvn
upEHNKuODOlCpKRNxdnrN4akXb1BFIiqo37Ac8JSHPoIwO27gKWrxoZDE+F7
wbW5fRnsLjRLtik0zHNRQLxeGEvBkVjidadOgTwidKi5WgC9fEAOROKF+1WO
I1A2T+jUIYrhHmt+YAHni/iKf5KYWM2Xfm9k4WNw+VDwqmKz9Oo0M4F7vhZz
opYS/+9eUlfVM8MEIjl+YSRWyw3gaDN10DYZEjP3vRiohZgD92ujsWlXy4U7
LBpCU/5V8SoDuSJZAx4LUJEPfiYdxVH2saTUi6FAUOkQbphVnErkp2M+OrJB
mzmfb2L1u+n5AQjof/mis8/Ft6cdvdMnmdHtKGcuId5Fupa7aq6gJBfDQoij
B7N37lOqEvhbPZJOC7ouMvTOTcwdE9eQyNSpgikblOuVhlY/w76kW4cuUGu0
ADEfjbBWeYJ3dNEabmk1fL4qdVm8VS60u0LZ+VtPmnjmvIwZiXvrKbfFWkBr
IMCO88esmLWhk7N1mdrpCVzAfJvS97kZ44ddh3xrBUjguz6x4jIZOTxdx3LE
pj3i+hDlfhfcV/kEpwiDtwZ3WX/VvkZSk1T6xRXFAPsyQPToE2begX8x8aBJ
g73cbvYy5sViBiVmvAQC4yxCD0jRdOw6gW00tFvHK3pzkslsRV6JL7UFQsEf
0ekrdqXOSKVHUcoSZmed0LrY4OE4+P4yPrePXfJfZ36Gkfw4oSyqC8XuRf4X
eEg73hmRpcm2WviGvVDJiPPqZ4zyHNktTPpeSn27CfExn5QN3KBbeagn3rj4
dEDU/s/Bc/sUQQZjWEvC3Z6AgokzFurkuzBIUXtlcXs7EPoWlMWPHx3TNgvO
rN/UuEkHQRSszwArMBPSbxmSybpMr/MGteajDOOmoKsnnJpDvp1JLBLH2/zh
cYeepp3KSD9fwoHnK/n5x7jJUiCf7V/VLI0ukbcH2rChRmvOlQ8876PC5owY
O7VnCD2R+6OMy+y47ULoOZ+1T6dzri/tmtmh1wWx13fwtUAN7WjcFyQmIlwQ
koBw+fQ/zd2ilvh8n0ue135TEFGlaKnVFMN70My7mNpuGLGEeR6mgdX5vOsk
nMjinj6jjQbFo1TeUmMtVgWB2BIyeTUt8XziFSKj/JEsxMCQfKZuA1nbL64y
rQ8TShmIXmJhycJBXtbbOQ48ROyiowd1CPbqoKm0xI8rV0YxJ1WsudhEmqv2
2Ak+l38EhaaTwCtUFTdWfZ5Awc834IhkJ1BflVvGVR/usp8BpmmYR3egrlju
whQU52tHmPmkKNfD67BgnRtADoeGIWinalpR0AYguZIuws2kcF0Jf6c6rsdL
qD5Ehrcxmzp7M0nAdX0abem2Uloorlx68KDBT2WZt7xahsyK/1esipIfOVrP
YbPa7osCJ7fDPjYvQKdJexT2Pj4rGmB//14e06t9N43+ob4kuw6nCaytQ1MA
IKEd5PqZL93tTuripf5UVkHqEesx+D1aP1VzC7utzVoFguJHwLW726pUGaOS
0qfQNOJz0nkPdljalOUJHG2y6lCA+wHEvHhWSPT3iSEt2iMC+IDCDDdQ/fAO
yc/xXWo5SLx40/stcuocD5X6i3sJhcJb58M3N/FjCEFozxuQlKBEFZZZ2Cot
JUl5PVv1oxD+9OlLczFpgqKTDV2yQzsOugri7P/cf+UhjtqCatwyurNOFYkF
ds8w/rOF4+7tEapGV0iqrqcplIwh23/iEG6Y2BMJJv9Fqb1yG7mKtmWFuMV0
OR01xLWIX2jEo9fqlxPf0IfiW8RbMH1QK5L0mDeBOYllx1gfLs96P8a0ZG+z
Vfq/1VK8ZoEA4jqX9QFu2a3AYfr4xJJ4WsQ9O+bBRoAALtMwgjD1nBXwJdz7
Pk/o2RMuLM6+BXYUVl7kCi9NVVeBGlnmtg4veMkrEGKUII3+6pmjtllD8Tkz
pWUCD9XsdXLnk4NMxrSfNL/eJmEosNWqQhxprD8lAeIWgLz6GIxFjB19ofVA
UMCUbTEtPff0eXHmuXJvRnuDmzgErRpD+w6E41C3uGrLHg/P4onBrtu/J+vl
trDasTdXTmNCvsYQffeojgIR3D5L3ZPB3BIzW8kCsacjTHJzllY6T+r8SXHV
YgiXvyYz2gN5ALMnwCOF7D1l6nepy+kum2KwZxt0Re2T63cMgmNPhdDUEQKu
8EUFofpj0XBbCCb93CLwcjly8fWWSM3DW0IKTymmFrxhjUGJNSXnmLfPTrQr
lYkT2IgZfIMvdvJYd+WIdhxFOAS3w1sGzQJp2joRlcttgB4mGHj/uhUWJaj+
jW/hbDLwY4VafGgNCacjdD7mu7WyveOUZgHp8AWaMFahul9T8pym5M8YayCO
vgcQYSuxY0ajVUmWGYIWcqiChcVY+yM8oURnMSgskhk82OJwr5T+/88VSI81
Se7tSRui00AanOPbTD+bI/1rRZTpC3fY7d/2WZLJgN3VhpQKZ6ePlQ5nD2vJ
o0lBW4SSLD9qWqWVUwQH9TrHa8cMJmNcdVRJNpVYKq64JSA8TP+e1cpNKAI1
DMWsBhSlyoqRlLDgI6IlnSzzuydL33eofAsXhrknIqWdd1Io5TeRAWQD02y4
p1K4G1sUUa6HoeTa/A95lZGVgqlAQV7akyTcZjt/w/QKYq3kt1Sv9w2V2tG+
hAXbE9LSjSTy8JJB3hrv0alituaStdZG77QzDxdHY+Z1O10CRSOKIfn6ODo+
XG8H2wtGK+Qtih1Twka1OtTwU0MijhCLOESCKN1aOg9o0DO2JCwZD6+czggJ
jbHjzqPMPfA4OzjhnxhxpH9xIR8Gq/cWASDmtXPC/Eklx+L8J9VMDXxRnPbw
ikkxqGfj3JlfVpQDEu/uXkYi/DZvayu4/HerfxmcyIaEV9VdpymX1gbCmcw1
9o2xQDkrCgsEwcVugFN0RnIrDExQHp2yKHdm0Eb36KozUvLuoA5yvsGagPuQ
bTphBvaNCRcTPcKExxElnymO/9WNEljqD89K68zidTfxpIpsY3wk7tc9Uflu
2coFmqsnKMjUcwUYM2Y27ETELnGch4SEPyjckB3QBCtkW0ydES/8pKzE4g72
nnqQCPJr/Fg+vNmOagKhZeU0+6MT8sIolGOUlhjyJST5m1dIZDfu2z9sAsLU
usN5Kh+66743H4mZTX+95PGtR3WYbNsvHTHiXZhL2NAsG05ynKC968hXXMFo
Al7epM/JmBxTuC9HC4PvDNqfTLlQX2CxWHq8WgqufxDBTQu3y7usG1cNrfwG
5DxSHHu4nS0E2S/NbXsKZeZeznOrjpL/eW3MwjQOMMQNjloerILrbVrn/nAz
+LS3MxczE0k38UhJl6U7DDBDZJMugLet2dsYN+Xzuqm8r1um3PT35PmSJgzL
OhLEbrWEDEYAubfrepEeVICUjWxTBc49Y94Y8S+QbYvA82hqdYOKiHq82hjk
OPCpaSTHiGf2GeIIJ9hjLTrVVTQiFJ5+IqpsPFzi2wehsYtSpCv1szNxtQaa
OB7HWwY/mprG7UMLML3kUnZVERkeDglb0s3c5JnOGhbzPCZwK2WbN6XOmQbt
XmpbakJu630NsyMJbJ1uTndWQw4Ab5XB/IwFpYsImE9B0syP9sXJZlus6q3j
amOtIAud+PLqErR4Y4a1g4ZJVcr+kwpWMjXqyAXMDDn7DJ0NZgVqNGaHFt96
sNLiqcXC+gmh9Ycz5lwXKMVG8GL+4H8Xh5G5GvTJNGS+UHYKgjHpb8l4qYdt
FmfUSHMDKepVf5/22WljcGV+WwQcT+64x35zZamBwRt1lg7il81ZLd6PG62T
WNmQNDw3QkKzVekhxerxPHce0/8ZI/TL/LQUWG7RonzTkQI2KNLwwHxrccTj
579Zqer0bPz6YIDkA4BJHgGmob+gze8DhVgTSBf5Q8JjKwMfdC0MaYWDCrkQ
GJD0LWbcsh6gPk4WZPmKd9KP7QYf7uDaIzGxTpWTqXU8vV8evbxIzCsSPJ64
r22kI4AGikPUL4UYkfZLpbqEDcX/jf91DuOcm+n/HApI45W6bGCiAP9w4SMA
b3QcqKAaoGTx0z0gG44U0V9jU/5A2xiPVXI5rMI0pvqX1XWr70G/imJ1fyYC
m0zlZG7oO+UdmyofVFGWBZhncBCfNzybaRB5Ry72JeO+01e+4jeIGkxqU1hk
66+Bbus2kM/aRNCx3/E303YK4dmnZ+5nbELQlOHPKU+tdUItbdcQcXt4Dal8
BnGTgB5ZrvomgJZJsboCFbcr1qnzJzlyJ+AMCTSUoI6EDnkmBUqEhDKnzgmv
efpJ+ASRBt2sVfFGZ1yZYJUHvksjI4PH1jiCYiAcE2adk1VHN4UBNkCYTUie
U531UTIMQ2d2fpIptuDkVLqLV+EUkMPdMoGUv0mHRiMbOwVij89qJya0jKaw
vwjaNjUV0ni4UA07qwj/eJjA/uRV8qGwm2jr8CrVaGCy03ZkS0Gw3PgT3Rka
0aNtJsKMX/YTFJYUhn14J+bMnTA7U5Ek7fpUdmvJUCeDHAxDbpBXADYPiL59
EeI79GFQKC9gFmqlFmIcI1CPH4eYvvwANeUnyQXAf7JMWcqeSXS66Uobu3j8
Nk4NnlbfbTS/11YVn4WoLgo/IoGTWRfO1U47/D9Nq9VbKZA6gxPZEjtK6d4K
b7VM37gpRrlCTZKFEDcXk2upt9Si9Q5mAH+bcKXD8xd50Ka+kOA+tr972e8F
bfxHv57HZjztA/tNh+IHe/LcdnYw2TAcc/X9NbaIoD2FHxUXA1+tbyEZ1ZQx
Iv4cSBpQSLZk4+yyQlIk4X+eJ9+yLnqosCe1L6vp+WcWcg7yRA9r6GAVoUob
IObLYPwSRJxRfjVxURNok8knUqmBtxnmX3SksYA16T80JFENU6zsjoBgIsJO
Fs2MBH8xkuQ1T7KB5JQBZeO9Jdo9UvVruMkxO+l5GDCy52r/lN8cYjr/WSXs
+TFt70LLXUNhMHrii2a6IZts2p9BFQlSLHVpsLWkauORFY5MohKmXU0ArIrI
3O/71eU5jCl21aDfDpjVAn4xDfGq7D3R9L/SEiItG1o32ATpQlYZGHagYp4d
lTpbUWUwH4UhHlbXMHGBV36H9HaSRgWTKklSZ02eLZtaVb02Nm3KEbv/5T2K
VUF+F65splxu00OQtvQjb2TVzc20+1ZOXbmMhc1t3sXQnHo4dGthceeXKKwB
KM1DDE0hltmU4c0ID3ELOq1m7MFRXjnlifXiae+4R0Xahp1nDN66WIO+ptx/
O7V5Pd2N62XlQ+DD+4BQKlBiuRtZshT1KkiIUX37uj+SPISVK4yPyNmci6sM
foutWHk8cl3A8CKH2YQv0hD/Fivi6Dyhr8KzE/Fb7mllDqwRKTh1gc/6JN/J
cC6khBeeNx5iN5BzZZ3LNYFpBG91Ys7YJ07ebkRQLieQdyXNBP0gUssXSN9u
LaAnrv8C3wTxjGlhpnne8qR0QhKJEOm8z8iKTmJEZZESbct6Z4I94DvZKXg0
Zcxd/Dz8+apn1ipEkQDoHq2dnpkMSOptu3zriDdGejruRuhdYDudzKYDSFGy
1yaV19eEEcy4gir+pEw/JQW3PcLzBg6w30cMcq7pPTNA5dBFKAJ1OqpEGzXS
ZFxHl8Hqs4NiziFIPFAnzKTNRPsKs+7/hAuTIz90Uc0UZ11Ui8/3mCTieUC9
LbTtXLsuDT1fVc8rYlP6OAs8zzcHbX97CSgVDUDi0i/esBnPrWq2d6rNCT44
2lfJ1oyFQvEfwiuI3t8drgmPmVv3XHikUkTxEKE9+XS6lxwvUXwhvRj2P7O9
SfGwE/6yO2m7lHOU4us6HBkW6VrrsVfeVApzAyi+YecIUhb3Uh34Apw0zD/w
Xe6M6gwGlgGdirXyNfaueFta6NQk9spyAfL8OhMHd+Z6dbW8LhpvXBfA5p1T
bJgXkL6WgdkFXgxe17PRDY/wQ2n8e5jsUVc1salFTDlTttFKd9Xr1OucNCt1
zD74ns2BJ4dbq2SrKh3jjVcgTq+XpZ0GMOqj2UlaG3FiAL+kunZhnhwgUsAR
KCsyM7ReWAh+D95pTQfRYaH5s5DU7P+cwteGd86pyT26GVaY5ItrbkVgUjus
OOywJRyh0VEJXEpWrfunyzgQzCJHMweQqYO4BSW5vAeDBl5n1Kq0gR79gdVz
3QuJdXAZnWsk1o3JLt+piI7+/cXJfB4e/oxIOPJs/gJJO5pGaliBEGpBWymO
NIj58hxKOxSzlHuRQtyMSaDq/4/3N5JMAy0s5bxdyCjm3FsgTkFJl8BSaHi6
ANro42QfqhDwAiT9rGoUIvLoqMZr0UnVGtKNtqEF4FeVE33KsJLtPOC2XhjG
r+UmkQ637teY2POPAxRSjvkNgaIvEJARL9tNavVmMP824GdWESUNpPdx8RKf
Yeyb00+WCujyRiZcLrT6lmcdA8kn/rObU9lrVdoUfjuuRqYHrnJYPBXbOjTX
mgRMQvnOVvVRlDiDlmGzqhQOYcC8fFHwJ8C5k08g0F8pfGU2UUR+EOBJZ68D
xHHwB7jr0ZAblS8IeEIBJLE0IlLQjrD7Ls1UL7nh1nVXYsdP1y88NHoQMqbx
LMtr3rtmRUsTpiUsyvGvtCcZcf02BSJFA3ZCxUe0zOCnCHRQYfVMP9WzyXdl
JV4+53rrQ0RzZHSDov++OiRJpP5wwUUHynJLoOXjIsvApM4eeDwnP/uXSwvc
A5obMJAdD63yH/L4WnhqR6r0i+wdySp1X5Th7FZBTEiBrvouKtReMvx+wQIy
WBULNvbAE0LKkdaNo45HkAFb2QZENcTBxNrR/Fvdf+haorBQvGJNm38oqKNJ
viUbYKL76VW+a98XVe1i3+bNvlYGlwVSU4qcKGVUrGN1M10KqX+A3DEebMuU
VWOw6wmBGSlxruHzXleAI/udXwaA0YAvCR3cydt7mVJNHWQqfy9CCh2v65lw
0wTn+Au0WlRVCU7o+ccROYO/3u5fKi7MjF/MxluHJUjPfip28jQjJOL6//Z7
ZDjRE1DRlQnWpvxonlLseV8OFB05eWgWYKtMZktu4JFPQNuL7Y1LiXaCZf3g
vmjQYIMfskRg/Q/8fNRhywnrR2TZFk5s9pCX4UUf95O27VYZPQ20PQ/Nf/vD
LgDEE3SIJRpULCC6+xRH7J3l/rI6/+QRqfOIPDsP/0v8qWKXTBePnWjyIp8f
/wHhhevFLtdxzsvtxW34OzoGTambaHhzfk87HpR/cXBNofz53otCLbTGnfYh
PFuhFIB0XwgXWizWiWssB6oN77bt/zlV1E79QThv4nDIxzb/URkSyrpVoAwR
BPtQaf1cC00CeRzTSIAsFtjwpmA28N6xaXt/yQPejiXN/8OxDnicxMCpoyU4
MFV8OzSAWP5QPIAd8XIaM+Dnq6huyW3//zeLPnwL3ogzKRv+MQf02uYKQ8VU
s3niP84YwgrGaTgzjqeS88HC3KVwsZlDZYGZ33DeLWYva+cjFb6AhZf4smTy
cTc/su9oEvJnbanhYF67MsxrAkDs90UWuZQzpamrUnOFLAne821rzEDcB27A
UbZg3UDMM3iXYqk91xPp7HkHDyLNQ503F/mxzcQNvwytkHGqMeUF0gcrnKgU
Gs2vkFs5kA5dWooxg0yOgtGusGTovgPe4CcT9E9CJD+P3LKR3fyYdKeQqUEY
cJmOX1iMcZgqzWS/PLabRct9K2mGEpJySk1T31mki1dkH8ssIqYP2+0hH15t
NwyVSGJ0S7I+GfXQslbl3lRX0xQ04udZFrGGo6vUpVHKR4hDy43Wi8ju/FF0
VLLGlLCEqFBcaoE4NOMCq9js/CBh5Awkr8rttRwWpJhdFjQ1M6jbmiV8Snap
aHLglVpwOv0frbObDykbsU0bR5x3ATbPk15PNiNvX2jhGwRk8feuM+tCp4wv
59B/KkeZpHA7E+hnEdOL7baSqiQ9AD1VD41foVmFrhB3r0KGjuoApYxeBT5j
XETUzuCMo54ESZvQQKT8Q6GIx9sQ7WSNWJ0CdT2GF8IssYRhzWPtpCQutRM0
Em6g9pAnBdt+o3RE427PRBNLPgUSVbu3KOw1H5zgqEZwnrwq1Wh/JzWPEuNO
SqT5VymYyU7fCpMb3VosVCn2KvPdWDOcxOs3tXk1Owsxp+51Figm51JuDQ/m
0JwIzFfg/AZBZKZ0Q/p+F0NYzAJC+hAs59qUWIFcY9rHuFwRwO3VY/ZL43Dz
gyIA0ZWKAI/6lEWgqrqZ43/AQ9egedHx1SB1sSrMTqtP5xiXtshvKhOgxrDv
5CdHvWzBKrqb7TVxdqRIBN218LwqFoFziAIJ0BN8G6bc3NvJECPlZVeLBNSu
3bFRC/EYr283dYfHZJnh8s0ZYjMouZjr0MCJUomiQ49mig9gjbKet8+SBCRT
WHFOLC8XeOc9bCzgXBqq21cY13Qv75xnA6MURdNNk7JhrO1S2G37y5sKsjXA
mRJ9Uuh4tS6DvEKA81m12E+O9ZK9tBT+lmAR3F15IaXCb9Pjy56LY2+1zD2p
q0/YsrmDoW7w+kyGrCiMRZTAPUmwpeg/JeY46Nab0VPKARCqi6TcrmRNatFc
1A6LmZnLH4qRa5Gzk4nMYJBEbOzoVkhEjDA9YKrJitTS0DweUuIG0lueSZh2
MZ+ewaOHUS3k/FGh+d9mll1A00iFxPc2euTWdI9u9vc1rPp90/PLBwyeOUbh
R3Boea237E+cYo4fre5tOvwet+Rrmwl27YAZLZWCJn5zwjt1PjC9DWAIddQT
Vf1UHtj1zY80djmYa7HH00qelBT6ZR6F/lzw2aSeOHDM9R1CCS+iq3OKPSU1
I2iiAXlfVlHcbRjPLL1Mcrq0MfA7s3U1FZwT2pdRdqyh+NFZ8X+eQhJv9/O+
cjoNn+vIoG0GA4cf6GykEy0anH+FqA11jWFwYeMLg9n8D6wj60EBvM1IJUkP
IrwZNA899Oub5nb+DdHZDg9STrTO9n7z0Z1oMMHMH3iFSoIftijJ7VR0Hvyv
O3xUqHsrgASQP+3s0KEGWSCe7tOlc9Snjscmgcox2nxp0fWOfyefVAaQ9rky
SFfn+9Fx0naJ1aeYZwf57Amd8AhdcysGHhnc+cA/MoaIrtvR6uGhylOndCaR
ZXUf+LIXgtjuZcw3JVm6FOSTraO9VLriHvXS28/pzUUnirRHIIi0XMWU1Pik
01UfvwXTV/udp8humlPic3/B0QCEJ4q3SBFNTYDI8JLXQBQI8aOEVO4x5d55
30XtsW1yDGQyQV0Gigj/3ozFZVna9Ktc2skU3BLlvUaf7mYjkctIx/wMI6vO
r9iAcuiSRxpRgOLalSiznP2PdcrIEkwpj9aaW1zsRlm3R6M9eOgGz0QiXNao
cBGlLaJfIV2frj53Arfvp/+vr7bSW+eWujiOE3Lf+I1gxyh6HKuAkG7l/C2h
GFHv95PDcZTi6ZqQROwW4TNrAj4w0EkinRmbqWDlSBNXP89ne7oryJMMobuv
7BNNuxKkpPFEUrecRYz7tFJVo3/4Pp3IHb8My/eyh8B78vANbrbRmxeYuLkB
xFEkmyBoTeXWcpjErMwprYw1U7gLXouLGcQmAtAkXdUoW4GsbQSMbDWpYs4N
erfshBhGYYxcibdwap+OWP2WMbhNgJ8gwZsYnq7B45OvWebUsHGBC/xcYjsC
5p9LGMStOHbbg5j1gTGA8arwqtTXNKRo1kS3wzyxFtrmfSF3f5LHFEw6ukDe
HPV5j1EyFQcWJGcnEeNBJp+DMPWuxeTz+o6i4gpxecoTF4TcwGyrL7GkIScf
WCgMWONNtJVyZ+hLUkULhnC9+caSp50WSKju4T6ibH9ZcU3I3QwpuFfFIo9C
4tyck1Yw9bPsblgP0WiZtChLiMtDWOBP9Y3mioadJ1BayIdEWEOpTR9TUXtw
Tzl9WRYQJUXoZyyK523J9yIovxi6oCSClDCgj5Mn2jrCpvDkVetct6Ry6/wm
JMwTlDxHUAG54gDoSo82uCR9LL/Lo2AINWQ41SKejZKaCMY9B06TdShDgX5i
CrH//44Zmt1rufFuM9A/BCnp1mXE1i//zZ1g8yupVjmvhbn3QhSRx7H352Y1
x2zypPNaGpN/8wagh4rmEoUgfLeveUNyuyx1nnQHXNJdBSXF1g4ERwsi3vgW
vYxGNO+fGg1JY+jo9dAwwgDN4vb3ADkx9htZrq/s9O/Q/4x+WLaXGyO8Xxum
lOi6P/KcvM4CtLTjzhm2tKsKZ5x1Zzbb09DehOk5qckYUxklb8iNJqa81WBt
41iGRHWVmglaAFeeDbzZA4rpidr5JQHsxqBPeIn6NXugpvuaIxrzInPSO7JW
CcmrnCkZdz2c1f2PR2Es4wo60gqnTwgG4P/ESURb8PkbA6JBx94IrPsHjLlJ
X5hDEp6Z3mU/aLcQDRCQQyAuEnysGW5kMtchtbcJwASbKoeeqIPq3kxAdcBc
BpqJ7upgfSFBDrjHel7H+fxcL57VVYa5Ku96JzvRFrWRbUNiWOckUOTkC9Hv
XUY47+zQ5FWy45QJBeAxe2K/HAr2Cb39rZvfDXaSTcznJDVNNHi8HnNnz7wM
WHEVa4s6YuB3+nRfUJETNOXZDhCq3+SmMizUQbhEfLfLkxSBsLZwKHyqX8Pm
t1ukJQCuw5J0ETatzXZGvRtyVkuFAg6cv8uF7USv/qyx+R9R5xMUAkgsqkm0
pIEl/8I0+HhgpjVOOLKbQy0xQM7rBa6GleVE6DjpHB4E3gh6LyK75js69OHS
KKtKoT/RL5wXCiBS/J+88reqfGBkt9DFKHHG0r9Z895W/mH4RGqfj9oUlUow
T5utDPwPL3pHuYqUsvKZxaGZq7+HHC81ejMk9dwZaKMScDxYGax6cY2hEtJr
urdqroIUlDEkjBE41jmHmoTClpt1WxvAJ+2qKdtmzfHnmUunbdBNHFyiWWAv
x22HLRUoDLDkyZkrqz3NB4bhAhqfw588Fmg19cPcEFaLYcAnzZoZveZYjxfe
hLDOG9AJe0YKJLx2iGMCB5TxSExUbvuf4SI3zU/XgwnBu/WgDSzG9v7hY5Wn
hJTMegvZ46+Ui0bJyXxBStwBm3OEn0/EYRT8IA3HVxapDW0IAgiC6EaYaRKN
+1KnyCqEKZj9w4tulSxfYAPWsd8J5zboaVp1WM4/8+rFjgEXFTqUYc6GIoV6
OHSq/WeGXlXW2DtEyGUyy7kxd6qrK/WjRxZNd/1cfbTosmMHU1LwN3KthR4k
ZNGfx1l/9o3zv144QEUTLi/69xvloH6rnmh1Ay5PJZP0g/Uo5YV5O0aoQ7Rw
F1Ap22SJOb9TzaOlofw47WXmEJqztHtx12xoquABxRa+vrNSyoPa4uJBlcH6
1TPVbG7+VqsIcMK4a3R+HeOFABYdcvypUNTL8RRslpXcnq1t1rxg7sn99eEH
rWBTfwOYzmKEpqHuCXnSQhQCnX0rU4oYrX0uz1LDAmLnXsErejzBahNo9BHV
Hb+8QeyqNLrZGOB+4X2pv4p5U36tSJnPRT/HsKmSEMqVpvaTV2uflLuuPPDS
So1F5dQUnS0+YDMq1D5cG5By2MW8NdlYGYVmBoNyVY2hqz86Iz001emOapxy
bmg/0D4UVrDaOA4DcRa57ZoJjHqmLgCsdgXYgaNpCuKFXcBGAyKDKns6qdSd
ODB17TfBHcdIFSkAa3JF9BSiKtMYWCwd9gAK9JtjiJj3KJEKB0d54AItPof8
lxNTkCEbnuc37RFdMJjYZBkNarcYVqz/KwnQ/bP6W87puFylTD1AFaAXNbdX
k69A3dKF8h/nS/TGFXV3iNkHsy29YqP9C/OtFmI3Xlwr70NZXL2MePQfUl/o
LGFHqoQEHhX1nM4VAb2GfexuzlTxU0gUaK6ZtqjTsD8aQO5raWTYbkZK7Caz
5zYdYgLHL5URdQZD1krn2uC4Xsr2+5uprP2sNaCppKw4zu6Hm1Y2V19w8XGQ
kSUl91GHODmKCeE3sQygaOzpNJCi8QpMXDU/9XXimMGR2aD8jnsdR8YShewx
cXmJTMjNvvhOyf3lj3mqMF2/7SRVSrMKQkXOEp9KjaFx7t9/XkS6nic+YuH+
w0aZbgAp7nXOGaRRw0i1dgSTMVHo2WQD/bAqmtYvoBKP/DmwxBVYc2RfnJtO
sbNKUE2mdKBda3NGJMZzX3ItlBrd4BiwUmCYjSc+ZYCJyUPP4y0CQOi1tQmB
HAqLjvVSd4HSjyNpp/JHjBWZ9ttPgQHrl4JnCFciAmYmbe2TJwwa0/JrzKcq
zOKTM7LYCNF0XcYATqTkyi6DVDJf9hmHWgCj4nhggUDhEXt+HqhfVV7+Jr0+
nZpCHLl/60JUnL+aW5DlI///o/P4f8OxljwcWCL464jJQ7ezJxSudtnk3ghl
j1IBVseGjEhf1mv9C6ALgeSlIOe3h+3/vjc3TkTxYRRfE+IbqaYTyEn1/iz5
TZP3Vg05t1GPSOi75zyQWFYYI7a5YSNO+Q55r5l+/laKCl+1UkXkdWTkg3Qk
iOZxCrApn9LEtSKVS7SjtuhzVbCVN5OqygQr/ZrIM8nnsPNJ3XQwvn8ML7wy
shiI5eXUqTm9LaNl6Hu7QKwyoo/L3bgGZPaOCghcGOqbX6UdUc+BQH6Vn+pG
ro/8HAyQgYR5W/BvdQ6Sig0N170Idqn8cUEP8SBwKUK7qMv3oEDm7yyQxpXl
vqvR+taDLN9cKVyBX98/csAcRmU1KJz1RiwuOMRAUnAey6m0uikac2ocYBFK
P718UyofFkR7+aAsLCO/WHiWTu8pwn6x3tg8XQmMRLNaTwkCyAqwyA2twPoy
ZzLYbK2Y9x0T2LXJ44jWXnbUrIrOphrPXu4criUjb5OcWWvJmLv7MJb1ANmf
/VkvZyyts+Q1CAuA4xQtFXr8zDmKrRkT6fv1EBs/d7xnBeSREBjOfR/P6Qt0
1UGmo0Bw3XPP/78aMhC2xx0t8aHROsaDjXmKj788pxOlO3qNJad+HNoQO3eO
PYamMjJXqnR4anFaItcUHmpdxW2C+PDALV94a4S96ABfQavoI6sW0zEVczrE
UnKaGJ3n3I2CHqgDbERP4XhDHR2pjrXztqrOoTXNomPVMFdO4k4+TuJEvtDw
NHFH6tlPFPy3MmfHQW2J3eLhn67cBd6ehqM/OjJSoPGdZNVDVnXYHRGAzorO
WsXS0J4/bKuPv9zrPwc1Xv8vUFaNGwFG4jwQ8TRUVyjPJ4nwNyvVDrBzFP72
uF0oHkttUb9Zejj1D4JfrhJ0aP7fujydawoLRSJLOaXVVhz59AuLG9KCNSrJ
N3t1nej7NvXyccv0caVLE5I64Afly/x2ObsTx7XDITyaV/KR4nWUWca9lOna
YY+k1tZfPf4HkLExOzOO3c6P7U7d25eq8NI2KVOHWs6q4N1IFrgQwrBQh0uz
DC3WfLHnSmt+CFXFkD/nof7FPnEGkajlznBANEodqq4vs4OlLnML7wB7Z+Rr
1TquGX46taVzJ1n3yFAPBem1sqcMJrSqwBmRzecBO8SHMVSsz7MFLBlfv2aP
tBNn5G9sodHTAXO7kpmFIMvaqkojAPs3Rt7QJXnPlMX2+Lcm2mczz/WZUG80
jIRdGmiJfdrIZ86CERd4fcaTCexR6PuCg/BeTy2+yoNPZgpFfoYn3uE6xgt7
yxo1C5yzxWmmsF/ClyvboDRsrj34UR+o3UETGUM+ah/RO6BeKcxjBZZb4YZ5
HIuuN6QZhldILNs2iaG0CGc6wqjdqJcKHhR1pSF+G4SEfVq3XTEkXFjaYbew
Eax6UHURq8R4q0fw4WetGlRHrClkepLJZxuJBOaFtbScORpeKYNoJAMmTiys
v+M+etDI5O/Bzaw+ENuHrsytrJfjDOA9UlxFyB17QbfNJhA9Nw3wCJIqDnTp
bzv3b3iF2F3T1CmOrKEIAPCMSMgI9LyJeBy35peimYuYoMsPym4Wlmj+oq/h
VFxEJ20Q6VAXjIjfr+87MRjeLNA5y7LacUbvBu3WtcUVcW4crGa2uhvkylZQ
WcNOibD2Fta/vXstInEikzTI4pLaM/nfe9ih41TukNH1aQqAbSDrs+H/FsAc
SdppQz9yidWJYk4EHDgodM6Mcynz+OoF/ZzLgN9rFyiWcsu+Pvn/ODuj/hAz
fUHnkQ/L/EfNsLhgBGYhKt2wZ1fPiXGEDB4uBsy/0P/6WFQArQiN2FQgdZjc
cNXKcMbs0sm59+2b2u/Bt6A+m1BjBhnW+GPmddI93EhaVQ/BcYE0+m+j5cpY
8cWCL33SrsmkAyE0odnD+3SsYzvcRM1+iBwqkR/z2gHUo1hoRqRy7QhZ0kOz
VLk5k4Nov/I2HoxzSr/dqKmMbDaMZi7qrHE32/EOnj7nnOIQEuFDdKtDcxSz
WlhNlllqiOX3cZOgE+iIUBxhsccu7YDjV1MnjHZ3u1v+d7z43Agx/1WJpPX4
TakrXBKvkcuAzF2FRQ+KknGYpKdCp9HvqavoI/993zz4vLK8vIAjCNYuQOgt
WcpZd85CyTUG8zeJFJDQQ5ueOLwP7GsQSfdEFSq5CLddqPyZf4wekdjNnauI
LINOVtgp3HNHC8G6ZzVSbEkEeq8ZGA7pKRV6MB5eq+m20SZSpl91KKm0pcxJ
YPU63h0i53n1plpTf8LnFxVpigZ8Cp3l04dQvzkLXXlh/kewsYf6518FS9Yu
mO9D7DVA70WEM3svlnTojugpHPh8yuSH5gp/gG2Zg4fhX/43L2OjOlPxUXMQ
0drQk8h7Fldm5aMLL4Kc/1twpRp8tJzTLJ/8KNBy+xaVfS8l1qHCLl/EcweW
sDSIgPgCeyZpKjSuIg1tggYx4STQCKtQHsCeRzkm1ZV7KcPYIlCxdUWncK/+
Etf91P9x5DfV7LYgf3TFuGiico6e3KzDwi3Aq25sl6/DOryrfvhuaK68VW8X
Gdq7zzKhEnuoEVnan51oUGYCygBdxTLAK29rcXP0K0dzl/uMiFuOrtYN91gK
kl6h+yAx+E+u1vJHiD6LH6NfTPGOnfBCyAOuMregcLWENfwfMv6wBxzmLu3R
qe8AfqsR/Yl0PEmqTZWppPgXgTpUz8go3Tg78G+57GEnkbVO7M0IH1O+sFeF
3J31KTE8frgoOaRPjOwJ9dJxOWtMlPndFvSc+K5qgoMLa/gNVk1rsyym/AQH
8OjZ/+aAREByv7dl8i0LQohWwdUNrEbpVkbMFJHORyj//4eA4H0Xh+2uMnHf
+Na9U0FLe7W2YNFRaYcnfl8LHVck8IWMYCWTratifS7pWBvVNXDvttMk9t1f
m/SSztkjiSyXK6l9fKnvogvub1mDKjKC+z78G9YUcCQT4SZYBKwthhDtWX1i
k+JHz/hPUyL4zcVr7DZtDs28v2kjJG9I8FdPjRyar7ZytfLxEkDtpHrznRbE
1rkVVwqW8IULvF9hJxnRVMqM8jwyNXkARQNmLgqXDTiqXDMNF35SkxSDUx++
qCzl3B+in80hwIUA6D8nXXwgwk/F7Lf9UF3KsRQNTEzleP6HsUmQJGAir5WW
BrfAk2u8HejOo9BfT2qOSKTnpRvUYAvwZX0hguJ2YWFwBjbCYXzY3WAkJ9dQ
PDSg05tO1dusxNj/Pz3iUZ9mgEy4606vKKjmV4U8swy2rgwXhJxRNIIgZXQy
FRdajPQXae0rf4+mUV4AauhLG47m3JIarXjqNmQeuDBJPcx25+DUusgqu+C9
VIyvGRocVg6IYF1ITS7l1iN/cW/j2tcVW0y/hlwF30qBtGy3Avmw17IUE8B6
rLdCSA7kH4fWO74HCiC/MlHIcgcdGY2sYEFUwYGce8KjHSUNIIdByMj2RjVo
uV22fWnmpr1vPzfIXCaQm6QdeG/VZhrMqMTOnOjSZuVkxfr1z8ipyLvQW802
fKb78L589D9dSwB5s93oIXhbt/S+dsy0CbJFr3kRxBbsbYakfIF49BYn0/u8
DlDCmGkbTwdRl5afHjEoJ6JiJ69BDnNCrYGRU9DwtDHYp2ZYyGInAmwZIzfZ
jxVraC85PdL2mzxROXsXoUjz/065P+uK0HCjS8+itl3aqljNLkCZbtDT31C7
WMNEIQb+8hQmY/7dlXgCsaq1EDjZRCeLfUZhC5zCSXG6SEGULvvOFCTgj0/j
EeGKne8XvJlT9s5FQU6pd4AvIeogGrC3r3DK1iVgHVFzlkC/9TeWO0kuKf0c
UQk9LcySpVri/UWjn/SPuJVm2UhvCz31Ypds72A9JXXhOn+bZzVjyHbbBLBS
bonYbtvMPMiuyFhRsJcpMT64RRGrL0XNKZef0F/LJErq66fekiFuRN7Tp77U
zZ7rhOpcWxyzMmnBzU1Od7e4Dh/6+r5fbMHaIbhmwK9P+epziSpwFI8iEqtA
pt7NllXRiBxCqOZgbqte961TfzJ3cnVdumGdpUzsHiET605m9hjRv40TyuHh
l+/++P42hpWOp8HGfs4sAhFwAL6eS9s14BsYkXHNcN0vmt6b/iG5FSCo8gxU
zSoN2fE4ISXbJE0ir5TnxxCz0qvIaud+cyiNK1XPSZLX+26kAiZtbQ3H1cvQ
1mAiBS9uWxx7zyA+aBIOB8tJv38vwU69fkCBUhV377S3WQvWEndt3l2i2Skb
y15zVhV70YARS+xzkxTKUhJtE0qPFMUWMt+kt+zf2xyGxoHv/s+uKuFB1xL8
tNyqZavNbfZaWz0d3fJsEAotJWFxAb51CKGG8QN8tMUeZosZk4C/0Kf+7vsr
WgG1vtDXKUzpxQ/qSpm2IK/04DQSQ0zGBl/eMtcIj5a4ZleZtIADEvk051cx
LdAIk7VNsppXuwY02XJJMrH7TpGe7jZIgD+CKlVZbRK1XzOc5wWS/TA7hDLd
JtY0L2dp4QuGLPDdFQiCSi4RWSF246nIrlrKF49sBG6ixLNIGQMdEX52eQgq
jZumfHmLhfBc8HOwS+u314vuNn06KuJufVpKlNXZGSIlY5yPkF042o7dWy5+
noYERswRb4/oQKducqCPDUxNuWXVQXr3PO3qMR4BlvD4l8nUGQnOmZN9yKuo
fx/DzQ7s0+2P2kuzZ3AoJAHSMp52jwy8eO0+yrAYvSN20L8+rW9ChKnw4chn
c/aaHNdL1Fle+NZWjMRXCG5MmmeLtXNFD5n6ZlRO3ZtafCm+QTqFsZqhuVm6
7Da7Se+L0LZKjG7grNQJ2c1z3n5f32gZ1Fb0CY4nZvYFRd81zeEtSy1F1vK2
NT3u0g0AgzsFKsP4PkEyNirwJZ5GjXMGgeoYWG3iwzCwFQmqFASoNy8CF43X
lob/NKiEQ5fE6Bjr/Lis3ziW3D6ZAYP0GQwA1cl/U5nTo1Xdoaq4AnA2z8xQ
J6NifxYhgp401mAsY7OtVw7Wdn0SZWBjaoeyLScwv95x8K4UKoocaLYkj8l1
aMrOCCMBWbtPzuESwsOpEbq3vA0mzHWj5ZJspwM9jno61E5IrHra77sjHfzq
kvy6xAZ2T7ebh3ItMG/TnfJAO5cJNl/XkncHAT3i7PaBUwGsH90OwqIH58SC
iBrFPY5S8e7fD9f9iR/Uecm/zu1HY7OmoLRWLdMZ5ukUuQi0A6iUcxS34OBN
uDEpe4Hpz7RK/pesMLqOQSvE3m+rj/3md77lG1PXYfxxMZ5dPv4oakul6hc+
hAVMIbCGE42TSCJWGBdoKco3OIffrVsZvNl9jnmBeYckBWnTdxhwgVcUScUb
Cnm0yqjhscJOLEaEFAdO8e5uwEphCHz1r60A4aeuXMsU0GTs08WNH3SdUqrK
7iwm8H3iLaNPRVn0/+25Jby5U90mOobSyGK5Y8L4A1tztg25V34DjRyLlQVu
Fngk9MGgVzdtzjs6nYjfFuhx8B9HLXoaf6IIWdsUQsnLwzA2IHg2vkiRUQSE
+fvEDJ6zr7Yar5GG4KMfeTVO4hhA+RgfIzfzj70BpGrF+TQlqjxfn6Ere5jl
yJXfKjR5BvjF5nuhSYZkBWaXdTqApvVGa//QmWkZ8FsDHRE35ttkb1EOE+nS
QZ8A/ZDo5hEpHmgbU1Wc4rORoDCi6WOcM6oeSIYtRyAsgJE0jQSCie2sb0MW
teoVxaHFCwWw2tcBCQ/zSv5e52kLr50L4IWWvu4afk7kY2D0mmlNj3/HiZBS
pfhxEHbV1ndPuCE3CXQS608qX8cWFs+9+fmeFULFdjrXkFADqr+EQv0eQZ1I
xQy9A290nb+lFl09Pxlqyt3URFgiWEATW55En8ZKlV6OAIPo4YHddccnUjR7
tU/BTNdQqUbT4QL/o+FZYL/3bLLA6jahKuKFBClZtfbXi2qwv3YDGUVQIEiq
B0tyqVVDt9RZAf4i7iMhHmCANbLGljLNnkB8SEXQA9GRY8NXUCl49qodQQbT
6RVJZRt4xh2QZb5AGG1w2e09D/jpXr45RBE6D8BvtAWnJ52XgG0YT2do2qul
DPw84Y1U4H8qwWGFzZys1K8n/KA41KhfjgPcI6uxdizYR3Ehe9H8m9rZ+5n2
sZEmP1mDqeQr2pnIukSQmlokSCEwL2XHcTPFjMLY8SUoPYXcIyk0wBiBUFuK
6KE+iBkK1AjfTgObAoU5rfdZ9SLFHi9qaRyo8lxNhyhV/LCNxtKq8M0d4jkF
PIdzs1JCpu39gIGLT8RWgPzylK1SMrm1NqjbSLCYT2PsLj/F9YVFB9xxBH/J
/FpTs0OWlGoTtG1BIuqCULsxa3lS5+UZh6hH99T63eBugbzsIeayeTkbF+A9
++bH3xLMuLtc6tP0UP3VIWeZrrPQ883Dn2xHL5p09GwTlRyrrO4nPbvER5pv
nszJJLW6F21Y3zJppm+kc5RRgtGXOKYTKXYCcV8tve7vsUuXrc+QArbwJOzj
kr3xEBqAW6gjLoIRRgmaEqYkAct1ToRdKXhByu7iZUftqkH19uJFeSObOT/0
e3aZYRvee76p6bBbFjh71FhvByl/cYKmZpYTZZntJ1WF6ffc1wlu3ongQ7R1
bEhssaDmflKnwOav+17zcMpBHlRN8XOte5636n54JXXM+rLBeGGCyjVXbTnA
DJbFOncQ1mg5lTXHB3ZxMNsgqO3/HxMYcTDSVRyRjDF9tSYsnFW+C4zEWUI1
CyZ+/rEmaylnwC4c2GsfAuyN3jDAefivliwyhrnKbPjAAk4VoOGLu4UJIQlG
UIWLfEx6DcM66XoTe89NlUsPkdrEqpBNPwvd47gLDcaus+KnAjDrlLDLJdPM
rLK2F/4nttgxkRJ3uP1h6zQwaGgplTRYVABLRIAlLuVKi4oUgnajmWHcKphb
q3FLYcXK90azGWLP4eml4N/oUzV6wzbaVHTi1mrUR2qHtffVjVZSGfK4MNtb
UwPixeiWTKPFkghbcoqdKpoJLoq68WqTxT6/vDRJNkw2sTuD0GaB0lUSAR46
WQPh1NSbBt777Gf+Vx/NdmQX+983D8JT1im7dwo3VIgl0G8UfelJCZ04TgQ3
dM9XHPnLtvWPZ/cPYtf1jsKIBspQR3pywY7ZsBHq9zHBoGsPa1e3b+Csjmw/
SdJqL2TpsruFXrxbq62jEA/SBwQSURonah/FVbZ6xX+Q4NewS87fUW59eaxC
jZhjTl2EUuYVgBIrqTHj7DobfMrv+p0DLuFnAkj1iekkXB+AVJQdfxoc953L
puDujJwLt3Ldu+TPgShvSc+0DRMx1IL4VRPO/k1cJI11mX6WYsXwALAtt5aZ
H48yMyc4yaDRKCTiVVKwefAA//K0ODq25NmaMy7VeKke0GS9D/U5IzFr5XUe
Q7m5+xZDoHQVkup2s7Z0P5x4WY5K489UxmNCVxIWUkHiG232ANyUzZrkgjth
9Coj7exwSMc0L9bCDJ7Tjf67nEOIaeiptWsUp/6zl8aZcaPLtuwW9ezl0bCH
9mnBaKkE0x3hwP85KWJ1B+YvoE5B1IysMfgH7uJT5SxMsF5AOFzOsVRc9j7t
8nQ7aycfh4F0TIMRxQMobFUcu5FkTJVAi9+WODi68AUDwsn5natm57JVLrd4
68IBJu+2Z9nKF3Xvkrg2VylMPXKyqH49jSFSpypSkItlIHQOjGgvXqy/8WvK
PgqesuMw5PSbYuxVK9KBEMavXPNO2YwNz6BHi7RwJiDI48yMDRe1PtO5oiIo
VeO6X9yBi/hgNTE8bCSkpQpp8LwFvE178KazDGc/Z/RDIdBWsO776k7Mvnmk
WfJrQ4ToxRDaT0YyWQJiQuT4kSJKDjd7m/uzPLdqQyqAMCTaSkLJ4rKAVkgk
JqbD074Ojm8tVSn8m7uOcQ1t+62tUgs9JloaVMNU0nLf0rSWkqQao9e+gS4G
g9ysgjkF29fwTA8RcSqD9qNTSFbU1i4b0/CUF7dshtZPl0rzHQX3MzTAbqR3
z+tEuuJQZWJ8Ruzwqd6A4k4UBQnivbF6994wkolwTZyVDKvYdHZ8f50xgDXT
N2dfufDskqxG7d059AafD4hYYcL+pTOtgDkwjZCBOBSQdiF4joSRzUePTc1p
lyM7sTDi5RxcL9ztXY7BGszMfRZN4UEGl04QyuTov2MWqDrZxqTGKQGvKJzN
jCb2bzX+Y5YKRxCC5an8E2NbXwxhuxAGivh3X3MfjXarGzEFqXYvFPROfPMz
nTaKkdJX/brluIzD2sFTpfcnaYmLkI/qVeveLuhK1fF2lAijhKvWH1rXgiqG
ygHimZexa8v+3w8adTZhXKwXPqBzJr+xiyfM/O5e5N193YFS9bIxkwn8T9Ow
nu5wAzgr80+AnGpUcivvFjys8cqzVv6OdECIFCzZZAWatvHEyNou+RPJZgBk
nQB6/yHr0/9qyLybMXL96c7RUoigQle2asl1aonbAn0LTfqNL4VqO3l/DW9b
kuXRRTEo8n4RDG5V2X6X4oNcnxjPzjyYWyvYJxTwvtPH3fZXGHGhvxbHvt3X
DNkodeCwFsSAZfuFK34WMyMFcpOiqmZjvd9sdj2TawpGZuHGD8zLOFGEqATv
Kg68o4NKF74BoYR9dkOfvH3ByZgV3q65m2V9JecgcZA1Qb7VTd8hZ5MA9cZw
vWnEHaCp/qtyugD6Wn4pWsVHZX8UdiCDbnKrIz7qePx1O+WxQftlGPukcitA
kmMHfDIBkYHbPoCo8HvVdmCXiYhP7wm4y6Ueha8e4kPsmIaNceh04vT7mkom
diOjuUMixj38EqujqtREd+4XN7kud+PulzewxVzh3NffdsgadUo3oSg8V2za
L+GjsNnahsFylPRCKN2oSa7vXeJ/2YpVxeZ3tD/7nNFz+Gr7l10X99nHkf2g
zE8hNj5agrZRQazwjXyjxwLa41q2E7LL73GgBckUl6j2OAPI3PAiNiO5rdp3
kU0/siqyt+UBC1RwOSGMrUcAsfWSjO6owmE4fkqSdrJPFeC+GN2+RyQg5xBL
UTY88cRddWcDP1zBBUKpD4a+su2KSgW4BIFhAGw98YddOKitlSDvf9r4dmR1
q34b44nMZUNgz50014erAefvTtgxpF/i9B6jGWlgWbgXa8Xh/JOYvubylQ7u
yvV7QhY5JbVJUxY3tXrsVFhsp9iNqj1kf4UO2KpRVP4Df8xWczvJDJ1kmEy8
Yi05fJ/aaOhtMoufI6RwdJn/FnSgbVnG5HorUrVugPcxF/BUZK8hxPw4Rcpu
2+aXsRKu0V4vMBzgQb23XQtcNmIQRE0mRgR3KDy4O4f5w696Kb5fB+T2W899
cJSLGcRPyb0N8aAgXqvcTZl8SogNIgxnxdjrW6cuXZuW/ilW9PbDBAJF15Lw
s1bAjYLCdXNrbIXU/WOnub7j0SCmyfcj6K1djacJYPE7KNDzxn7ATsIoVFg1
XMAsQ0EYSgRf9qbnjwvwVFqBkYfAjxIZB8S7Y2DMcaZ6/pEmZ9/CcSVsvPQc
bc7IMKbwkUHvqxuk8LZ7D57Glut1siHYmDs3pUfKq9qH8vv26/e4ubUwcr+Z
9jaDkbZMfZ2QnSov49KFZoBC4v6c727rxTUAq9x/ZHqC3sHGSUFhMOoWxP6m
nJwbDNDju89Kw7pN7TnK76IeeHwtDujvKm/mSsRSRIhL1mPobdVmwUxz9TRw
u7hWeKzHgW/jIYuoU5yopB6nzf0y/NZ9CSCCbM88pIG69vNigZK8goqNz9Jo
LXKgEaNvOJZqILavjx1zpv32Glx8lW11ti6deGAEiJve6zt4A/pjryiEx7jl
WxpvPCKFSjYvzl3L/tmSYhfak/fuB97PUSORVqAQsx2ExH8Krz/MsXWzcBWf
BKdzAzGhl+YlbrGSkakNPF7BsETEzr3/1rDPRYdvaCWKCyscjVqYR6DTWM14
Tcz7tuUl8aYglKJ8IHvEW4gOZrgMY3EneAPQgY2mOOANDLHTy7EFL8Fu9C8X
YUH9Mps8ZO+Bja42ldwVtqK6yLxSqNYdUrgdTvQIDMCTThVbkIqYjxtxevsx
JYynuG+NR84fwrOdzF4TqjzXpsvwJsszLNLg6PjTXLjBdTRmSIYnoLtqKu5U
VrUYdZXFSb3nnzA4rUiQxw5coHHYhRqh2T8qbOTN//0JkiaBCIEwsmRF7DZj
u9kNnyb6/JIN/TWmmfN3NSV+cNmwb93SJ/sCSZ6SdjYu6Azce1tHKkwtz8CU
muXI5PGd+ByitsQtSnCy3XMVdRjcFuh+4t9CvNp8Sb2TY6ATgmMRlGzymjHB
hbv5i2XvsiS9hOJYVKW4o3HDXqt0O4OFFgIepE/BZYfdQOzKA/6tfmqQZs3U
49NXLqqRbwd+M4Xqxb37aSg5E8revdZ7MUeYK91NBTGYJCQte/wzzxHL7h33
guhxEZTIphR+LMv4Qy6SnHqugkcu4hmScUZRKdWiqjh5WGp1xCtP2/yP/eEI
w7zcVP55XRC9x41s+4aYZxB7yRrfozinneG4QsKiF0lxAkQRAvGts54Q201z
826x9RMGqHaeoNGU7XL9+EI4fj+R311oq5vSbEHBMOVg2k8nQi2e03Y1hiBD
AaHYArBtk70LMp/8sbTeidoWRsinYJZxCNFljqSCFCLjoR2MlAiYScpvfoSp
Y0r9wP96usLeX7FjNYkWLskQTlGL49UiYdUH6+EEVmbJiwovA9B4z0jqabOu
Nedu0VNY48awKqMnDpDtFuigjB1G+Q8fnNh2FmdxaCetZMMjj8awQ5KSPKwI
EIFN+AGuPHBCkl16lfxPXwCWj0poY/zEvrLhWsbk4enj99UN5lBVZ/7pIyFM
/yKb48UCxxVdnV2yszdVSvMnHuOuUnP3Lr0vJ+eSy+grsSzWfOF8LRW9vRXB
Z/Xwm/N0HWDNCAEGrIRVj7Ay1X9C0SKJo1GFlysKbTxGSVYFXBEOk/hdiHgL
pheIB+psTmUTFh2dGoE0K7Gw9Qzmq72+kCHoe7JUNZZ5AeaytvYvbxzREtY+
mfdgjsvrGyRzCHJY8fViCAcu6NeLzp2rqbgsGqxgsU6VjmrL5nq3GnvH5a7M
QKsBGzhQosDqUG3rVVoHGf+2nnJHG+8ddKocQmTLssYmHvlYTJLJbI1ov1Ht
KVRPgiYiMj28xsHnAZEmt/W87H7PNdTLmUSdxNGliqpvy06DF83L/BHDGzT5
3vJa5VVaX91lDgZLBUArMRgnxEubl85gUnv0mS5aZOlxmr4siGEdTuwykfqD
frDYLJNRPHpjZTKPHl1pmMK7gQ5yxZLXjZXTGq8WKs9x7QX8YH3XI8TLGhRB
VgAyNHjweDbytTQluIS+ibXLz8VBdHSKdLrg4gX+KErZFlmAlVeCpQUUq8Hm
2N+y4jL0YhU0uEO6ua5ZQHmSoDm99+IYOzPqH+yBtSxE0Dirmf04PemkyU5L
jkdYmrHduMficj8HXV1LGxja721BgV3mOPz6yIc7uTyp8QWgrGOzYeHRdsoe
X66A+sjDEkO4hxjUV0CDcjJliZl3hjXbHYvJJBg6yc1+ZkgG/tKpnNGjCgAy
q4HYF1HcFgdRPaiNETWj9Su0Tkks0gP6SqUNLj0b1k1GW/IrmeTMSu0AtdaD
efIZuHj9nK29eWoukXll+VYeJHUlQpNc2LWpWUdY+ehSDK/6xlcaR6Lnkfed
xjEhHKWtk4bsWqNQa24Z9rccDdWjVwHw4vOqcCwjwojMN4TMi5/IQAWR1jZo
aSMQbigpOlNnafv9uovKZVg6ErpjfwNu4qk1nj1GO6fxs2C/9p0QtRVKpqnz
Y4moyymmscfGG2RRHTFXh4T3eHYMeUsYaIMg1Bxl8UZ+lvtEaZhJWZeHHSPu
MW5wdBIGw4KHm5msk2WtyTFBVrR1wCCCn8N9ZMoVKyYAclA/pHXknAe8E8fT
DNbaQyyGqIZeI7TEGKFVJYQtPCurZXN3mXM4az1vQ9QVLjb7VJaOmJ0F15qL
TrDlOyXu5hqncASI7czzG9sDBcWA2f3OWokNoFvUmyaTmvarK9N1tJlvUmtR
BEgVjzHVFBl0jycbXZJjtOqVtgEoHe+Dt+Lma22CDZRdxueRcCLZOwlJTubr
MKeMsjba81HRJo0kRmWlAGwnVAoNhqOrlZuF5p/7ubJBAy9iF2sP4iLIzaA3
tVg8ofMECkcXdcmn3p7EEDAk59iMGBWHUbwXJAiBF6C20bBSmzfKZwzZRJKn
n5Lc6OqMMCqz1dSw+zCVTxB58zLdRQ/gzclGAaIa954wk8uoFocrCSjTtWJb
s3inR7dyJJRXmWsy4SKfUtCrT3memk2ZNywHU0iTVLxwkPTIKz9d3mvt5CXP
V4TWEnpuetZyDQVwEejByt7Agdm/wMW0h+D5+B7Myj9Jfxl/ZMGCFwR/1pC+
68o+IjkgL53tc3CsBL/dtdgnHw508zYIIodGVJyky86b0d98QHjnyU0zQkXz
SdOHzdJJ9tOIvgORB27Tx3MNidM8FJ7Q+y13Fv4r+lLupOxTfUifLPiMAl9o
iE0RD6cMXDV9d6QsXc02Ydem8JLw1429/Q2xynpEacKQWrGIJYaDh1RQtVq4
ZIKwDFa8ZRwha4FScaT+yNTkC0YX73I11i3+BhnfOvGpPHa0jFy8qCoNXwst
TMx57AZt9KC7wcZwFHrYVv4d/Yp2eA9MpLfM+LQNRNEPjokJmG/YUOgvz6/5
Y+mtDEtpPE7Cz5AmmpJwVUoWXwH32XVosLOw0/kNO1XPb6J+JdtnpmlNPBWR
B1s3NtORxXninGpG5CuYI0VVmmwE+kfeX3SDKE/HusXe1DXrCVLgokOwze2z
JmdOPblXb6LOuISoDAGFpgyL6fVO9eawZMsNdGc8H/0ahfd5MhNFstB1w+1D
WZLZ98xmX/zU40UyT8amAV9PURDVRTtekC6n/cCrVbAYG+dc7tGQZYIYFwZO
7m0VSfrlAPeJhg7Z3Z4NBUWcyd0AfhKpVxOMIOt4+2jXr8XlZP3CCLUFe9c5
IMLywv3o7wxltgpPSdBQImIK+RQeABeXiI6+/BycTY5g1CVXHl9Y/+imLITv
v78LYlEskQVA2O2EOmxnLt2d9oRS6PvvCggNSYySJ7L3J0wQWt7P0Zss4dSm
VCJI2ws/UMcU1giMPYGoze7EA3Mjo+6lmqR+wc0jdyqAWA7l+nJbqezi5694
gPe0WlpOFCxis9YL908ISrb9IbpuawhA7HygVsQ/IrR2F9p32g+R+nKk3I8h
jUMCNXAp68ATEXbi7RvkRd7pSCaGyt+xF3os1PUo0tXHieRR4WZpuY6Rhiw4
j69RHYkjpSSHv8aUYJbAsFvIFQ087qVFePbx7agsYDISbWWjf5UPDTdrPUrk
hC7vL/0fUMaKANWnBzZPknZMn79r9vIKiu4N1tk3dX6iX4J8FO81/yYP27ps
hZxlzEmKO5tqxkEPU5cWEkryZ42VCv6nWWAEoSHGOUHIpGzP2tHxdBTY8rvO
i3V0aX4UzDDJxcIwLk8c0NkP39b5YmL0jW01RjvlF/KeSbEOwZcg/oCFm5Kz
XM5FQODqwG9WxHHv9mOOo1KaoujwvB7trEtIBrh87gAPQNTXlMkGfYbSFzdU
XvRKMqDTafrI9RPfVs9pzqWd51+hzi1YdyZdfWyKYqS5vxXIsdU5kHOJiOsw
5oBtI0NoqEtS7wT+RtmXIxzOMWPzbpHC1kkHnQDgWeErRu2hRTIB6+PLYNIq
N9BxehmUL8PasaNtHJ/EkBJKs9ayr8DCvqvmx+Z+/d8NHpD7Hic9IvQPmMZi
aK6S0SPefCe6PNp9Yz20sltSDK0dN86ETRK7XOq3SXAJCmdUJ363c/nNmiLL
mx4RE4XNT+jEIoTxM3OYQ30nADtxPjDv2qZgaCxQeDSQl9bkJTIc5VVORSWn
0u77ROvsDipRXXmSpEWOYIsgaNrE1yy7x9JyGaUIZ1vCI6+sl4Cs5zss2FPY
feO95jEPEzBYKFGEiUU7ytgHyGiFnUb8vGk2lrl35qpCdWn73MahBwQAeVMz
bYPnE1xPw298ekRBL69TJ6FC+ZMruIkGdlV6hol5iMa6cVqIyOFIcqG7mtgz
FUxMPbsn6AFnOOY+Hw1jiGRRFflaQDwzC3aEb8J/ifCSmryuaQ8y4GB3sJzt
g3TWowzoZmfJHtAmNAnDf+TGiwFn0aec+r2EELfSgY4H3mmCYHotdpLCp9PZ
AcuwxSwh8QQhh2zEeakwDAuoGLNujkTFZtlW/a/dxpvhrwibVSsenhSWfMec
o86or2EAkM+/cZ/VVgEJYHCsbpHETnzbOuu2aWoGT/Ue68ZZ89kqwFhd9HeR
TDoWj7vfn3SM12PvTJreUQp0jZ1oZ0oGeN2hHUN+pUIKBARut7cspC/AB33D
TDbms7D0IDAaBm8byyMhu9hZ4NsWTMYRxH7ZBw90N6rAar4jC2uAjRGedhQt
pa+RjWz64heG5UhA+Q35IGOnSwteoHXWEIcAMUnFgWdj0nba8aHKivogy/d8
WYLUs1dSsvNGZztXEhApDcX8JKRaYZZPjM19uuPSUCqF+PX3QiwJGfueVpCp
dpLDMjCGJbIXKKn0YWt4ZFw+ZCx29pLiXcfNjcO++XU4no2s5/wdcRtk06oK
Z8QHu2VvFdtUvIUK1SDcvFNQQMCS/Xha8Y5xVEYCRBDXxmGii7eDJ40PF3/n
vPxcRBioeESSn5pi+woQ9Kn3zSILSvjxcjudzbL+WWL32aU1QMWUpHHj0Wzi
t7RORiRabXHDPAjkmeNBS93r/AHaJWT05Jqt2adgR/Y9UXUAv5DyvXV4IJJm
0hCNPeF3MbmkqcvU2kgPrhdwDMbWprut00fIcWABuh06pik0Mwg8HIrFSbH1
ixc+aW+SvnpcEHEkkIulf6GMtGmmrcOWZ0tUYf6mi83SsKAonpO4E4sz16lv
74uoJUBbCfX4awWLC7RyjAAE/3fsnLwJSnJZHpwnnHhqRz7eRThdX/4D4wHi
5K/PCUVrj3JUu090tHxF8yVxLWYOgeaWGcPBS1hZJufDaU2dsBTjWta2TYPC
BTry99liaVjXVIr1PaNdx4daTpFgymIvYKmPivFhl8WHUK7pyDakhRVEtQIS
uBvMAsYZqXdun8HR2ghN4g+z3UFWm6JTvcfa1iNA6wEJUZmuAOIu1TKQ3v1J
1DvRayZGTy4nLJ45G/aC6D/NrzzhGVGUYXpnc93NN2GQAgCU3dc6YdtzjALc
3aXqZna113gfU8bjMfxhFVSUOgmTXNrJ6oX6kNFU5UkM8C1hPNI7d51nzHzl
U7odLUQSMSJa7fgc3L1P+5j9GepbrVckz1s2x0cm2MxDb/UB6z8HmOvLn/Sc
WzCcjj9C5ssj5XD8e6S0+k7m6bmGlwFHzTBRjcukjrLYf+RS2vmWb6eFBlgl
LRusvFh0nxWw1mCrSP8VQ/ZgKrRyTdq+riwf/TgIhN54WPgCv6oyHDd0KAzA
tnVFmXuS9ZFfax1n/0pjBG0n5Sf5vJH3I60VYicvlfl415gOGhN4r2lwAFnw
khym8HPphRF5SHw6XUiWufUKXmao6wDxwgymX+Y7DX5X/SYW46qzNxlAsnuN
52WhJiHeLkWxQ/EAXwyJTEATj3bNntEPqgeXk+A4H+RLIEpMrb4i0O877PGE
aKigonRijQ0jB3J4T5+kZtzfyy5Wd4EG0JV4ZrSbFeKQA3kRGLdjWvng0RUr
tJLkQ0dKcOC6kg6poR7C8ZiRupauSjaqqI9XsEaVz8y3tN3B6RqF/NNvbs8V
O3P8sREGnkN8BhNzrHkR11lll0/LhOfoUwDYCUn4ayD3g/pElVZhaGTdoSh2
VtGLf4w3c5iKGPhhLdFYwTvftTtskW3fzk5z0E7UiM0Lp8NMNsrXJP8w1h2q
xIK+XF7ajGxPampgNIys24o7Uud7qsaJnHJrB7rzxt/khCzEly8vY9Y+Vb1r
pMJ/7ECd+P/w1sCaEoG7oMflpZ2OFBzc039KBv+T7b/N9wR8pg5aROLxDBC+
LnHE/X9nuD3uB+Qf6pyJxZzvLGKKDql05SsKKlTRLlOkQZo2vs1nSWdPNXsA
bvys5s/IVZ4cUMgKB/VyariU/0Eoj3WanCctv43Gh6/ZQV1wZUzFKMCDgpC9
Lfkrl6YvPHM7MDPvaaci49kSZqrNYr+9mqAzEOp2bLZOy3oxRsiENZKjGnwz
ACVtUe9xhUxmzynhZR8FCkZ5kleAFYhScI/8KmYZG6Ab7pkYmug7by4KzqnY
vKaWdkqC7HOkYy5WlJS/6a9oAu1Q15A1mSnygPHBWoT75OgSNDB5JoY5vNTf
y8aUUhGwM8tuw+ohuOXd3HKVkPsexe2uQSTxyARJOUMMDuMNTcwRTqY7UCzA
xwcD5SFGuKBBTX5FIF9EUoKWEpDXNd7Pyic63kF2aQJXVkLCDlXuRoYcuUzL
a+5HIPuNAborkAEsRe1fas1/n7uA3gA+ltiIV6R4pcOWmDDHKI/KySKtJp8+
a9SNYYZoko1JtWZ/LX2p56foQUtquP3sdNJZ2YJanzISTkSYpZsExMk4W3lX
9RqsQgj6dFhbzAX95e2RYSjHghV5P4gm6nh2Rqf3MMZLfCRkCV52gsoBS2S3
ej4FvqLa65ClE5aytUZ5dWytl7dwwAFMctPuXZGgZUxIz323CiclSJ01W02G
i+z+yD5Z//lOUvrwS/EcTa/5l7CE24KIuHTNYcB58p4tIn+qLqPIWLjRFO2u
TYlADwXk1/nSnSXD5BOjZtciVqvmeWRTcS4fP55rBpiITvqrIR4lPq2N85Ld
SnnirvcUpL9J+WycjrO3/BTjMZ+bJle9Zi0Lhbc03jM4UXD2uVae4lgXTXIM
J1i/4j1aYDRC0vnkTm70ODMfusl8R0k0O5sLYPKvUbmI9VMknkjWbv5Dxe8S
CJlpF3LdVxAikLbbQRoBMRiF4eK9QpGf6iXi7UJ7msGyAZ/gGNiOWyB3VlpU
q9xzPn5QWtiOmb7Pkw+GcapobvXdq7FLdvQGj6GEg651ERtiDuFL0CfZHzbu
ObJ2EvsOiu3G9rApPTrGpqfRvl4+vuotSkygRejYggoL6drJUZ7V2hI8pFCr
EUVZ3GorMzQ0+WMuTAqE2WRRhAgdawI5w+La9wrOpmE3cj5yD/RTLOutKRv2
teeBMgG7xf8FJPRM+/mOJuj/zaoOX3vAYpxMrs1Og6qpqErhvURGVwN4pJHB
lp1jC4gNloFc9Ukyyb3UPXWjiE0Mg9z/rQgUAd29wfeNKNqD86NcxQNyGLCD
vzCdyi27OsOw2awUXOnD7lI8/qLeiLFx9K+xyt55B/pAG1rxdeRuW7mKVmvh
w4Eq/xScRgRTxhisH0n2k3G4eCUsUXJiSkEMaGVbdneX2yan4LzVXY9X6rCo
mgXzl6+DuEZHonEv7GcZ9vF+aJwi3xPCK61VDfoE+Z06cTOH4V/Ec3rh7X/V
hmlzi7BM8kP+3NidFDA+DU6VfLqZipca2qHOKm0NdGTM7RnZctOWFyyc49TC
OF1TkTup6lLW1MkoiZxQK/Z9TMyiT83oqVf1DSYyK0FcGB7fA5MGjIqGNeke
kMfHjN0a+Ir+lnToXwMVttrABpNzeQM+qly4aDBS8VirURCrOsMu0tHMrS0/
ZAdL2wZZ706ouzYUFMeR249dfUcVImGG/aKqL3aNowOak2PyIPk0/7aBqPOS
3xl3K3UC/QU5skTtcq1p6v5J5hCPEtagJmaEvad0USOUJqtNQD9ke28DGtw3
0BjAFx+J+sHl9qx5DKPFg2AZTFn5hL4pEofcJ6xM83+58PiJvjLgeLml7qFI
voOvfkAU8398y4s/6zETrwMtO2QlKLlsXOTVD4Rl17qotduI4pRERwQV7M0s
MoLGr5SIcMBP98gNqB2UtIDOxIdugDV+luBizJmT1OvrwTudM5WXs5eJIws0
Ot/CeKTE1H8KQUJPAAw7TFRfOaw92C4tg6sdGLYa2DQfU97WXzWUzMMu33k7
UsxT09YLrymfu0zcnrXa6J4TMMZlBcHs50VGtgbf80nf1nWiRQRZtysNVYfG
2A2p8xGAo2xZadj5S6hNLfIqYGFwYKcrk1ZHkmFgz4jjMSXAw5aKaMoxZhg8
ilECtWdQDXP7leFET0daL+pfTy90BOTd7VwESNdrq93E2KIPF6dKmUAm+d25
d/AAat5IxaAZOGagZPtDlveHdSX59TA+FB+hiEbzA8Wi+CLbVVt+eRQHc8VX
zBUEQDaToqkLOavP7dg/GugyplV9T3sOPGaebaQyWf8T0fe7Lpx8XsUj0qs1
ATmNoaADeUX9rKLQtJt8+KiEfvLFgu0bTCz2rBwKJq8HHWg8sGUaetCeFHQe
7SrbpJ0dtQBVbcDptHDaiGspqLRbTEgZRNdRAbg8Ptgu63ohQ07g+iyVoE0O
WW9AMr9PJwryCoRUbimWgnzTafTK02MCvnV4z1QrOTw5qjjcEriSNSIouNzE
FfTM3WfKpny7j93dkna1kBw1DAshYjUNYQgIWvSCyjg3gJ6oSZhQ6HyVBuR5
hVBKED4G8eRm7de7yapflzLRW4dAq3mRYyDK0JKReA5tPJOrOstLF2xbX9we
3NgYVjGAI+UrUCSFv1wh6rqL1ZWDzXNMkj6r3lutkghp5IdOA+bGIn+YFKQi
OQbPbnNzdR8rqaLXn/8HnMBGKMIckRO+2FgqNC9CHTjT5kT2SJRRJ9rmGfgN
swnGFvLzqgi+Xz/E2q1NEOSI1eO/LvKgg6ISM1094XaeOWVu9A0JkXRKqqY2
PyZstGfGw2HphIA5Xc5YDOz4SQNzpwwOfSwNSBhi5vgaPKuodZUuBlUi1aMi
rfI8m8HdMZM6oPvDqf8AAnDnRFI+ZfkuY37OKxXOQyLunCf3NO1Z3knGhesa
uNDsropw1M502Yw5YyyiDbAoNL5yhfH29QwnJZRiO+1YWHPLy/oLQscY4ViU
yHN1APMLzPpheG9Qngz5IojGYYDtNMcsd9qA0aFsGGvIsmJOqYERqAGG9M56
50Bj03US2Ee4mWVY1Kh57/z1B0p5SoTsEShOmN6noghFmfg0fSdOzkJetva+
MTiViAhpVSiWSdaHTDW6W5ccr3ZchmcNUTwz/dbYju5ZwffQCScuwISraf5G
V0ZG25zO73MhDR1hdFvz4Pt7EMxXRN9O4I1HjQAIvyqUHR1K66WZzjPPH8AJ
Hf8z+4IYhp4hO5K6VrImHVwPQS0nz6H1Jl6sBQwd6YTYsl2uSBgm5athO6Xo
KFSciTQ89k25Bea25+J9TWq+WtEiihP4zstMpJusgJGtWtbevwyVY5snQmZ6
7rYMGeV7Y9u5rZSybBdT5LDgyv03mts3gATrEqTopGTBSYelLzytnuW3WmI2
6f41NWhqb3CdfZeQajxdUPDwAIkyRaMbBRcvHPfSElvmYoUUKzB6dr+L+TMO
4wo1cCwnWU5U8e386FigCqsnVs9darT3a83CatLI64OqxZv0Ld0TTobO1Ygv
vuZu7CUH7fveKsqX+MyXvmWSnmHD4pwmx8NUe6RLTVIzd9kUdZcdkgtw210R
jnd18EfjpHylRK1vi51nplX2HvBrs7HLXH7Mz8SxkyxAMKOpBrK5mmgZiFht
eYycoG1+1SRB5GEuC2X7qeJuLLRpkAiR0JvYr9DtYaxXl7qfmmpnxT95HRY7
4QznLMUaL4+qf1+Iz6s2++NTM/7s8FS9NAyURqPEkoLcNB+Wz4GA+XVY62so
056z4lg7E4pa9f6Wh7t7ugeTOLjrJzGgtGPIVV4zxjz8rH+BLAC5JR5dK0Ov
pnJvaxWmgmLINGM9WOo41K5NA4Z+yt5h81XkzqVXVYuSCpkHvDnMdLmPPWTq
5xomuBLaKy3EPQmnNmqvefVlUAnKTA3lrAHxhZ4NvypQyqdvAtbNXYh+KPFj
gFYBkvYFamAOfB10yH8svsHf1/aIFj0ZJyeqhjWO5DScfe9yk9kDUs8e0s69
V6+1SC8+e1zV5zm5o7JHb5CiaI1kptqgjiLguaGQ4yD5KQ08KrL1/aDNs5Du
c6+fQjJvPWTOQgqVWG1GogPXajh3VOdkkQseRKTUj6Hu7WCefNEg0GEDnZtU
/73o5QDa8vhXaceh0cgnVPxgCE64sAO2TdZtYi6lZVBm5LOBHYUzdNtv6bXN
UwUTamKuib+4qOapbZPAICQyj1vW5vo7dHcFEymrLuIs6u+MKMDx6fMO2Rar
eNtKkJTMUys4BGQJ//TPL8Ml56hNq176hL6DT/cVFtrCiKl31s1WcSlzLd/1
o7iJLfaC9cYQzmAAw0p8T1OEjqtu7TrYAoPeNyPjgfF5QmCrJzX4Uc0Umlfm
oZvM7//toGY4XPS4vg6OUmyWFjo07xPusKs+DyVzJo/f/E8i/+J+UEDZTfts
T6+Ksk4+TO9FWKcK91d/4cTe3+FhVlmXAmtjKMpEGWn0XC+6BxCTJKTdLKeK
omsru7evkJWGDuq1Iof+HGkHQ1zKOkTrF99CwoDhno+7nc/ivGwhzobe1Ts/
c/8UOwCxITGtyfYqdOTDQBQWIoAYK1V7B4MD0hdForBEsRZYibd/2eF5KufY
PNVoKjsx+b5o0Q+XmIhGGp5dtAPUIkEiN2/4zY/9ezPDVwDh4FcUYrUIWbD4
MZkKBZUwWwI4Xi7mjKvHMj7OGn29XAGqgHnNDSU/B+mmlA8C0zy6IKEy3r8a
vQuRpSseWoJ7nNyNQ2SPSZ6V/vFEsevW+EYvidkTxyBRm5jzvC6Vzz1gnHzW
NIt3pA8L6OX+/8yOx8MX7uh1xXk5bfn2L9PUvgtIMMHbrku3XTbXn9ypEUhG
X8uFBym2fiNoavpOOXBVPOV8p5hcDwrVzReK0NoRY9SGOQ0oYhGgxjPfdRzb
YIWaM8FJ2o9RSKsEuo9aEm6E/lwUioGQqImDsD2avFqapjyw/Lf1A1A8sM1J
pT8ziAiak9FZzNPSNftxNhNamxkNu5U0RW/5XAP31VpEFTprcPTyVoBVQZaw
jLgBGb1yg0U1hLrniXOI3YgOxMxef9DLmyVfWeWHgxu/HHpoVZjaZZVKmr+e
OCFyFhaslqb/NFimUZ48Q6aFtJsCaP+ZS1pGIYv8Mug1S1PPp5eEP3/zmAIW
2jJgMsFdeXZikFx5jfg5Is4XBmmVlZGBGqsPnHf1alX6AL/t2f2qgg5H70iv
eW7KIWEnjY/D2P1GSC8NfilFMq5V9Eul8E9SvvxowSzWxRKqu8Sd/r4arwZK
LHvhdveOwJcG5p+HQmHNnT7peBdHhYxbG7z4cPmJ7wKfQ7amdteQ9yi7ngJj
+5qt9ZamtLd3Uya37+5O98Tus5C+AT3oYOiSxTehy6mX5Kx9hd5l5TVXXiwQ
7bDin3RwMdTszi+ldfh8b/mqNTSeN/xtiZcQXrtNhs9kj4AA0iuzswouZ3wi
qD8p8lRe3aZaybQdmdRhM/MrFRHF8GixP2mXvhMZGn3pj0k7CdcEI+KbAhEE
+WY/NHXXfZ+eezC92jwnQ6c3sAoHLbPzGTHl2uHFHpc3f7DpAlYNlBLODa0t
zdCl7edvfIdrhxIMliSYwXrg1DoCgSRu6bbezsakR+UpaRiaK75ZhgXGoEa4
IJZMJtOb/m/AVC24XzuxnuE3CpAFKdTpPcXiVM2Ut8Dd2Htq92P83S77mDFl
Uw/8M+OUqsWc7xKZPxWu6iK2LdS0V1009QPb1uiJ7buuBgj3OkoEiKFgOLPv
MKpFeUwCBr4kAmZ5d/yr5A7sJEz4+ECNDlwMEcxogCHqnk+q/VnlGuh6tfv8
gM5eHDcOJFrxuD0WcotdaIIGkJ/Ju0l14wJOwcAH+rg+abnXS+WflsjngdBL
AVmGkq6xWWTYBMj7yg9XF6w3hfA6gVZU2mwk4SEi9ng6LFZ6MI3ua4cCsTs8
OHlFMvSUaTs11rxzU80zB5VtmxE0WKvijNcUukx/w5D52cgDdZKbe7skzDIB
sVQ/VAGYrX7ob+627jEQjGTe57AShZyysGdWlVDyRA9js3F0g3+/49n0sc2G
DKLCde5aGNKIq7JAYLNXDWaihtKKorlK+yEwPtUyLEJvWEGatjo8qn7wgfk0
2EteuaG2SxTZQ3YE/qvxHx1L4kZIwT39+XE/Dkxtzd1oqK5IgUwd+nJI+FD4
vSxaFy9sYPIIuVaZKWblbg1G4RwfFTMxYm+lPr4UknDyxtIversQdTeOJjJS
1gsKsgUIEjE8Lj0rIkHTD6DX4bw+t8Vbfi7+RMXxTSFG0SLEqESp8qOdwknE
BiOD5lDCLiAXBvcYA9kbmC1YB+SurTri3i0XqbXNtQArau8HrZabCgXPY99S
3mE/j1ak1TQu7dIJtLIx4l0093xY+Lzx4SE1oNMtG7JB5JYvTRwCFKOBXZ/2
UHvbXsRp57fRGNRX2+9tombLfAUAWiWWXOKVKFmdDf7vQbBIDuKlOozh7uGS
jA1LMr9Bx6qMpSAHpyiyzCTLbXXnzaJkK154yFYsnTWVPqGMq+56EJOS9xGR
+TJoNMbZD6l4gwOGeiXvmWZ0medTx+civLhCw3CUXP4QZLcZUkFb5RH9c+Fm
R7Pfl3J03lgYhng1C/1Oyp9DRuOgTUcO5RqC9mrfxDI3v8Y5bAN44JwxwBkN
kxd+/nsBh2RpyOztfiyzSY/+5f6VY7T0pcfDoXYOlQNTYqzRpNwaYrLsTh+T
QhS0ckxyn4oPD79khfwVa7JlBHPRTv4suxS4Prh7pxin5kMEh5mVqNx8jdh+
31ZtQMQUYfuFVjDLDB527J7j5xSV+4+MPR0IEWB6/IHKxMx7gIFMe0UiLxkx
UFbAWMzmNWV6+TyjJZ2gHXgnuxmBh+vk1hst/nWAB35j9neWLAynukBVYhH1
h1sc1IkrYdR8vne1M55hqJVAHtPooHN2PdhpLgJKXOZ8bXe+dUO5tNQR5f+q
MK656ft8s+3TLFLE1fbbw0kjjSFB5ypTO9zKPRMcXuL8oOBOh9QWCVj0c4Oq
l6xOpXY+Zkwa7/5pSFqwf67VB6/6q00DDqv5ebOXy9MxdWCU4lz21Flp0P7r
FSBlNoB7RiUqL28NW/UlCXlfwxH1WoHJxusywnuoMM+Ua8B0jhwfkAeKt2Ar
kMvnTWceyR24HMva6Neq6VpwkNGo+pilpSEBTIDPB+gB8QW0lTFySBHQqXMw
U3MjJkt4bClDnvNE0MMtY4ajlMDzKieLYGr8D1zWR0mIopONqkq1n1QWsVSk
o6Kdn5owW456B3C4fnS5idrZQdkWhuyendVZ+XDztZEX4LbLHvDbvdJ299I5
o3/kCmncM8bTvMQVvZNjeCEwONOv7hx9rMjE2mSodx83rr1zJFHiQnjgVAgu
L0MS+TupyU/UEf0I9Tbk06OIpyyVp7i0uQumXWGehFdsEY3onOf1tt/2ie6D
056E/vKD4uXYqtT6oP4kom1OfpgavWZBtXNF3ZgzCVFXZov3vsCx1zZxBz9u
7uuDpXrOBrBCXx365KETc59staxmPbFTkXPXTesqt8BDtQrzZ70HV6Vy5+vc
zD/uRqE+c2hCaNifg48mOdpQ/PJTgpZD+7baA0ipIqlpUTyfdqwBeKQrVNgF
zyFFFnb79HclE3kaaoRkEuCnVQCo6BwqjCi8jYgkF35Ye1tIKfU8U/UB8h42
cVbVHc0D3qlgh1Nm5uPTdgnGqSws3cQ7wI20PTeEfzD2eQ4sJp1o1whbfBrh
PWhuO2OdzmjYYS8UsbhwmRmLH8GPASky9oZxEQbQUNN07pTh2EXWZmIN+pWl
8ZaBSCbwu4DycQYMC+yuKC37KYbBikAr5OhmcUyKmRDTbj7adJIJApQdov/d
0CvqCl70NDBU8ADIBQ7uhpcJCymlryTcv+1uWz9LakQg3oz6wBFjkoaMzpqZ
H3kfFfpzycN2PPq57VSA6Fnw/mRHA0L8LENP4S6E14wHMEY0NaSpAjUBLgP1
86tWkY3n3VAOyqnoRFPo7QMyk1LlGncZFlv8CI9p+E+DHsneLnagZOJVTRE0
+MkCCVbGALbcslp0E01IyQQbJ3dHBMFH53KxMXN6uhJZZxLI6p91bqyT4ZGL
MDX+H8GATV5PtxKi2skJ+M6ZGUKTXFt7wdW2ywEAmhgX8E5zPksawslSGHyG
ZuZr50Hf9GOOUZNArtV3br/ul8C/1tFHoN8rMe1BffLZEAP4FsZbfAnaDrsP
J4agxAxm8/+Oyxe5XFZUpXZEMalqbVcowj0jsg2QnS61xKtWcPI4inOEjlap
jnXwL97hCmzci8WBUFgJHfNjPA/qWXkzCdo4KNLMkTB36eBoe02u0AjTCnzM
F/oKsQtp1NSTC+xHhac2Jfgdc6EV3f4xd+Le+Tc7DFwToa2ZxlAzIxL///Cn
+Mta3wUkFJW8FEvEkDlraPtCqHu6o3DA+S0njpsCVjcKAcJ7TjGbdXKmtj4N
0e7iGiFF0NVyj57/KtXRHJp0pEHtCwiNF+u+rc7j/q5cui/aOymUlPPrYXuv
bk7Y73Psna2NUpSaTvFW3VxUtkSVj+UCGDoJ5w6V0K8udBYErFWEvkp6PvZ/
UES3UW9BubFFhZuOzIiT/uA9n8w/oTubkahJmWskJuQFYnQljWLCdlqzp2hv
pan+Wi43Qd7gBdg1B1yLo+6uqHP7T0oIEUxGLUdub/Ge3jKYnhQoMFw4uhMj
cTybmaxCgw9xrbNF4kuk3+TiuHs1gTDxfxHugZTF8dCkVhALMmaE+24zkxKi
nLoEf08fIkda8yHyN+tl0fiWt2LLEH/6/6FdKNImSPQNFKHFPrFXou4m1cD3
iiuh4diF8Kgq4sH6fLsn5CbUoMhwUHMSI7h9MOcVpw7NQtAtO7BKiMk1kmuj
gcqrj/WUD/7jSa8TzWkeZWrSHz8pG/UcUC2NkV2FvYbOdIHp+CMIQ4UrcJN+
JvjwQGljbZaluAXWvI8AelBhHtriy2EvGFbs6QK1+71nJ5s4FNYvKcuvHt9L
2TdPydsdTBHLb9+2q1lC4caXt3Uq/ieIYBDvYdA52T1hk6gFYOJ3wUndA2+y
nW6pZqNCnWJrl2jtZ3WO38aoF4dmvyB9O1YLmQZSDjSvgY/VCMg4xyR3Ujut
8KNqNcUIS9rGMR0xqbfKTZFJyovJy8vhS8D8iQpcbb3GFBl94hI3Pe+EPKgI
w7g4BAt0k1TIZJcAngm4/MR1t5RuDsEy1tohznq01HO0OIDcM9ey0c1bo7wf
AW7wzfqs5SHkq9MbUsXHFKtGaVQg6/PyizQiSzaUEH7lH48mC4xnNr9KcAsG
quE04XHMBqQI1WfvtCZFyTyLMFhVmoje+BVw8r7bdNfldrrjZCOfSXQT0Vuz
VTTNjtCor0F2TB+cVer+QiKL/+GnIL3qiuVFTVE03hsiXBo31IRQwGgbl5Q/
tW50M7iO2bSr8enACfg5UpKrEfcNAFs10sxU0ePDDmxTdyOvzIxa5Z4tpyM9
kr5Y29RUrdYSfaSC4WDDrAzNTX+zDyCSa+cSqVLsnACMYglzGLFnGMJi2EE9
GVnm9SkL1rQBQgyloLQLDROToTh3u+Clml7bUbHsMxxnFT/YWNsiS1u1OhPM
uxu/NgtaMfrhi/7iUZL6eIC/v2CpU51K6xmVYAm5/97KlIC1E3E8x2gjzBjq
JW5eXJEN9boEZ3EmFQpmwhslepCjeScwD+Wh/sHXkgcqvg9FEespZ8dFWX1Q
HwsMjOOARF5STg/SDy7MwNAQCv0fWp3SYyJE1fvq+TVXR7rHMajL0tAP82sA
+A9uepD0CQwugLar7RhLQvqBvmBJe7mhrceDuTo9nz/VvBZ+VT90ipvhiJt5
7p82oXF4+ny1nnRwna/4xt8bu0zeJctFm4C3gPMa+NRz/QZkdi67h134Euz3
7I2BdZ6QPjl3oQMevaKSdv5+cBP9SddYuH1G9BMq08DC81ViWdZJ3YZDu+5i
VZ1ZyYnRsJYCBXLv5NTnIJ/CWhNm7nldYJ3FvllJ7t2nNBPvm3WiAK7G14H1
OH9YOHvmM4umf4SSxwdEW/xmOCLEFMnWrsseYcN0d9KeEngfycy1Km4QduF9
9GSMy2cDpWSuxBACB/YFiMquSTkxQqqfOP5O2tSS3wGVMuaBtssW70BWfmef
oDs6jFp5UbL6oxpr9SWQ7Jr41vvlU0fsZtzrSJxMpn7dT1JaTxh0uw/T2YwI
2tzxkvy/aXZjJpaMI9DQdtX4gU+JYf+iB9GWHcYtdVfHIfb2OJ67qVPC75TQ
E16QyePPICRdzCSoOCBLhznVIrOuSg25RYZ5YTGC2DQElNWFb77IpQZZGNLH
j7VWlSy4oXKzzvJ68DpgFFDCJIZY6PTHs8IRkvj10eKTGmwxJrxKoQc+RmDW
DwHCrN0NFfLZoxlY8mJphfADgeMmTE5RHDk+qj4dVs6MxLPwRpCkhVw8A6Nw
zAyl6jai/+Od+HyHzcZGPGe/xGz8S7G3jk/p/AWn8/SdVCdu9aTUKkTgmevT
IrkYEzo7mElvQgNrL3oFE+rQfapNAuWh8sA6puha4yodAKyu9UBeS3nM30wg
yOZXlbGn0xDSJ94/MgmD1N81GR1yDBXt8uGvEmZVSsyq3z2GjFF25CTg9lZD
PB13Zdzt9j+aM0rbaVwnoJXTNRSyrH/qLM8awAMCSBEwzftvhG5B2r67d6z3
4H0LABW+P26bENAzL34zBdAH9n23i5WQp6vNINauNygQIBhkJlXYevUcnelv
A/9YaC+Xu3C5qZAblP1OR6mM64x2LXCJcw4nHS5q2ZY+RdXzYeMbvOlEY16R
LOOxeTIw/XnB9ftF14VuUoeqIrZ+rzE2rlnI0bQGQjMF+q1pzWEeEieAJ0DP
zwJ9Mhh0FEhApNSjnkLbEs/nOafPUn5b6kDTeB1RKadwva/VKzQfaiRUIxbU
b04zAtWQdE1SaL0G+oUEFnuTthsjtA8KHzJUfh9lpX6syyE7pXUTct/Gs8bg
YStXCp6opmyxmhc1gD524rx9Tnts1apzgqGlKlGOZHH8MKI3+gUjgdmLa5YB
8dOgWHYpTuTudZSs3mBAoV3YFwk4xS4pcrcFPzUHqoq/7apPdHCfFKlmtAv5
1UAnpFj052N2VUBXxBT9Ok8/mBqluujJKqyHMKkUt2qL6SOxI8hvU2rD2lDI
smAKntFjsXWC2SsdUVQlg4X0H23u6Ce3TZAhblq3KjZ3W/AMqvg7qZNRF7C9
ypm9xpVuMFXlHjn5BCKw7GoQpkg2+oAF6Z0+Fsndoj4SNzAnvrJcmrhESPDK
SCPZIF/jX7vT7rbHxtKOTL3kvr0CWh+D3LURN0kaMIX+PV98h8SO4dTavINR
ai6z6k0oXXIlv3xVaE8VXObfPswNJ3FVPvrKqP8ngziwJSqr4UVdvIQzx0V5
Gdot9FKXPBKLbyv4Dz6gyjQZlX4rJ+PyLt0J2r4pcpvWCMAY+Zww20Ey4SsR
ko1oFEZJ39+VVm4PJuj0wYv1PBdv2KrSzdtyeE3ucgLkEdc0M1mfblEZjf3m
mLKoS2BiAhm0INh6AeXAaO3RJnikMLSpOt0krIrqofgS1CkwqcyBAYNOkf9/
pfHCokqzc/01HxKjUPqYITgtxpbiLJGzVjwx3pdbFz3gLuJn7maLADdZEmPr
6f0EBEKUZOwOSJUU/PU44KTVtDQlN3Da1nV0ypcmgBTaq+mj6vpRuutFpdAY
7dVXlp3Hp7GGrVPMWZWA1Ht7uFCGNnd0JqsGiXVQhjmzVaQLT0Q2ud7kiSI7
RiTo7OfERF6E+DOU+jvVMu2VHnIq9ufwIWci9XtkR4RA0auz+H9E9yC3HFwy
z2dbotEjMMUG+0k3YLUzRRq0xMjuk2h0ZTUdtYd6reCAF0Y7CEBklfu6AgEV
0qVMvLQYiHexJo10du8/9d75vqmonXx4K16OV+AkBohoE3+Mu2w1XCc79ML3
o/DWLB+jm1twUbp9GnLZF6QYDrPJZIuWCnpjZYBIgq/hhUUtJy8Gtw5uzHAl
n4Jk3ED/coFw+3IBnvrreI9gtL6LhWBPwaSpw7y1w0HlU+ODVw9xsgARK0zI
1R104Vz9zoMlp5uQRW8oc29Fh45Vn1WPJpFO46Axikl3ewzGG3mc57pIFYcW
+ZG3ki6cCbX8kQKmvuYFn2qnc+/tyGk2vyAWoUcFky3SXoKM/wMHJnOiKIu3
4umMLkVjEZ3C6hhevlFoTcCmXkL9MOfQcngt3igbxr9gG/WAntRtEbWDntad
w2nYYQaEehI7Lo1oc7/aX1714o0ynbjTdQH1RpMYt167rx+0X5LGxJY03bC0
bxXnHp7ArzQS1RaOl8XqPgIbdZ8u84fQZJUJ8hRuZPeKinFKFf074vjVFrsx
4I6l9FeepJ6I6VgXySxyTci/RgdI4pPr7TX6PoJ+cOoXm4cAmLQ6U03GgYIq
Ixk9hSGRRG56o05DT7RRxbbbSjzrruxdogd4DSfv1N2hf4BNpMCsHCBoKOG9
FExhHqGe1G2/lZqIuuzuyiPrlcP88dELUFcAY7zGaZmJoWEeB/SPmkiBHfE9
IKth8bK4VfrD+bRUtliz9rLwcMoFnAlvlP7qK9VMGKEy+cUoNqmnoLsZ6tXC
fLE7cRavskgWcheNztNoO14lY+FwYEiBDS35Bgubo52ayp1fv+57QCSlavOk
D0gPFJxTfXqQf3Xgm47o6qvOvGYgIGDm1GqZPu69SNZVkllqW5AB1kVVzdDL
vZHRTboaSScSfrKaXpf8BoHz+qvYEDUfITy/fNI7hHEEvq1Fz5bTRSp9B1JO
eT6eR9vPyjIQ/rPXUHaZbzGt6qSNjafI8sxS2J2ohHbp3a+eydou0EeJLmyR
zxEOdC3ccEzy3c/fUnSBaHn+zq54tQ1fO1BX3g3YtPfpCSbXFx6uR/O/kmRT
+SWeSEt1yaos4kIDSS8+Tfb/aD7ZhhPIHmu9i05T63j5VutDBjGW7StS9x2d
EA4XXXma2t53Xfa0yLxa2QDOTXx5WjVvP4lxvEmlSGT4iBxFCuHw9lcEgPqi
/N39Vf4rDtdUZZJTQQXJ28AJex9PiJtIdZTS7zOoWAi8qiMkzmf1cD+THh+c
iQsL2Afmv3bcBJ+Jsx6WO4UTA4SVLiltQhB1T8Wh/H+rN39adie7qg3DOLxU
Ao4JqQfssdf4AgiatGPTSHHxOC/3R0GonV2a/n8f9VUN2s8hQTyxZhwhpDl+
5ReBldNIWBdi4a/sGGulx4/L9AZZW6Ddth9uUEny7hosBfBL/jWkGI0JxwSQ
wx1f5wWS53cLvdg/T7oVJP0WdhpCTCQ8CiACpgbk/xqpDlETo3UXu+9KjXWi
G0C6R9zveBnSXkinYWeJalC3ETfRI5hb2VfQydHXbitDUI2H+Dq9dKsRrgcA
cGjYDZHdDEksR/LjCrqjVJRHD4HTfSBgCqtqQvghFsTZ7EWfFqf4UaUcGcOJ
z2nTgz9iv8OTBiHUvVlHlA26UMRspMsTVuN/DOV8WsS832uzF7IIcyYwTASw
lPsTM+qBXeB0zhCSiPV9JazfiBEiztr4UZycLMK00iywwwlUKSSFI5OrLR3L
wvt6XSn9cyPy3cIIVPezk9jm1pyluYr4vB5GxuhiFbtmK/XGZfdo2eyI3sqf
K//dPiGLYDtFEgiyDjMquVaufqJhMAD4O8Jwqnr7E0j41lWUqxXGLkA0HzBK
gC7sWTApUDWWm+VrAkQ1mMLeQwbcYG4ufcPBFSc1i2a9a3igCaA8JrpgkV7E
CaFQJaGZsO5kEEIm1eOLvj/Q5mrfMgSvQgUXw040j5xiSxB1uNaCLt1OPyRt
q6ArufsAQwhMspA2DUs6MzU+zHTcp76yEsAw8Qc1c/6OWbDKCxISEX1j0ra4
MSB2uYEUrw88PWHu9+xlED6CeovXrMJGAVsXsNqdd74Y8yCd1rQIqbYDyija
NnCsqi3ZnsR4XiIe4VdRfaZEL0bWWu0Z086PoNg0FzUhVjnKtpPz75sp8cqU
pdH8IexACwolWFy50M6Pmsg3oWGtC53OfixiNMR+F/vcflQxKOiLIvprg4Dn
/3bFAZavspgZ//USPbxEkp6qtkI1EdORLN9ubNDnnQYXdpTOvPWrZHMV1skW
VeoB014yFnAvqUr/QTGAwrzvmKWBVHhNySKOeZjpBmzDtUL2kJwsMYZm+kaj
iDYShTjHzZkE5b/SLI/miDnHdMyS7KbrJ5CVejU5omAMSNVrgZJUdIBCyd8l
x9j34ujEz52wVgAqdY+M/+owIzPVZJtRB9XaVTuiXwzWrZWv75EormRJNoSl
ij2g4FCTjKbzFp/MctQWuKpSJU0UKJBJHPfMng+XJHOQaYA8JxtIUmhfDPST
XtC5RVHEnjJA6KdtZs/HH4FxR/X08BxDHrl7q/O/sD3sNs7WBbM+OLFCUeIg
DqJEqafbPmkjndTpq0Zp1fOMGguPyomCytrVbscU/j/apFvGm1vfCnNQ3kJk
zL5N3/E9zU/HIwVadtxCp98yjy+lJEANVC4cP93l8Ov+mXDDqkP792DFAbjR
/MZzf/IrO4Gya5Vm4fwwuZbb68KOhnJq8KzjWpxonR6Fyexfzbi22yrMQnCZ
MY6AWufsdcBWo9Eis0P+XvrLTAVs5DJaquu+NjHXdpNqn7jku6NeQ1oXRQNj
3sHhXQ+SS5ezsFOdTlnnmOAcLmY6IVqdFVpUDEXNIEYeO+MyeZWhQ6Pd1uMK
Y0ku9MaG/qey4v9/bnZtG3iLAc7BnBqVclZGITvKjcFy5sNBz4Sl003EnArc
jlusSK8tC6CqS5ofLPYU21pSnQ1tDhOvq6m7WtwA0je7JnmIB4rdqY+Lth1f
98AlMB6rfQVsK+QJeFz7mbacKdohhghzn7OqXB353CHWIFA4mVNjE8ZhhIZ4
IMTvMlSDQO/qGFMziIw6/DU4z3Cu4PZUSI2Gh2od6sJpbARPnUBLfvF3XYOX
UsWaI69u1KRKo6Ilh1gSwmbnroQKn2orNxYOcan4lwwQW/lfHG0NA6xKqphI
SvqWQdxdmM8Z0jd4cSl0W31Qr97FI81B12SGI60JCWEtQytxt+GpGs6SexPW
ThUk2MB8bOnzjP35UJF999HtiT3lKz4jxo+3V8x1O4DU8Q85ViURfIjSleWl
peOz2YDkJsQOkAqKW+LK5s8aA8K175erwnJcI6rSG8VgO6xO5jcslWARiq1s
8yM4OxO+diXQ55Ohqf6C2XXKhS6lUwDcmHbWACe4iUXXvgM0XVGJ3JhZ1KG/
tTw+TNduirwDW/ltKZN5+3Hhv/segzvaoylEWljlYi9BtQIgLC0gg+DgpBr9
GHoR9XqXYrOFD9jJSWm6hwXJbiI5ykxPrAeDD0MT+k47noBmKyDFGbrne7vE
vhYWzPObaNtjAsflArn6WkiYsDJDGM1hNe0JU+iggR4OJN7rsAhIPYtu9bPE
RxRou7DGdzJqm6y9HvKyBSz2lkTLZ5aUcYhW7k3WbmQNbUcmgJrY8OOdCg9Q
+wy1B/YHTGbSn1br917D6EN31WBtTN8STUIDgQbUa+JkIhwBZWJLrlGL0uOm
RvffS1VB95od/8PMQcgnjcWBCm5WF7jpvonF72DDg+qXumcWGBYu5TvbKeN4
y/8+Pc/wz5/JF6AauVylGNJ0N/yUMx02glJ1zH6H5PixzR/E2Y7IHjAAWebS
V7/ePiNWYjA2J8ptduuGdAqbWS2BpIXqKxbyDPvNW8eN7bhGUVYRm3VoRKGg
XIs4bBuFZDUFQ/Fd+ow4SX0veo1nJ/vAgpU4XZBq+xQHW/VjMUId7Dh7K5ma
eLlu5qERqNMBzEYBe5A2wTc1neg8WZEv4sWhrgymzKjN8ZsYU/boZJfE1pqr
4p9o7F5njfhn2NVj2qfezdhuUKVAOsbbTA73dUbZupjCKGTGiqTP9ivyM0yJ
Xw1D38wY0IA91nQR+dSq7wazePFeJFVr02s7vqQVr0ZqZJn51EZ5LaCtCNI9
X3eCG+dfxT2QWOFWjDCwLRbOiyJAVyXjF3q/AX/6GahDkSbse21lSSE4Ldml
6/jYp3TDBWkZyaynsD7+8sLnIpvuT1e5j7MRpwM7uyAcJ7ePUOWo6n6loeWC
3AN5mvjScZyVvZwkMTK7hnu1U1SaWnDdHpEd1VTP5SFKawGgLD4jTshQta1N
MH7ZSeewC12jJEJfwQ5d/RwJnBn3Dpd72bBTqFkfXGRWzMWc8uMVmLPhE2aG
LEn5jG/AxebDl05ydiA6AAwqc1U/HtJk95toC9IajF5DtG226CLiC6SHz2XC
rZ5sl0G1GYaunFzSicFpvAeO5JijRZCkHAVNOyIn4iWFSleWxCDtbYXsgN+C
qzSa4RMMY8ep/x2paJ8gp254ZKYRSuq6gA85ssc5WTg9fzaDRXlQBJeEaJCe
q+tGXnwzDUctzK8+71ZS8IIRtNO+Xef0uao/VMu3bM5cx6MTivNRvz7B385S
5z5hS1BecJkQOfZVFQcMlJCTSvKlfzsknCIMPsvre8DGUC4basXlIYUY5mVg
AGyfiEM6MhaAGZNSOUA88+4syUmh1Pj2HS+5vYCc+5LzHgbMDwKrEm5Fep1v
ERPYoMdCzrShLBG/9UKZMtMTlxQpXrMEN2b6RmlMM83outMjbGUAvE0Lo8KR
gqjyDWsliDhW8YkRsisXaIDPYhyZZ7b/THuEAzXxg27Glv3ZD8VK9u5F/bVI
NhHp9CdEPS1MaOJMwKN+V6rpzwsIkKIUAhK/+bfDyxbA8N2G5Xw/1PT+Kbps
A06BJXENOxuAWcWOf2pdZOeDGgWlxIEtkbXMzpZELpDSmxTkwbn1FaY5tSRf
CGTm2TG8xxrm4r4pxLLvcMo8GcDEHXqInHabbYsFzWMFhFNJEb1Nl/vfe7Go
OzxtVFNlTobsZpKi4SLTn1p4nhiIUvXuL4FRQSYaGDrc8OVJVw3eaSW9euH6
uSA8rXbxtx+YghWXqMAH3xAaLr+3ZSt47TTMiQD5UAkSb3oQjK26dXGr65NX
tYFwMVRUKgER0aoI8sunyGiVXtnfIfzw6ei/lwHBCCq1mXyCapnYP5Qbblum
dfmfBK8TsZ1QX0zJiGxWu3aNqA6zC/EjcAy5JpkWmfpz/Kbt6ULaKsJdnCYh
liWUqMh/BKOy8LiAOZrizDY4VmGk4pcLJJATjhoizwSyw6D3uOn12in5fpD0
ThfDhOCcK/fea/RQ7B+deWlbxlyyBg8xXkMBMmwASLjXhIfuefkhHaSxTJNy
cdzEbgREBPpb5WX037WtADo5qhzAvt+hxE/I1bs1RvKeALkKyV8j6gQe3kgA
N4mXAuF2F5BbcRO35N+unUxCBgYvU/vcuOO9VBTSdQYMgPtHF3MM/EpMP4I+
ItiIX88hgtX17zFk7DxFDKeNfPpz6B610s3SQxds0/AhJLlvwOI6lru7E9es
82YMz5LNa9gpkiPl2GhpM5YBoDIuE6Yn+gCibfU4RbeFTjw6LfunXfmyP59k
bMdnE2tU1x7pium+Gir3mCXzmRbW9haUWRW5mSvPg0sFM9qTWHJfXGTp80Cc
a+KecfC4y7JEKXCHjaPhlqPDVuJuv8DWxqUZ+zS0lcm8PBS2FU0yO++eT5qi
jFIjAcGjWwlvleaMONfYS33H2UJ6LVATSBoD7V6OaCJrmuVVTFhB2FYEDn+J
smWH34GEjxkimQsg1Du4zEb2JahSNcMyJbQUwgGwhRBW0ZxZRsn1aE/seXoO
avalxajvfrPYpdxGG8oKMKhiLOJYsK+oACoLPjs3ylSAvW1a+3IrcUvujLLL
/Lsnn+Dn+Ifj4CrQTR3oFR6PabV0MZ2ccsr5ABp4/x+k6Of3is2fNOojZaQj
vGTAY3MPjNBgB33JnD4G37roHjI25dyeJn7CwcUgwi4iVJ3Oc2cOw8wcWq2i
u2TBVE2FQIceH2vXEeyjL6u+fdJw3YN+G9HZtkmHU18dcKY0TGHjvtAvbSnD
3tKNVMcexH3I2d1ifa7nXKrI0MXlXxErnNnZwhSTuo1jyRSGu8NxTjtAHP3T
ZEG4eYt6N0gHv+n40VzGOhb1grXGoysSLcldJ4sqS9e2jkTXsXnpKnxOVwlt
4Hw0FjUmWpK5ctfJ8jlK50moZzB+WLS+7zBI/M+0VsMt2txc+fpL4wXevRaK
EQrU7DR6mu82jNHB6E+Zhx3xvPS0PVi1Y7e1Dt/FnNPIdayDv1OnDqiFRded
LYDXqPEGe0K0hP2pvyBBML1gwSrXPmR+j3m27i/oQvGLZ6ennrhr3Afmr8Mn
wBl5aXh6/weg9pz11W5vJgMmYUQzo0oim3oTkB+aHHCm6PNtv79o8GFMOeE0
xEczqMuZafQgQQj27xIyOj37FjdSr8LzLUCzYZKMeBi07I2ClIiQw487C/fr
FxVLodAch53LTE5f2tJUbYCZj9Uu9v0YwM18eJkRjtfz/GOSgHmBYgRnf+gm
xW0Hnzuh7cc0chxcEAcKCQvKRW5TnyPqv26MyAcv8tKdjLGZn3WVXjwEzxtu
yhCjFZCwrm8jKBsbgg/6dJMJsiPxAZJbPXolhoKoZnUqHZf3eM2YGCDguLrr
sTkWDs9J1PBmneV2pZklvQu8tNON1/i8djMrPJRpwKjVWzJodJLxWtscD59M
aNZTTur81j6F67ZARBKxIkghhEkxtCir/EBfz6fkPETYD6v6LyX+kuffELkZ
yN21tx6f7NC7uwfOsVo8fQCJuIZf11Vo845mQVTEu7TU4osB60LCyUoDHvCl
pJcIjwuQOIiVvKQRJ6kSFN+j7YzemcbfmdYlFu7PuS5Ax0I/r30Jp9kR11j6
Fd0PfjhwHtJmGmpJNLdp3Mcg2Klze+BDHrkuKD/W7X0eSeIzUj8D+6pirOiO
9RNZP5iABS9XTIrkKukDiurplF7tGF29h8Jkw6pwO2B8oNfFFZbIlPFEP5/O
870PCzfZsvQKYAP0v/pnf+zNqnthLSE9Zsn+vhHJl+D60MKo9a7KiBLsmkCR
40g4mWGU9uMuaXs4xzNQqgLEDpbYY7ipdPh+DZ7a/tsaBGXRzNMA3HvMtmOd
5NUNcbj60wcy2NV1GsCJnJ7RnmoOcsRkr5Dos8t4uG9JMpyeFMiZQZ+tdTKe
/EJnWJyKyC16jDNAltqUzRCM/UnqrL+LUc+zNuaIo0Y9V1Ud1dn8tN/CqY8h
Kib3xUq5c2pP2mFYRJKVj7qr8xBgBaNHjKO6tQPaWiIvcklFZDrMfA595ipk
3odeASXA6IBs122MxwgbKcDKW5SrgrmQ8VmmxuNMQOsBlcgHOgkaBgXnvObN
HBHZyURRBa0Dp2rLQVG6QBGRK9usA8/4adcuM6Gcu029CfnLzo2HuY6+YjAI
q7FT8SljZNZ5IF49nsms+a+IDiSsRGj+rQ6q8wmnHU7ggE+rXzRVLY3IzTFn
pGdWgP7B7vEZMXJYmcsAPD6DDzb8Jmp2MHET5nn2QmDGpSmt/wgNrPG0S34U
HaNHITku9COP1qN80BbDdZXK1Xw/u/yEt/350Di2ny2WonMkWr73ykVe9j9/
9dOyMzo260gU86jM19YRgcvJ7Sy+v7yYpkeD5jvXwf6YAZkllr1pBGzlvTzi
Usdw3c62IFWT2AHzOTjIipxfPB61+8s0wz06rIr4rb28BeYRIfTT2kg3wI3u
L+FSDD/kbaNP5dZYIhqXRBctB51rIWHFOqO5SsHudasRBVwzrQsDQgLabL6I
cUV/GgbKDmdG6Ig5KCRGVBJ5w8BRP4BLrC0naA2zMwYW4+sd5abObMxahOXj
9mA7zlSNNQoi/YFX3TS+0dD4J1iLJO+/SlJ/qCLeKepSz3Lv2K/bLSgfkbUI
bgom+4c0TOXzWOseE5gb1wTkNwbwO6Bl7jNzmCIKYak2UcNCGJaL2VWmerLh
zTtv5qQDyiFKvNaoQ9pRxCKdaEOhp8HC22wLGd5LtmGF4mNx6857XC5WwaxG
/Z2/qKbdRdTpZqm3TVz+DtgUmq9JWlxHeytXQSk2aZ2Pm0pyl5auKfWOGC+A
a/OGWeu3r+EcKhfbwcQfsfw2+u2cEMAQT7xVDINlRCDh5ZrkC0sWx8XYufoF
207FSM3uj2LDoP+lWWSwnmsgLIcDRfJzAVIs2KS2USBRLKjpcPPxm5Tr9QuH
2nX3S6nuuYMbsf5j+TgN8gioIBd04Y2REUw5yPbOg0cXqP5LEoMAprseFgPy
C9KeiqOtPMJ54YUuJryfseWwTDqwEa36a+b77VMrFrfnAVBjwa4On51JeSZD
oTtcrZwjwh+IPaaxyuwniFObO3V5umF+QPzNon6LIgS2qM7eA3A3/WeclPgG
MR13g8xS+Qj2L42duSWs3KFaqb909JWQsM0IKs4Zl6Joa8I6A0IrE7ANZr0L
6DX6XqCg8JFci1Anaq4UOJnpnBLk863/QGwDhgjXSquLFsZEXkw668+8ehpA
16Z8a0fEeZZhhOI3B8FryBeD1kqp+5pxJflmE6NWXiANAJioBwHt7BgYF/km
PNn830bBEmHSHGa7RG5RvYzX/Noi75mInmWZ4F4a0yBfvIOyt7bPc8IHr0He
571KT6TjNdHlrj8JTee2VYmPV/nJiWBQcXhAleUenirGaBe5cDsRDym82QZ7
xMeuVdhkUDVYtyJdjgi2FGnE1wc8RjwdOT9iluvftByPw8YXKFgBiiYEz/Wy
r8s9rKW4lgUotj4DYdQUbQw8xO9HM2hqhIyZjku3l16s5LH0HRHe+fhKoYOh
X//2fkqHHwP4GHUB0Py1yal9+EFyc3pguUuTEOlI5Ia0+sJMadYmEZKgMl2f
615q5/R/j2PWzCFf34It/B1D+lNHCEjJazFKIKLrkEsfmcVMpIZlaJefzpuL
Y1n5goMh8SQ8LraXHFwP0pnRdJSWbpegsD5QpE6K204rvx1v7YhiJmszkw/h
cldUsQFeOfsgRfzLRvlw1Db1o5IEt3X0Xi1nuX9wMbHojAUWbBkNxZwD7m+B
jWshukRgRGykmU3P8oY2+boJEp6G91jHta70wgooos50qQaBsWXgtwImtRnf
2dGkkGg/QbmWFvbKUofG41ulS9/8l3PQnf83SrLbpUF5liNP2MS64UdY8j1K
gj2xiD/CH4kOtrkKTSOyeq0jMdzGPHhcI3x1WuTRZITV42Ba3fh6CfHsyOv2
8FGj3dzJHCkA7hOqB7POzk3Jd8uo0Twaa76e/P+miJibPyhmFZi72VoFwpSF
Q2t4JC6OKTC+ajE94WXAjZN1WdHlFbNDxSY75CDyu01CV2DmzKSIlA+eY1JS
Ra/5HblbLD8XAzIr/WHuwgIOopDmFli/Aexw7bCpl/PKLejxv/8Isx/RUQBL
ljP1YlP8boUH0ZR0noZfSpZTycGdtPhNy6lAUfE1YlJv7j8HY2C2DOhl/jFN
4+zWezqaaeQnWFZKOk5pKH8uo5IwbM1gPvvpYD33Uiwyk30653fGyG3AovkH
2lnqLbkIX0QqEdOBWWcWPThIajQPUznmU+PlCjM3GJzBIKjlEaWQp/G/Y1Rn
DQcNLdeWHmzNRvjeIyoqvlJQg6dTTk+rbUNKHIev8wpGta7x8dBhZSDLjI9t
Zc/rHQiu/SqZpn4OkkFaJUbpQ/UHU0Q4OJL0rFHmeZ7Aqxlmq6FZNM1doghV
xMpexwzwHuVQD2JQ8QsivStJskWNvX7XAnelqTzAmHRolGTY2/UfVYQHcBPu
awOMXAmubTP2NaIRC5xIxOWVdFR9Q0Pp50OCQ3Zif4VVj3nBScr3S8zeyfK1
PFQI/mRtRK5GBNsfBsFbf7gNpYGSryLxqQj2Bee9O+4rSZ8C5pLPswgRm6De
2JEZzNNwmOM8XA0Bl536XGLeCRmg58yvxwsiBD+pzz/BkRs/QUszF+XsDXVD
PGIwVKSW8S/bnFYwmeA+QwpL2q57GlFZ43BoxNiBBCV6OeV/ZK1R/xAAZO0e
iLafZ5JqTAqDAPTFMcOzsIHt0SU8XaYYnpa1Ceg8QkYyIfqf7jclVOxTXtF2
i3xLMNt8GPm80OHrEnnzeEtv2oVKbohWsg5aWcLbj1PWl+wpb9ZDk7zwDFNp
ET3+G9s/d2bettX6DUCiq1kYYn7rfuPkhjOLbEEpiCpyDqj9tnGPuylVCYQ0
Umv0KumDvPTW/X/V7zlwd3kUhjo/daMoS9HDMGKHtKpKZSHQaSQCpJIfexZa
OWJi1rauKQlkS7wefHjHx0YfeuAevhNV0ohAMdSLodDC8nBS3kGb+bYtK9A5
Vrso2xoy4JlZA8OtR7z18f5jNphN0a052pRHno+ttRlRv8uUa0RXDxOYE0Vb
uEL0C18mUgTvZCa2OnVw8LEYPnzklcSMm3AD769ZDLowU42N6xGG7bagFXsJ
Tu9UkdqJYsdDD792TAtSSHrwcMSl7BlaYxWnKzK68mgdpri0Yir9iDrKA+Eq
mPym76nzqYfeIg8vT9z3/ajZN4hHVRZww1M67Dgi14laI36oPSgzp3nSo8Bx
ad9zetLn5Kn/qg0lkOCZIYcltmbWaCkuhBXwlF9Rsj+klTbqN2i4yHKo3Dab
YsoHgCLNZgsV3RAzNQBXPnydDGkj3kQyC6eZwJ2heiWu1RjJBRC4r4KT7Fp+
xRQjHrEWO3e7K3WCwzJMobjEtQPTVZZk0jUw3KdexcDkstT76Gdv7VMw+UhM
TkScp/j4yj4tHPxk9N62ixmE87rE838sDtlatp5Ly5FmkMI4h3lTHaYS//IO
AYfqwkQN9E6ewfFCBw0Bp/UBNJIej3CvWYHDU1amUYABU56ISsWXmoZ40w6W
/6S4FfmXoMvfbfm2t8S8n47jC/py6vyIZVmd1MNEFqSdGJ9dkSY74t7zu0iH
GR9KRi7OHa7XDgzdB0Vv9YTEnq76pmJjwovsAEy+o3g/oveiR/cVGFNbbZng
kfigh/nUj8eJ9IRuqRm+9axZVeq748M2MtcvZ8Q3vtuCLD4ogc3OBBv/N+LY
i903LWnYclYSL68p9kniOY+OL3woGiUx4/qGBRgWeMr10/yyKryIWu6HbS/3
EbbVS25ZdIHS1abCvDA0YPvwFxOCeF1fTIhIQ+MblkTLmVzWq8Gh6AFYIagM
E0QR9uy4A7eaEuOmgGg8WxXT0S3BFK5QDCwN7Uo/H5noyn0yjN3lGIf5W+A/
FEI+SqdK9rbQAO0OLZaD4BIhm9h83MsvOEix6Hd3QHIZGQ5CFCsb2+F7JwTk
IR6vZivpjuaYLa8fZB3zuXKyQoMTvXRleutN9mZrsnDuKXozIGlCuJ+u7SBL
KMq+RcidfxMEcH47OdeiEwmtifp0fd7Z+6q6LFXIvRvJUePycy16jgamjQQu
pNDs5M17BNKRivoN9e4uP6X9wZvS4tUpr6HCBUoQX6HNnapxt9oWiqbssrAA
X7RU4Ah9KdVLr2ocUQXKPYpTmvORqJtzasNCHstjV1cFUuZhyVc8mo+5GD2T
B8zI8U2fFSqJnbrKeyteAHBBI6ST2HSITpucyVJUx4UAwpAiKIzNBGBW304w
Cn0dJ0HSSF2fmi/JFzbxyH8POmvmC3sdRHIUchy1lm+8uPkAkuBpuySGGbVv
OoHKGLAP/oQOxnlJMA728FSkbbk7N2XpvEiIY3TFkmoYRPMWewpxYgQoC1wd
M4B8f7agF8WWt0YvnlWH82/PUmeA8R/gKyne94njdzHkaU6MyPJGaZifEC0h
9ZrZsi3qqoor0JLcZBbRz0ufQ3xXP34FRP/AAaMsr9tViEwfpZA8KxiRjnxq
ls8zIiF7lyHUDmOCeT2zE2Z6z8jPrPAEltsk2MYQL8ToMoD3+L2ai+46nSg7
9AvgaFbtINa9LqqToNRFaQkGA5j+WKwwcnSkkHXUbkWEqYjqLPe1X3FjrGW8
dJBmVB1xjkUpktnUvRe/+HtPwtG6/c0NEcU8QZ7XagICzUxuLXAGzlvloFTl
+a+intMbKfBwHUNCSpr0NCynESCj3KJa0dK/cWdyRblGITa6cQAn336xN9jn
SLF59J8lltrtpEsb3Enz7q+BqHEb1wScPIpCAEJolj6XuG26GecPXVdVrEHT
dqSzSs8GCjMOg7ecuV5bvFiLIhr80wlTyM4yyUM9ISy6gHp1tp5Y/emQbj6K
sxl9hOEtLewO+1+fC1dJfIqbXX8Qn2WvIFcr1wuWFigxtBB0gM0nf6KQEDu0
RanjK74PVRj+bWUzBkKzrG3k5d++4j2zp1sdH1DDml3NcM2Lr0jbt+4sXTTL
8a6aCAmFXAs+InTMcF0RnYaX66mxULR42KgM1II1V4vnjWTSe5vZIymA5Vml
JmznBptHg9td7BMvsCOavhSaKRlxmtlWBfYZ0O8T/n+JbU3kH8EfKw9xj27F
ZpSbmuKLpWmTTWEN+0jtVoskMq5DueAkmvDyLdtbom3ESMsJM7WQBtUvLhfa
hnzSzTW19u9y0iYaqXUXHw7FV3rAZYbn2FWrwN+YJrCsYnYEPvx+C2w3c7Nh
Ib/3vAL8IcdyW4hUxE/orXZVpxDsqy+p6/uBkLdJ9qq7ZVFMgU7bOp/3YUJN
JgTyu7uIaJzxoGLy0k52PcuH5a9KzdzSS31xcjniOjIO0DrxmN1AYDlMS7C/
uP0V2RcpFQyNeqn84G+Gqk+Z/HeSvErfQjJQjASp8A3FQJMiNF+RddiuzGBN
tV8a9xqR2v47RszaLlciYTwaiEHh4U82TNyVwEZsFw4zN0uMmNEpQOt/Bu9o
ZiBd5/M+o31UapZivBF5Y+2a460539X2AP4UvtbmhmFNxrPqVO8p016AX8y5
73K95VP/q610MJOxXJdj3GrohBVwGu8XqvtvFfEMNVXj5/GpXbTJ9MQcCA45
BsSpR50MDGMepUbPV018Ou2nTyqB6wGzSNBADorGcH7KqD8H2/zgMx7+5i5i
GR6nT9THt5v2jmfdTQ0MOnRue6F3mhdQG+FmOLTjthRZFmsjQTkRLGfEM6Gf
GCuDJmPeo0fYUNTvNZhZpbsQ9wglwcJFm5LB37On1FUkIMKZjExmlKqW2Yhj
PmQHEnn6iw0/fQJUS+NEA9Qgcz0WNmcDDGXNCPAoYCQ0Mks6U0P2TVU4M8R6
Rpz961MH5YXX1LHQpiDT0QQExUS+lQUNJf2yu5ek8yYiRx88ZH2coZxGvP4X
o1klTjDqJ3gwLm8GLroUBIsZLCYbJr5hD894oy28A/gySunT03g6+ohjAP7k
NMXSj4jZ2BUqVwLPB4G7yLbwDn5O372OpBi+l3UjLYl4Dj0YHDe9J+4bGV6t
mCbiVsyZDZ0409cHJ8GOv3jEg7fKJvXzV9gl75l7lXnG22O+X5cEkV4PS1Uo
c33M0a5Sy6aiGjJGKYVOfarxzgsoLbWCW07ZvrJQ2Nuzah7yQikOWGnZGF58
rUrrJ3MIbkbi6yzXd8FrMNaF7rFMNfaXTQTq+97L7HOAVJ/81YBn3Icoynmw
2efIw5ebcDIIKmDvRZfmYs8vnU6XCDD4b0BeLAqG7VZDYNX6tB1yeUeRLzuC
//6M1e7zpABWE9rD7LfpNT4Zjunbfo+3tgc+qOuIs4zHKSfHdn6RgcrhdFSZ
K0i5hQjAESsvUjERdIwhgu7DqrJdRJZmpOFQwNJHBhyBPgUridjiald4OyMW
5syBr7eyOf63Utkj6eksNlfWXp+eLdbJa+GgJOwzTcRlOFadbrOMJteu7pr5
KH+bR/ZNbhnOiNTf1uPa63aSlIcKgyQsXxzbSL7KeiDRPMLqcUdGkb3jxlsJ
gK2yoPLJfFjjmMJsYEiLjnTxDi2fk4+PjdnFXsoLrxnZkw7TkByyTN2sIxAO
RaSPxtzE8hetUNz83Q9qT1dXeOwEuohBJ0Gxw7l4Jfw9bF+SlaImk0gOd57l
MK9MiGoXyAvlsPw6KCGg9i8UwO0MWk9h7QMDxaLLHJKLHo0fHcAuc3smpeCH
MD2zAaiobK40Wix+dHcA7VKcfyekiorBnulkcKlbNAlZEIoec6slTm1hIAwz
RixEsxhHgOqqFcx97II12iiK4QgFyH0uFbw7OD7XxVjCM/Zux3aQlhqr4lKB
1HE3HLRL9/Fk1pYRsq1OPLkJAlkh1H4sqz45+Zix6UEeQPwx+QtLhoKPEqkM
vpR74j986/9D/EKCVhRrotcjIEdSvH1jTIzPWaGFW1MCuzGh7UrMR2sM3OyB
gUVxtxk3zPmJwbciDigfdouwysHb8wL8VLAQ8EPu5bi1PnO99L5hCrcL5dio
qBJy94PjSwFzj4uJY4f6DBGLK0URqrCqq8uR1Q4x3cM3wL0ezGWVOcVugiAT
H8bdDql2qt1hJq0V/CGvbKY/YbVAiUxWfIeLU5Ae83JlPU5wkewHGUmH1tEj
bZBMLLMK06M1MJs0CbFoDrx0f8kQI3H6esNkc6QRF7VduzznChUboDS7CNpP
tBBXZe+deaYU5OZ4/x3kCzt4y6O/6rQUkgm6CzAwIrRWIi7j5rfx+g4NN5Oc
sN2p632hk6oonvlGD/tD0Ps4lk1xFmcprn9jvUgNu+IVEj53iU72VDm7Sjqf
Iehs3dhJAGCJ14xT0zuPgUjTuYG5GuGrr0eHcMWFWatFchC1YMW4lvHljJJj
RnZLochhuQVuZwOs2JExZOTjzbv6uCcfAee8um/pYuwYnPlyf/1XhUHVtrKd
0SW6WkFZ3bF/oLrm9wPPEWYPVZZ5LXh/Sg0txhxPkyWVyeqcIHxPHRi73PC3
910mJN3YwvVETw7dgDukIbY19C6lHUOH8arrIlfUbcKiLwSemsCQHmr6T9A0
wGb+ytMf15g6Ltye/M4Zki6msXcaPl6+DffMLZThI+mYAxARD/xSf+idqmzl
5JMIPsuF0FwRPkelnv4ARixiIH4bKXwzxgeZVBdKiSc+d3R6ayQAe4AbjZ7O
Wb4g4Eq/vErNDQUlLw2Y0XyXseq79Va7p+VBIS46tDEPV1gZSzRrTdMV+WP3
zKFzl7DgjUcqTW+ucp12+W05SK7YORNI9uxCZyqZKp/P1M0jAmdGWH/gkXzH
MJk2Fnq0UNQIeCaNzs/y99MKeoxpl/0ZUxT7r69c0du4T6u+Bb46gB39jJdp
H4NR009t2fnBv08+i4dK8nAI5lJgkb3gLAFDI6FwYVpLQI+bew1Q7LcnL9iJ
X5kCsBXYCBFhK4kdOHZduGAYUsAXbT6Y572+lkgk1Ntc5H4odAgpi4rF9dFl
wKNZAKZBWlFFQGIEhK7SlWdbqXJgYgTOddAxdWuzGu3FLluz0SQOaupz+AgY
Xc71kzl4YwsK8fhrYpmS0jw/iLNKb7huRQ818WvA4XGoMtPxgKo9ho2A357M
qSJLQM1grUVs+JcLim8T0XwpoQOg7iUtqqoqC6PvYdTndZ4JgEPIzSDuYGCM
hlIrx4jAxyz//3E+V7dufXN7ZS0/0pzoJkMOPvvSMU/M8wzDlFd4n/3WVZrv
JdqNgfJigbZkDBYzKNgnSHcuXtQWn3HYEwfpcSCZLt8sVPInrlWuxxINYZqi
oLNh4Z9V6Rk0gwNQFMn0Ug4QofPj/mnKPdXKD4jBv9K0oD6Lo74vAdhuDnvP
0Ix4ZKjbFg3xSXc3MArWwh14WTfq86ZZ4TyCLBY58srY5OCuR8a/kZ5AkpCk
N4obp9qiLDzq2phuh+uUPjzu7vf34V5q9BioDTffQS4JrFa/bDGlsAzK5tt6
WVEIEI7lQ7hxMkYg2ecaWiVfOno0HGKCidFZiDtBX2RZ0S2HpTsvJxrQ/jyP
N1oJrUowGGWtxtbfv66cOumvnoGw5U3fJ4nQyf2F/WfLhAglywaUJsfPkk3O
3iusAqJJoQTXl20ePBe+uEFGYUHdYkMFNL99GaQdLbdxHzicHddWNHOq1U0h
k8M8dU/gO3U+GVWNEb5MuG7bIYCL9XGP+L+PzXw5YCsk7h6CQDpNKXt6wv2a
Xz6UrgOD6GvUpHB7YzreLKaIhu8EY/jWmyqNlB6YS8E79o9WrzkGwagoh0/Z
E1myWu9YvnabD5RC2HAsIGqWJHskHAndNZmNdWhHhD5vXOKARqh2fd6l0j2b
vnEauXTxI1TKtfV6/SKS5CmUpmrI1hes4ZjX/beH9NGo1/qZXfDjlMlq7PVU
s59Rt0yKVW20k9C9ZqI1Ys6lSjb2yQnsaJKrstM5KsWvC5a12SvVWum2EiRt
mlYkSSckRxZ5plm37zcIr2t3jIuwMoEJAXdYmhpUmNYGcWOYCB9ofEbhfT1x
18nxs9cAJgGwRnVMPPRvuhep9gBjyqVNaaGCfmDqXukCK6ILov4cCJSr4bCw
/f5y1yV7KShc3LBvn23TehN4S4zNjykOEuP1ibEBlFbGxUHJAPT+8g3AZ5Al
br1gFU+p9hrF/2+k7EzTSlE8ybYGs/Anp9Pqsyy+W2M2XYxSiSvubqNyvdck
XKBV83lfXFIMmEbVdLRwh/shgJBcho6zKCq6BkQEmnCAeO2y2D/1LOo71+dF
qxmOiIuQarRPzChslW1mCfbYZvZesA+KC14FAz7e8jfaIKkPTpgoKZNGA1b3
FlBhCMv32UdfQjWAadCkgiK+oMlxHnbqsXpV5r55ehDr/6NfcIKyy82SfZ0l
TbEkW9v9yRoV2tfk1BakaiIwN33b3eBf6VI4RNwvWyrlnopkChxxD0tmaUhY
pNEat3iYBpRiEP7tdZlmK7YYeo0UqlU6L144cdcU4D9BQPlf5G4h0IF056OM
sR0c0EFTG75I6Mc4Zq6XGZ1JJ8cnvRYXg7dfJoLQRBaDFE4C029V3mIS6aU7
XcwUqsgLazBJU9bUxp97H1uoOEf72dxqhcfNteM8AV6Pw88Tr3GRjyvlDZ+Y
gA2uDi3qfcSMxg8m3OSmrKt7QX7G3pjCj3xAZreVEqBJZfJqdiPDvYsB5uhA
v2USCZFr6uXZQw8n+LZ0Qw4ms6sBsJykChNMFX9DolCzIvvLhzti5PjT8DDX
lGLeglQSxVbKJM/TVul7z23ah10/M3rylyfDeq5icYTLlljJHFmKjc2uXtlH
m9bcjBa6KhIvszC2JL3PJQtfmeeNn7xIo2MvuE7GEmblntYOJGohxLiDzKEd
ChgcOMU9MVJE9Thz3BfgazLv0vWVID8QOeK7VkwhCd1tZJt37NVsu4/5DQtk
PFi7li1MAbId/+9nAxGq1yF3HOB4GxwsWToRozUYqu6FQHc3sMTbhGMAD5WR
oTM3NSpZUHxfR7qE/21TUI4oVdP8YkXwWvEo6XKCPLkVB8J993vEdWASfqUh
Jkp+ojTkmGLpJW15mJ0UU/DE0bZW0PTiTmOcD+SbVL6g4CH0UwXmdXAb2YHK
tm22PqjI5mVapDC3mn51h3EsDoJfw2ZgKQvJxy9eW086BaeHkpBD3REeTemC
9T4WvFvbdWwJLdnrtClGx67qRQYg4J/sXifCekKsP2SnK2OdffqRJG4jJVBc
psju9AH2H6AFEwGhoEWK6U/zbtqayHQcaeNFwKOAb5I89v3zrjXbSUXVsYPa
DPk0sbXjPah6QMzWVGvhDyhIPRQ3yYlp1tYwZgW67jONFZ6jrUoziJVRD/Ro
/EvQqorCIsrylUa36nc/uQ4uymZzqa0w9UI7Tp2aU7bt/IHh7aI6s5gg/i4X
+96C1KF2Kh4ilJ7mRy5yK0MxE50Gy1PSJVutzfr7owkgEnuc4eMftrizewAG
YaK1k/zeiLe4uQXNW06Uh9197QU/gWvCCVzSY8wOvI9LbotnUpgUkni9H+Ma
fRRCiXWaqc1wNqRpoAqnLu1R31m2g3ZJsQ28+2G7bBc94GTDEVniISEHpznj
KoVZGYnIfSILmKOY/xRBf0/2E8P5sPNkHXkSlmeEMcCKSIR+Y/VbEu47CUo7
V5l12GiNY4H7xFUYsrPTY9rtxyoTDjOe1iNdEvB2cfE31rZLvFVbuV7vtLEG
byE507aUaQIt/cbTOhyPksJFLpn1PweGtB/TpKJ67Pp7ovAn05l7ouaDw0e7
3EFxH0brep4Eh8Tm2XQ3RmhTk7eJgxQ+4FlOzXk3yj6lhk7Pjg7JD1GrCodA
zlF9tw7Fwu5ZRNlSB0rtyE20rv+kZrXkB4d6Nm51l1XIVTkIsxPDNUYkI2km
gMt6wZfgj6RrlG3na3Drf8ORtPG/QxOIzLzgG4w4cvL5uuZdRpAOZyrCzELg
ajoRUgr9P+DS4Oy+va92VxQ7/efTEWG8lORdKaLIV40651m5K/YMasLI23OY
q2IofgF6K/OXnJhajBmWztXRNec8q3o8G4RRU/BDTjJLe4WfGYQ/nAz0jkOK
RzlG5tB9meTH56XSafC1/cawoMuM1qFUSJOAdCCAGP94WnppweaiTgIrFZSE
sD3/M2qsN4rv8drXjD0nRx24Fgbj/AMHIDEWnp2JWYvqQS9pf9lmV511ytWD
Nsspf8MylLB6fJ2uO6siOKoVDSoF3TLrjBEhLEEGTZ0RttVNhQrFsMuzT6sy
Zj+qPrlWdXwTy5c4eQ/IBmUeA62BQV6Av8RjoetMW/aSkxbaelCMZY13BjQ6
5/A9pe1usI5OWncyNDWTC9W0axYH9ePJzjc07ld2dQLNtfy8MubrBMm0IyWq
qOOiD3sqnfHOq1/SU0W+uezZp+awmrpIcQS8nnVfkcrE8zXc4QIhLJAc88N5
ykrnP8oAzHmKVEhyZuGtMciA/Q4gpC4RVyCK5wYfRaT9hNqrtYvHY3R6qZ2E
2Y5VmEhAHUGzAeAonU8GKW/uJ/Xen/1j1zvq246UWGmNrolCR5lrCmWOz1eo
qvsnF6ZdQiBG125ADh8u4VrR+M8ASNoQHHeFCXBCUyWf8mVLm0a1d6DlOiob
P+jGcy7+Qmh/zJmyeBRdnEFTIReAwOeg2/AIHOXZuHpr+2lRaYirDcOEbgwB
6D/geOSfa8vMIUZnphCZT3B0re0152mstDunSfSKzQrR/y8nBUNlpzj+PJdZ
xfXKY83Va1ZTkX8nJCtgM5oNnrLP5l55i6CxKwQklojjSspwDC/Dbg9+k0Lf
dYuY0baNin5dTyXfI0xqBgzmMvQ0GuPB2+e3s63QxPeg0Sq/ppyNeoWYenB3
bjEWFsq3eeOfzDsoyt4XFWs07f76IGN9KyydLAABykR9iYfAy8FlKvp3a3qp
KkE/kbA8O6Uv50KsrSMv7kfh0EOF7H6n7ApkJ6dKU1VEFrWtgE+li0M6YtOH
YwargPqA8MSKG1xMn7Fnebca7nAwXZ864j/GlKOG+nC7nXti/Q+GzzL3JPNv
S47b2L4AtmvAFjJD2es+WF/8SRcKHLelkbVD5GgCThwnMhw11oiAFSNvo8oP
ihMY/eZ3kMUFQBzg6MGr+xxaOPcYcCyQIY6b8lowxDy5hq5pyQuvAC42tv9H
6wgSQ/ltKODUmnJg/5cBYlkgFeeOrOhM0SoZribY99c1DWT458JKOmpoMPYs
Qk4Orot2t9Sl/Kv18kghwbULBTds0l6FfZABEsdzqETKfWxYWpllGFMKkfZD
AKyAmbI7+2ndIV2Qjw/DzawjlhWPoW21oSDFlRdxMfdbTSZwmvg7bw4s+mAi
iMXB7O4GSyPGARwGjA4Zba7jLZB6E32/txqdd7Lbj+fKaQUmQO13EC7gDvPD
+w59QcLwOqCA3hPZ1SAh3SwYXw7EvgfABsz7XVhsEjeiZxx+e/9/DB0aJQRL
UEcygRADw0X0vY4eM2CMvigQEv0m281B4WU3xbItQDhZ4PSXGO5/TnKiEu2t
jpfun3TrfybERSd3Ki21kEjdEd2Xo7O1NErYtR/4gEO94ey36qPrMyk29T7E
Z8OPZ4QimBKX/XLucYXfi+MWhfcu/AprpnJslSWv4xwjmOXFwl1GKcqJOD0f
WReCF9ehO8la/F7cwi5Cyv3pD/oacSrABsC+N8r0tSVDANzmlykfLKD8G5bd
2XjpqskFA33Hur/oLiXBtpqF3j93IMMZMqLi3uWfkVK6FMMDzngXRCxtWhr0
QBfnEe3S0wMn/TC61lchyQR3mxVy6JNgjuaR613m9/i0DPsEWWHc7+lcG0A+
xpYGLh5oWQIbA6G37+rYObscVnfNGMJsrCgXX6acnhbIKzg4hYRZo1OEMl3h
+Hopgbyfl52a9wYKMN5o1quopzo7h1UwaiShdV+OsAykjwWNSJPmPCvAuCLU
d8TT2SGA2EFmK9yVNoSLF0LA1JzwsqlUgvPerSYy5HAIIAoawAjVIvfSqjHl
HyZbE74/z6I8r5Y8gowcVqfCivqw22ukkd/zkTCWB0hspjGVcqtkXnNfozTY
7JmgaBrXKUqshXqZUZpsy5gtG4Jm9j4RDiAmmyJFVpH6V4E7IwEFN66VfC63
oB8Yr1WZy7/xrG5PJAW5ZfTF86rh1mE6c08QhHx4cAMuHNsAVibpu6HgvzMs
ChFy9zmI+YiWBSCyGyz0qX/WU2fpPh6SglCBoT7OCN8F9fnBb0mqDGkR82jc
EMvYCNfZAHmBe830w1i+pcksHb8c0yfkzx6atoum/XwaV5CLC8iNuTaucaVJ
fJe1kIzUcxzYuvuMxK3LHU74Dwn/X6rtIIkwDbc5z1NsOBSOn0atbeZaHmSc
aMVYE7/saNSAnkSwE7a2yYH+C3kUvnoXnggeIm2U4H0hC+rLW61oQH1RXONZ
5vqPQXnYTvU0ayc7nzV3Qlh/P/zDmPdpc1HOCenyL0taAFPkLTL5Zk3L8tle
scjYhFejO54gOjoNuacw2VouBrzsnvMeLdzUlXb291uNqTBzH5WDUBcd1/WD
WM0E0bqiftxWROp/khFqNGMcF1CwXriA8gAZK2LWPtFanDPcYjnGGCXGgKLi
RT4U/gN6Hcc8/wMYry2CtpkHEdsHc+9pNy79SmUKjlIsMPes9Nq3Nk4Ezefx
FFD2Av9Krd3Ldvv1vHn0cnmTAzI//mm/Wa43NRUYwuRs8yvkEC6xrdrsMqsZ
jMkHiObhnmBtFxOUJ3YnR0mBXBsuyzxHSI/PmhFHqQYbxLfTuRaT0Dj5OnmX
adywa51kEednykZpSa6f5w41J6eIlQCGRQcSJ6I8QpTxP9fsBhDa3o8A4uGb
8dG+QAAnRvAuf85go0xyvc6mLfU2aAHnDnhgk/bUgPJrBcgsviHbIc8m44et
L6loTTJepHmQygIJQzoU7BCrVBYSokY9MdF/t1thKJaKjByvgbNjqjmFEnKR
HAmkgV5isjos2yviANooYCzi/dJSgpTnjPTAm8nt1YRRVis23zyelGeT1sCG
hd4diV1+KCioULR7Qlp9cdZJjy5OfN4PQBJZct6vmb0SOnKttGSGD8FkSIIO
MWDIsZ1af7ioiRl12Zs2C6/KDRIWfmnsKeUTUMrjJ6ZQKjdW4DvxI0ssq54I
x5qZxaUZ9b074zg2yoWmFi64ORA0WfyXBcY7OaKhdbsHly7WVyis3XDnhvPM
b18KMUTdTG3Of5aIYSqrVa1gvA4yQiTRF0jvrGwUSpE1ybvIiQQdZlYpNyDz
qSs8Y7WiIHytzSXaTIYGoA+VrBc7JHmGClC/ttFX4ZFzdS9Ayuh2ZenV/Utf
gof6MogYyEqKyJRB7TeQ4SHTsNfqsjE8orp/hz+xElnvJdDYgQx2NuqygpJz
/aX28/NEpiLYQ4T0J/Q0axoL6MjldKi5b8tlkojQmxcRZwZ/VlKuUeIu08AB
Hyv5PtadepUYv/hpNRRznRSC99bemSw/Q/hIEC4S2cmvR3KFn3mr3v1KeZZC
BOKRZeVsDYSm2W4W66LmeewHzs6KLvOuQIOwoErQK1pojzrxFVuIkLw8NDuE
FeMNK880mkRObl61Lw8kZUnxNx3nIQqECs1wsuwRkyC0LMhHbS9E8VeYn9Zb
HBlpAsG7CvmBRfezxC8MJD79scp23g0oqYC82DmfPVSrQwrZnc41BkIUcpew
+Vpgb0qkREE8OFWg+sCByTMlmNLk9IeL9GByMXKP/QNWiuosBm+o+8BgtZZ8
EHL/vX3q9i5UDnpkRh8uYo13+/SfdZRCFqSIwdqwqvfphjtROC7syEKVftso
QLg/nnL8k5ph1nkj+MREtK2JvMznDD3pGYOA3bZM1Xf0L3SAdh/YlX98G9Sr
u9vq8WMYqNwcB8TcIHR3qZAFv1NHrLisYE+LSkIa8Gd18ejLeyYxShVxBKLP
MhDWVXOkw0JyC/+uOz2aWoiZukWvC3hsvCB022pI1FuTcAJrrDkzXeMtoY/Z
VQXvRaTjBgX+Fb7bW3GCpjzPgiWYIvcAT45oKM7Ms6Ksv4iF2JINJ0rAEpRO
lxNyoLTkARAbcfEWNwHqlAN1O7eYcyPBhoQHBdTYeGjohj2NzXwMc8v5KaEn
Sjoj832tvvgsfq8kRBKkZ5xcmPUg/4hTcVglyomJ+x9GoD2XsA617mCfho5m
+B6N7xwE5NBIXPz5RC/vIUBYaAl1FgH9bHcMbT7WLMopc5CEsfosIpfsO6AF
96x+xBgnduEyA0utDyGI9MgibGdDaxXT/RTDwA7l8Fa7Wu/38tU2mptiKe30
UIqNxY53q66GlLNAXeyh0Wyp03hsk9mCmeHpzEMxgtdHZ+L4c8C2/qUoE/zO
VE1Isn5+TVovXB36i/IJn5WRHQ107xN0HqXnkfjYl5A+IP1kaQ+zLk76v08J
c7lHOP5ihZ7Dg/cJdGV1pmEsXOfKUuvlQt2EQHowHQGyMw8XFfAX5O6FU/oo
8gdaq9XMMfVQ0QAQ7RaG+iSAHFy3YTQJHVfRq2V1zLKNyrWY85OCmsD3wloP
Ac6SnmzlnowvE1F9jTjaVFnJdsBgjZ7KnahZQ1TvFfj/rDuFjid37qiGwgz3
OcDzea0DwZhgw6vuKemOoDyS2ADGfeBBu0GlqrzD8PE3F+PWMraMg2I6tA2b
kaskvpXNpafBG9t/uIAJsNCDaoOGuq+IdMdHxobjh8zboEN0YwS59/nezJlo
BIpt1VF3pfNrdlbHucoMAqfslGeUremGIOXgUFN8TyN+NS/zCG1d4Rz6fRPt
qfByBr2dxeLq8tOa0MhAALz8tK1uWiAqs4lvC4xv80JseqsNNurGdOhZ52jH
HzgeUmTFitHLBfEXDRad4YSXWgahMJgOGwdL09eVs9FQXMGSDRjj72I6CCsH
NZmla0C3yUfY3lUeFwd9KoARHif5b1ZbVJS3cQrX63j3P1a2IJJO9iZHjuiG
E5g6Ai03GFMDSvOpqPRYkPChwZ1pi8mZuIKB+FNBA5W2WHM5c8XTMtowvAcm
grHhQYkGiQXdpoKXBFrskie0uHeYyIUfmMsKxy2xfCQDtteuP0IW6k7ouI1P
nE1qeRtFQXHPC4JfG6eQdE6Y0W/ivQNQd2J02wKyCT4SrUXgympBS+9QAev3
SCfV78U3zi5mdjO+PCk8MkPSB83pYRR+/vtOtDTXJVi8snVdA7Elq+CcreTg
NnTUPbNLt1l1i0ubI3XzjC5Ez2ghk7NPT5/fu8v760YfgSM11k+zJm08xiWS
SqGvWVAczLOruoavTcR9//vVWzZ4VgOo1XnotXLqP6jBJhcbF4VIaljLVxpX
Kr7+sZ6K/Vz3hA/IVRLa1LWTsGEgzAFKX23rJYwyYv5QYl03/Pg0IEPDbzjr
lVR8d042z/vUlmP9xfwJvVzItbEbBk8DEfI6WGpus8G3EHpDTs429Bc+zrPS
F/p9lmZVdOovttZvLCTQx3VENU9d8K2XL2FAWU9JM4JjtExAXhgGSK3tsXBU
JDZZ5bme1v0y2G5TTxWYcsy0KJBVjL/tIBP4Herr1Asuk9dpEsqPi1xLYKt2
4ZLhAqTW5qzqgojZk8Y+tnPeNSlobdfDTWZyQQ1kGX4+oofj/n1la9XjZdjB
+skSlZ1+EFedGATQNaAdXU++CEaPkm8rm4fTyZXiXbren+BUphOlVh+KpjkH
IupQ0LaV70hy8ztVd1nOznc4ZzNSPHFAFSmiIm9vNNndKz87+JqiQZezCRap
FUWaPoqRfVLR1vzg1IgQLlw+WpaZ24FYnWleJIqjo7PL+BqQZL1MaRSMSCHB
d1qDaDACRxZICN3EFDid5xKSl3uoLKygw7asT1MiA8Qjr4UGEacacyfQM62R
EyRUP6a+fkViVRZlgoVaWA073eXCiRk3q4N/6p8JJe7Xl6k3v1Y0iS+U6orP
aIVD9aw+AUHTQrw5qVkEZBly/N5T9qMb1VTPkOZHGQ7fFDhVIehvmhw52V9/
KSBgqDGCWKj5NGLujtma0Dij9LauWlMwZsJq2KXacgOC9dJissrMrAafb9zK
cVYMfvwGQ0UAN0WlcLrjxt4G2PkjIdliF4jWPPUjFHb2e3t2IcOKzEvRyblI
qCbyzevKpgsAK+uHBBFUp78jN6/uO5r7W/TP4WjK/NFSj0FeUxang5a7Vrbq
VKXNdMo/mtgxebu8Sv4YCDC5PF0uiT2pn2C3GvObrBi1h4vVPz3owOKLjo6R
CGT0JC1ba1i8BHSiJmlkDzQkz8pNisxGGuHVnE7RefHa/FW2s3zgToNC5w1G
WcQlmfYGyxqLv84mWzs/jfuzo7h8P0k58lo4yuFrRkP3g2XDkfQywTsuFzSZ
31FCNVUEEw0bLtms80ksQDyz+BiqwEpYwvdtSiuWZJD1MedvXQYMsRs074Xc
3L+QJSDASHGB+rh6suAGU6d2Pi9rOQ35HzsHwOgjZYnELi2mSLw2HUfNmiy+
znNxW5YJvT9CQtqN/ZJTpb2hr0z4IlGj1AfbBaL15CIxqkFH6IfJe0hMW+Jc
x5aOi/dCnwy7lSpOUSv0nqIWLRa3OPuIzfSKKe8gSKe1MBeHgh8xCIaXm7VH
KPLMAFVUPO6/lr1yIc5lQcVBjU+PJ/7WTcPnr8a4GwRftJxd/EIletisimXJ
aTYXaSOVPPUFMfMdvNJecp2buY/89UqiQlE/VKdg2/X360c0VsfiCBez3f3h
Q/weBfe++ZXfzLSi8EaWYRyHFUzxMo5/LT6eMsOHjxTJD3/k10+19rV0+Pv3
/icG6IKV509CypDMWhDaNkogXkA/zUdykn3NJCzstnwj8MHli4hH3nuWCyyU
NQz2WZIV7azkjeGF8xe9/Sws9mEQjSfOPeRYXvPdyXO5ZPvskzqdHUn+8kJl
ZtkE46va/mcRsdVNTT7LK6uOSAtwDfj8vlvd1wAII2bS94GU41uQIy8C6T01
W6+/CaYEy1NThGEhVlwcOsefsgiHMdbJuI0EIUI9hEutc7nUBn45sggeY2r2
UMZFF3gQXSBe9L66v1LDK5PTQFtwwJM5B6QR2pA5/MOfnbnIKEEafl+kD5VK
T4432eD0bFniKs8ir1jYHuFIXnOo/yeNhCzrnNP31AOeE9zzLrQCmwCoH7LT
1SsSQudaMXSKT6Iu8Z9sMrp0FBYLvqRVJ8RFGjf9dl2fykoLXjY+3VcHYRpE
FZqbctxGbi6Zv6Kn1G+LrKAOlactyNaSabEv21TD6EoA6IbyNC6Y4pmnNctA
/C9hdPrK3+YLjp7wY83mc3mvG/E2a0AUKAzO1GvPmmi5StAyAtI/pD6fNAjx
7kd1gHNwI4JW+NmdHURU3lgnhdQRD1Km/WAaBrq2oxcZ3JMEA1eTu6dwKTzE
y/YN3x8JKVbWakD+Cgs6aoWiQ7ByhN31ZDt9JsZ8crR0mVd6TkXypnBntiij
DIUUmxWi5wk61ozoKqht0Wlob9KhHz7euP3OOpZpAlHDGz1XM92lX0+wQV9h
hDaQC2Jd4CjT+V3v6EODSIAFr/9AZRm92EBMgTPQm7QlZcqiYXfCkwu4QIR7
+NwAcUpw53pmo7wjSprA/Ki2hmwBmGAyy1IFxzgQhU0vo7YldkiWZGbRJdtE
pwao2qU7YmN6HV/qXbJWRvMADUHRxSu61IVxdh8J8RFCMhxmU4Mqc2G6DKU2
Rn6oLRouKzm2kRYtoG6FJop34caaGiFmmrd6qSRoWGK8dneo7MDr1wvJinM2
9jwr5K0qL2oKYS933CEts8fG2eHuv4ETgrJUuQeL/PXyqlKrQvSeE5JXzO7o
XVGr8TYM9XGReBk7e42W4vyylxE+Nx632fc0gtT2e3qWc4K6BuBcHr89EXYv
uGZ3h/QK4FGY4kCjr+icATSUGKyagDc+viUqOgcFEapj0IwQcLaSAGACkam9
ZhlRho1b8+gpA6cwCJ7jZvNtInId0TIvrHUvRQuoQXd6kohfppoT1XtA12EV
Dv5ZLNLEAkd2zoPBwgumqYGlWJjKRFvkzbj/gSoEmPHfq44OahbetVfBI/kH
POeoti+hdR+mbg7cMYHnWPddsu8lRqeBp014THtinRLdDTqld8eHJFbqbq3V
uZSbpet3aWGZh28GjErptcgLOc9ipZqwjY56LRioSJBINEOxy7/4wSHoRqGJ
8RSG5Ybg+Pz7JkXkRFtbZH9UXz5MjrhWTGMgWXVrLuOIriCS14pbcsDFI7sq
tPvcch71j2HWJlJixXHWXKFMnMJZkMc7FtvVOFmlxpTiSKdG8VUsU918nIYl
7afFgNVUMUgJIMmEOq7qf8RTXCQMvlacigxUNfEUmq5rfPNZ69ee4k/fi/gq
HLA0/i/Phk+LI4TpMCBzi/gqyJaXj9OZcaATJ7pYZh6EKBwvi97dA3TIjxeq
sAS0sLrDHUr70YunhfIAfPsKhGWR6mgnr6DaEAWOYWjdTKUyf+8LoqkKQR1B
MjIIi7JXoVoAGckhP4T7mW5cOjiwdsnBvXcMRu4obXaZPCrUnVMFLOADLnFu
z5dZQrJtHfZAplmBs2VfaWs9CsfGp8auadUqJw/fDwxlHCiabAIEurjm9QCZ
IMGrMst9VwdVZsapL9QLDbqpPSPnE/eCa9OIvkZd48M3ZPWLNFTZeCMlxBAp
txPizHELsM9ZQNib+ZgkVmkik7NhK7WmnURDbK8CeEchMaOht5lVckKasbhg
DfqJ0s/EcKFhUj7dD+PlUjpbT9rWjpe2Egx8lWZ1ypT2KKrSmpR6JWs1Ujcx
prm6NRd2ubBsiONAgl0/WvAzBsRvXcDR0boYRUunr/yPs+TllEnyhMrcg0dS
zubXtJ79aWX9jbEX/1W95X6wR3MpYCLIreQrndez9E/bvG/BVNd6tF+krBZZ
nLyxRajigOH4xtTHpt59NCtsV77xqnLqgt36qUgI3OCujl4o6NAKcc8Om0i4
iY7E8PYwqXNqJGd8EmZ5LN5l3NwvfCwGsHcCqyNV7r2LCGYHr2v1ukyVuv9Z
6eX8imHtfMiZJsmORUaw391psfRZ+dBwTdjSaXd0lMir1k6DDtVGi/kpVFi6
nZUaKkHJQnK67d7EPojrb5nwDybkuW8z5S3HCimAijBoPIzFfxf7DiJa8xGy
GVVo8B3X4lYwcX1GIJodtYrVOR1dYddj4CPUO7bSpi3+ZV66SiKXEisdIenl
YSKisgpl2Kj4D2meAzqXcmqqhxkmDmKo+qjvL3s3NQZ+6L/6XjM5Ic7c4G7G
yxK2XbvClZmfvVVNiObnIQVcI8ytU1JKRx9NrABmEvOcl20e9/WgUnaikBfz
uHUVTAQF780LcBbbKbmsyPfCkXpVz2jyDhVyVXFezNYy9YvRQIWu6PL4CCmC
0Ca8/hKDQ3l+gJ/QGGtxUNU3v3mQwAw0jMPrXcLuXmlcroQ2MDeD4YO8SF+b
caLP54lEbCLpmgbW3YmZlDZS0VtkEgcj3Tytfcgdj8t3hL6HtKmPx9e625Ou
pO3vcKAG8mUtofxbDcNoCk7EvCEf4e0tUC6g9Qjc5aZW/cTi7yW0spCymVL4
QTTWH6+Ev7MBqbR/CoCl2M14kBZ3AzCL8BPla0jX415UAJq8CoOGCWUP+jaO
3XS+jNUtzyuwJi9Yl9lj6Ae32xQ4tIK0mCsh8VqnWczBiU2csl414RSFYVHi
dgQSqtB05BiQGe2ywX4a2/hBHiz6WLCTC+6Ov4GpSOu7UqYV97SWJmvlMrsI
rqunwdGWthwUI0gdGJCxqJ8kJidfuFItw7XMsYAxWMP0QwartUzZDEPzQ+CI
MjtRMJdRUPi30EcGAnQQ4ffQi+sY8homU/E9kWy/kpoOF0f06xwGuzPhZEAe
uQI7Pxt/N0NBvhKTC3gv261re/sxI2zeQv3OcpAIMjqXw8E8auCJxw2UQzVt
6iG3cfYVBJLa7URrgAGk0WM0vt2OrPpr8BBqI8TgAWeayf3WZ+hAQvmpdcVF
jtml+GEltq4kNcvFbpJFdGh1m4f26tqmQmLq2f5+4CzNZZSKBbsnrvinRP+1
JrFbzsy/wMhLfi5ohefxHkKMbolvcboHhuGX+PJE6nSVdUff8WeeF/xn8NWu
R9YApEqx/9Q4l4sl2zPRHgTLUkweaEVNM2jS8O5/N0UuTyONiEQ154PpmnrY
1pR47vfJ2Porz/qss/P5FJH1iBR0JQe1Wkc/WX+b8HCLcSvX/pQm8F61Gh7I
IwqS7jFhW9wKLM0S7A6XhSFhGPS73e0jsU7+4+cFvtipVyhK9PC585rzs6RG
lok1n49Md3SghC/POpfzRa2gxLEsiLjNAh9+k+yacS+8TgZZ5q7zgOXrLKnm
0H+U0UNz5oS8g93nrSAmv4iztrfi+5DcatiaplPzpkAegd6EbEJNyXT81KZJ
2qm+aamDWzouLn34lz24cCIk0y7ULm/Ev+r2L4m2f3vyLIWi6E/VvMAy4A5o
40GpwWYDXFgEsKa5U07tsF3nZzyf972BdcF758uHaH5RI8kwcT7gMqad7U5k
xkjyT4YLQvRj8drppYbUe6CTYcrLHq0D65/3rd5HElbJsNBqdU+ELhHlgj8V
qO0IHsn5NayYRa24DGpaMfWaaBTAxkyTEeaC/KUHjgCksdGmhKsLUQLOhhjx
vjm70XZg9RK7m7Kk2SBWHujhyCcWLOZj6JZujyA4E94blA+SEhs5AjLBe44V
7wtWKU86U0UkvvRk5g6hC1Tudc9L2Tgv6d5sW/16jffQ/Mhyti40k75m7r88
izTdwD3jQv4kAcftIW3kF/tjqzkIe0HllgB5l/rNgDIBCqfOSijUWuqSL8FL
SfoRYonIemdVkNRTBUsTaU3QS8SNvHQCHPJ10zuMosRwo8QPjNl9hkqjz/5O
5R+6AAo58r7M47ybxyuXjqPaZ8LQLDueBLfXRfPsr7GcZUL3NSyeJUCPKlrB
ab2t8NV7hj1sGq8nNB08gf0Bn7E/9t9Nru+ZqR5ZKu/00kGDKP3HoDiHaXTZ
BFpvQMB3c+q/GoIJgFLP26TyyEzw/BR4H0DH/GjBduN9tN6hdgztD0i+54Ka
d0CP1nB+l8uyLiii0pvUY+3dQQkBYw6elEUz5dfiNInP18k4oO7rslRNm9uY
Ompa/s3PWe5Rr0z/01+DulYjHGIotVX4kv3LLbitnPFy/dL0j1H43DrOH8FA
Yow35dlaI6L9H1qyY82GWLTGFGlcZHiJbfo2klzlpWgeTHgfgGb91ZUVUK5A
lNGpc3zh74vJ5B2taQPO29a826jJG2q7wEK8K/Tk7BbftwG263ocajh6Z1Yv
qyS6lvMuLpeOrn/b/nPe0ToMWH6NuVOCUnYWuIOniPB4a5O4iUy0/MN7ZRLh
yWWGrTMf8GaOm+47eC5/wCtVPQt2bUA7Q4Swk32q/dKr/FHw6yjj/GVYUU44
HTQiwu3QzYFmFNBthvjULh814lzk/YVyyOILWVmBsSNUKe6+iCoMQw7cDz3/
ySNT7Jvf5jOs91AE1GRnFeC13p9PF5YBt29QBiNaBfm1pijISg6cz9zqiMHk
L5bp1Ykcu3q/qFXsej3R/llZWpuW9VVne2uJnmHVCnqG7We7joXBdC2JpAB1
q/UvG0L6xwV3xjliJU3pnPhBStZ7WZWUHpitU9hFsFDOgsK3Pj78B2xWPaJ0
0nZGulm9FpUgw6JsOdIv4mQtOZOTX5nKXAPW4+GoCrS0n3BUfnDDFqla2uHG
0CEkp5K8nNyyebDvtioz3QK4skW8d1XT9j8GnshHZw+xfb0J0QPAcJzqW8T4
FAZrQ4GV4rfw0F4dxOaNNZasqHZwd6eThuYnO1qr0y12Y7OpuAfAXFYhNPK6
TIAgotNyCYiCqoeXVNe4564QocOPCp1PmDJ8HGL5ieaYMCpCJQ9ejaa9ZAAr
Mbh/5ZsE9feEeGeCPJH6Gk7EFXlfjONRqF12f6VlmDpJHASp347/nk8HjvjY
IFZnF314OFE0FvUUC2jlMWB+kR98qE2RN7ANGIMGNTkEyryBtwLPBz9OnNsv
uz1Vf2lyl+jOczKYBaOGLaBY89fqNHYYgjZ+JvR1wOplL3BwmK9oA/qrP6BS
53aZagTPsvxJ1FRmU4pEbEi1GSXA3gW84Ebl9kQA6J1OlM5Hu56gO4Xb0L+c
FfIsmr2AYyr7VRguNMHeL6YaITHFNKrng+KtQUz+3DgWJobzfMrCUNF3+t7n
dddLC/NkIeErszoEz1P7MykWhYQlNbQTZxzuh+1Jkn+HSNVFMNRk94Wx+L/g
+fY6Rm9ZFRA/cD2exYaCAhVjcIx71L5F9vRJVS0IagiSRTM1QLtV2Q8tSrul
+3hUee1073SHNtVgiUlXiD1yt21t1QIuGXhU0WD4N+g30yvlAq5FMsqK1qxl
pAVRZTqDrjFKt66enVBT+v3pleBV6YtJ7x2QYJqLyDVhYYqQCFrBPNF84/fi
PFLaXuUOV4UV/j0DtO2ZstHRoMpo/3KlDAR3lskI2Skwr7ley/kenCX2Ts9H
+i/22oyqhPzHfQVnQKagK0Jk/UMeOHW/Okt+shvC0MONrjdQ+BnhbBMc2jOu
KiOhP2j8sgQnEhUsWiiyGQrlJlRrAYzvYgoewUcG3DP3pEcqWhzVJRhhuyCq
qAgFryMEvtON17aYB0oK2YAo5FlwT8OieGE/3BVGrFBaxhnto0uZ52V+cVEh
dlfM9WylOR65dFSD+awPaWsH0qtlSsenL7U1qC2yGHSe+nQ/gss62tfj5zlI
VmTTKNyuyyeQ8HsbEZ90VDXsAJ2sXsF0jWo8jIQshE2sHkvJG5gx2k8Vd2kH
/SSFV8losk5wlyvUYuW1Jbre6x/T0JExhGUNOZ9tb7V5vfalzGoMwGSoCf2M
fZmSg/FF6epkdzOrV3JHVAH8FJGgCBhx97wVJ/uyDB9r0gbSAR/gXPiBzplo
J/Of7j8QdRHQGqVuEOGL5H+XP1StQnGSf4PiQAREA9EiDjxscKaHCptGa/P8
laTXNvihiZk5E3MTvPE+dFnU0FI7bZqc/UqWP4UbXPsqAv/Kj8boHdlUuplL
pVkvQCj4g022a6SJP+dAsnSHs4PH0nl8RjsYHNJlCmV8olA7FzsHoQ/37j9h
2Z8ORbJCJx9whYGAUTAyPwz2IhaSGDapynv8RnFkIJZqpamQOoKbDH+lMDcx
uJYO5z04EHlX+58MJBAMZt9NsnWdMhbQaWGQHgjwRIu0WWKIs1cFlMdwbhaM
qA2d/bry4IMitpL0YGQXQew12paJz0vPcbDaKx4vxhdmBi2yocXABZ1Q7Vsb
T22lkfw5Ryo66h4dQKKr2tDmko63itFYOrn/hU5/DOqz5o6kDzplUFtzb8SU
IzGbmZoh5ig5521urOxKxLH+PE6JHj/chlnrd3mAVrpbaE639M3xbY/vlHm0
fvBgQ+KLCm2at4MzK6bbUN5zprtlEUQNEmVnYPIyI8ZCKC4BLHmCgUeNz08d
fE1q+iw56RUZC1FomOtBIb5DZDv5hSW/kxY4b3hss/5pqdF3pAOgoEpLeENE
PnkSLPXQL12AHFa4VHSjz2akHXMYHie/JjNM8W7MlQcXjpTa6T2e4oAovPCv
Hb/HITaNk5ZdNDhyBwleNVEXlireDNCvKGF5Cc2jzf0p/kdNteixcUEiHNwz
zKX3x7AtIjEAOgLa1GutdVVkO1dUcar3zPHjEApFTF4UzUA5shmuutbDJPY6
vVpCRHZR20ElA1jhkfRYawPZl/K5xJ5mMs0+1lqQaP/rqVjNzz2etj0y3UJ8
jkhdagcqOtTHSAktZV26VSOK4oIVsjcjGkhKWmL80Vm/qLvgLCKXVOqgm2Mg
wfsKu9s9woU6O8WmQfGLJCkjG3ufOkVMQ/Vaw0dQhcVreLBhL+6r2vllSXT+
bCqFx6jlJ29VSxqXx840pRI7WfYtTGg8lheqm17go3/r2Y23GwSBPPR982F0
c0P1mxFIii7MU9D3E7SPRsfNCmTZ7Joct3DDfgyllH8j7PW0UTQoxOkEYej5
jts/o6H2Mtv6PRIjZk5tVPvhFmQ/RShO0ZRkwE/kCW5tPjBDvsASZftjoWh0
vqA7d/poK+i6cI8Ul16rGKcB4XQLs7hNTdrHxKYZBjhP9AkhpnF5D6lTMIJE
k+S6r4mb9jv1G/zwsp43Yd4er34e8cLefzSQHLVwDYmAC8jsjSegeZP7C3Of
t3daoMIX8cZ9UOckPiPy9trCRZ0utuLMgWXxotW1eA/zbgy7ptDpb/6Fbh1O
tllzKeaX9caddfU/YE0ctF+EY9iEyMzMA3mK53/uzOMGV2SlIWeBNNGN4LcH
i2DLzvM9ChtMHp/Eq8M7nt2oR0hy6EcfzcUCtLh7bR04fn1ADHQlqO6gmC7P
8xisOR0auHSJ919PmHwo0jucI9poiWqq5Inf7SOFPETP/qB6NmHGmRFNjFV2
Z0J7wNXv+DpPDhQvlhfLXzNoeoru7u4n5Br7TiEwBv5nuZs5Ce7aoA53v+Jy
5rIdpHrC1KsSyULvnC1szmvi6QS4CIs0nj3slGw7nhu1h7ECbYEMCKTM40q+
ffOI0dUR14F4jbXtVJQ/NtfGj7gYnO4eWHmWIWEvIZCAl7PxapsRXhE1eOM9
sPwuTMPAttLcT6NxLROv1bWv9+Wkz9VZ3543VpDnvL1g2NjbvQIbwUz12Ldp
0k+88MIt35Yo6hp7QA7EX1cypSbg5AnBD6M9Fv43Z+6gDcF1vVC3p2+iro1D
Uzood1mf9jW+IZZQWLDSo/ziY/GVJZ2qDAPrI1Sf7sMtomaa6Ds+IPs1RksK
xEvnhQZxoFzpkuJ/CY0ZBVjS14s3GnhN7rDkk4ISto9k95dOEbpQuBggR3iF
kmumCfCXOIi8IPakYRLVZs5FuFjtKakXr9BODvGlkRiWcBBWH3xl+Rx0ruRQ
Y4Zz8OQwVxyuGgzqH7/QE86GVJLSMKBo5Ph+RNHt8wZtt7j50hBNLtaAGQaW
Ceooj3GKIOcjUyl64JolVXcxNbL6B9Qp+148kTTipwlvYN6moChJ76BEaVXv
t3OrUFjiPgIjifrSW7FehGKdRDWfsd9KrARPbpKd7d3OTXakj/fdJr54QWIy
fl8cz2TzRxwtyy3daOJV5ZOdEEwB2ZM5RUZVuN6t/NbINhwlcHMRC8KXxW4E
kZHWJ1RlTWmUqGduhndlyVEh//nyNwBx+3pToEbrSrvIEEEyId1wgiXx+hkG
+B9dHrCMFI7zgzhbFJyCjO9YWV6p60yv1dBB83OAQ01VC8LX6Mc6bWKg+jpQ
Ov5raRfEPojiRRQCCqpWJH/TvSsoFQtNE5UX6VL3W4Ibs+hvbPuqhrmL12t0
mBpnHuqm3ItYad0xbiqjWyDWndtGfAgMVWA7NtjxoVGiaAG1Ni5SRoG8BgD5
SfulBdjj/TjtTXrIf6PjpXNKJAt3T2AoCOtI8+R2wf8c0e25N8fjRcsR0TQn
RbMC6pwdA0DVst0UNZ0tTxlaQchq53b30g8w0DcJZ9ZuKbrqK2wQb/ioYamw
o7B9pzYYgqkSeI4YTmTDfcYvvBj2ymClPWyW1MxdcvAGiIkuzR/TuWqjPdhJ
E7MP0u8bTXo56CUKeboi7dD1nwVpu2TDZlbfZg+Yf8aASORYRlB7d/+Rn7KK
0SBSsu99gxsmTmZS2IKAS+FznTeCDx2eUdD8LdWm8X8WN7AYjmneFQwxM7w1
SzwdJ8YxrtVvt9fuFmhJ67j+i+anKBuDvFB7cOwVzkmjHSxHfdU4sGuI4leN
UhwgDIqB7sTwGRGJB63HZjV4na91wkTLkL10ZBsTRRk1dLkyiIjsPXy8WnpF
E7dMIBKdVKfJIyGf1q8ZRiZ6n2rZ7ckBZWoJZBNF8/EeZaQih+/QxsAE0SKb
7HwmyLmhuY+dBPaJh02rnjiH55LHp6U2T+HdLbcsOBJocKoU37LXwM94QuOt
YxUxP+RfJmrcX3rF2+LD1TUTnFxRpkEy6wev+GtGcFbPaCNi9tr2VP3f+Pp3
P6eGy2tqwxZvrMU+NmEY0wTLonI5cmLu4lcgX/mBilsEdEmTTE+Ogl/krkfk
ArnA6gimlH2KUvZsps9ClVCBbFh8jJEjDUlFgeOdbajp+MlXi76SG+H0rj4c
4laaemgN9GpavvIMnfeWMhh5RWboQAtjbam3Noo088Q9ddfsZMXh3paxBOlD
19VNfRrlV7XvvdZQAk9cSsa6r+zPO0UCfxL23+Gsb/lYgci/8su/7smxyPUl
qiy2yUg1pPQEtp//7MtHVp0hXXKMY/ptZAxa3kdC9GwNCO+ASwxgdN6jMwie
9Q8j1vLsdknCJSYvIF9ar2VICXnSzwmffWleIlcVywYqkG7s12oy0rI2gY6u
ybyJADu3TPErdB05ijAfL0xy+ySCg76TREb18tQgmM2/za1lf80box1e2gBm
ee+e3w1ELRu4igZDqsBsoZda+qzFGdzcc2hl/7cx2VZtK1EhLhJ4Jq9Bu15I
+KeANae8yj148pSZSaKPimEWEdDp10RT5x9co7naZShCavB+kqa9sONrW8ZF
zY4K9BGDAYyfIA3pp306KPL2fJD7gAnoV82cnt8JphFnhR/5MZqmBQmv2yPt
pJNw1Dvc5oMd68jdl6Q/UMdgHg0UcOQfn3+L+iJE2fHC4xzxQlSjOO/SmbHF
EJd9YDDkQ9WKnZg5EePuKUHo9PTlQrWwc5HUysnVeYCs299hT8j/Fz5MOBr9
2HWCX+QNv8aWf+8s6k5QWDFJxcuOq+eM9i202IISIyg0AL1OQpmDZ4QK8cuZ
hqnRei16zertOUcJ6PNWajoShM4z+WX52EuYRzcCEtaRnlNkHkHDFNJyxup1
afRluVjDZKMPDOu2YGfjhXHZ/mmbatnkT7e2MqWdGIr3BCww3vxMxDdKAHmH
dq37JLqyBkYqePbNsFUN6dJEahDQpVvun4xFNljCWIYYqVzV7hFbZNAyZQZe
6PvNLrw46E+unw1EgDzhHEYrCYASyY/WX2YO2sorlEZBZWMQhsszjfluWY6q
Def0xnwwhoJagQlOicaZGI+U4CY1WTqK87RBkpus0sYa1N8IcYCT9YFI02UV
nFcjXA+Qorjmpy9T2/UUFXRtxaPyu85eTLaW+US2qZUjoRRsOiiWcyQMZz+H
18OjCXSpui0R30HnJg0EJct3dpsPBUxVWozKWVj+ofxsPBYdtGeBQOfeNiQe
ZZAtO/tjwP5mv93wEowK/rCteKbBYK789Htpz+ao44KOz1DsYwcf7s/SdfEk
d44VmVKv469ZnFKUszDcmJ1kHP2mjic/nUUxZTvTbHpGc7Us79i3DgvE6Fam
cfmks+ySP71rAQNc/36BGx/ITa5O1qCqpWgm++nbIjXochQKQaM6gzwkS6qR
P36EduhE1jFqWbKOnRZh3vIoXcn7V2nxX9LgqKvjum8gv243EtScxRbBJeWY
8qpFCAe+PGbJXWqALrkv9be/psPhDiv0ZNPpKlQ12I7mIM1L6uZZ3BtXQAXH
BX649cijdP8Jwgi/Nuj+3hMcZrGjujCefbGFVSDYFDk0MNwU6OBN60rATbYK
RN57CXz8YC3z597QvB1jI8Aygch7TsYbEV7HKJB4WAIZr+L/R0wzbORXsvfZ
RQjFeQydZhcte8XgUZcCwmv9hRMD92K3QC3BtyqiLi8lojKzMOOdikRkLCmR
1afdp896bRxKlysj+I8x9PKNnd2rHT7SzeMBywul6RsgqUOzlF8JwTF36Uop
1rcEBv86gKciyc6jTZymp1I9A/AW3uxD8WwqzHZ2ox+1VmbkXuzbpu19tUQz
40LdvOBubGyTTH0Q1yQXcdi2ul/m+zSJVAz1l+UzZAar/7BL+xXQ799LPABS
3IHHQGLqJ3M4lXPMZz+XtISf6wtD/hgVWIDQFx9/svJAV1MK8oUKDbWtWEBQ
lj98K+wqLJxa6XZ3wmipMTz2Zps2k2JsEQylDCG0z5vv6RbzzZifAQdoQ4sH
uqGKFKNI+sHG8+kIKUbeIr3GuKdCuHfYeimwkNepuVCwM1f4/gfd/L51PD4F
jxHX/A7+RVJCrZPzN5wIbrVlBzEQ6OJsB6QAZ3GyYIrHIwiJLILcJo+5Ne5Z
ZBCRXLh2piKVd6RmEepmcjZDzOU2b/ebFMjWCOVJrZCCPrleWXV300CCWr6q
Ycm7LvY+Az+KRu+oEqgv1DlK3gjP6+UrSU6syIX4E/tB3OwQUPpcO7wK5Van
cKpKKGWD4wc+N5fOQT5bh4AKqOU22bq46FTMZHqR+acXnICk0eT6G8rp/ojz
GkAFSBVXKGnQmh3rKImTh2GkpE8cYUxdo3Syg7oNqWC83jdjY2mi700GWiUU
9cgMsG8oEe75/9WGdtArw8WJblwSAZu5w47rlbM34PPTvLjKmsgQY1xSpHaj
nFb8/VXH5osfTD6UNCkZ+ekB8ZzCOmf7MFva3tDXJHiTqaAkr7jTaMsMediz
f7Gk82F6yEKI4O7/eDaTE/kSF6gZ+u0L4HUkdgOFs/3ZpgcEvTqIBGWWYpfI
/QX1uMgcKG+d8KlXbZxjG5IFLU95NZLgqH5KSx/ixvQpNbFc54ovNaoZMQXr
2IwXuQ29nggzg3A3n196vLKbbIBBzDmXeVxNJRdQRiFeUo/na04F8WxAWcs4
QZs0AIRUv66l9sXrKzb54j0T8qpWys9fCOXLdRq0/o+E2zxrQDRzstH/uo0Y
1Wbc/mP8kxnJazqWLfK08TQceGAVIEOj2Yp61iiHo+NzqoYO+SlS239k72wA
tR4ae0MeZrKy3mjWQbM4m9G4TYsw+rwoPYVzNl00hEVsGf7ke4MIQSdaAsv7
7G3cRlpmcvJef4vwWa34GOU04ZKkXDoa0jvfgTghfDV3cmfJlgb0Iw2pjb6y
Uj0bMVq380USPYuN1Wav0/4LycLz2GhXJqfdpb9MTk1y+L2yfKn1VRRe7vQK
F1QAdZsKFe76Fldy7c9/VSSmgSYzM6cyQny/r2uyDZoMdFGbJG3XNVVPYa4n
cVgpr1RP8aNs/r3D7qCcL2L1QrHXPjhvcKeBWkMuy/3xN48C/folN/0raj9V
mxcUZIsE8fruhQ9ZslgeeR/q9OyP+ti9A0u5qg1njbqYk26ihuiFBIFBKFRA
nTlGG7ymujBa6HkNOmlD10hDH58fDrwo/7TYwCK8swrJ4QYhHaopQHl8Fv8/
xjBG0Iyxtsva0vXTLBSBozLEl9fclz3KuYnzW+r0UPDRbzzpNpyk0WvRSjAF
Mj/wXdozcQCSnBUlW8lfvVCwE8q4xhC8yhO1/JgccwU6bZ7CgsAtp2O4syUc
U3BT9UGOIJzvaLS1Z7L6oRwWZRoXEgivSUVeAwiKF1ThFSVhw2FSEHLLzKOb
dnwCiXfJ6GqZfyN50i5/LuZALxHHL8kHWsCvxwUBzcHI99dPx0JCIBur5Huc
Xbyf/vGkRcbCr2+oqAKd+dae+Yd2an/lNWm0U7tuPf2vGB6yqdi0a03k3c5t
zvC4Wowmolgi9XGqL557pV85oLawWqs/A9IzUZpcCVFomyjTlnI2E/5k2B1F
Sfo6Ke+s76z1+wOnKG0Il2Zfa/36tFTdJ6s3Zyp4P6me3Dm7xn47ijuq2Z6x
DVS9k75vfXejob/8dpGMJnqCoFYzDL5bmbLSvrLS2nzcNuertBIUqST7WLls
0LF13hmY77d8ZTei5u9H7ssc/D+adXNp7wDdzB+SD94TaM/yQgaYnGhAYQpa
m8ptWabSYmxCxyBIw0p0VvjtMOMyiZCfUJhVnVyvX2/3zeTABWSKcVGc41hX
FpcAA1HSdUf2PrC0oYpKIPxA/sSJeviNFOS7zxLeBLE7pn+WBPzM77Tapgrf
5EuVXB/dnGbrJdJfkda9ek1f85UqyFb2xaP5Wbiu2l+ycRe04rahBD0tVd9u
zhNtgorcCNhJM5AHotWyZ69VRDCFg9UD8Qlv+0/VwFm5/vRBH6/pOBnHcWDo
kChE6NeBQsvUNlj3Si3Q1jO7ENVWVeZpEkVk8gA+DHddaaOcB9ZCPr33JuAj
OG2qZEdAzy5GEroxVogOOBmAB2Fhw8D2HcqVTV2kZwEI4icqjQSsznhsFwcn
xdXcPMN9nLXLGY8GqC9JiF51acddcSnw1GsyqPBSDGsT7sOinIUImLh9bSLM
5vHOGioMeE3kQPXqTxhZQIzDWa+oDKoz9tyTk75KLWjNX21dMcNQTsCZ0rhr
E+c8w3qUdLc/pjPcQPl6OthDnhWw/hRin8Kot5mvuUQjVsNkE1BqbojItJi8
culkfNmaeyqAJiLNqxfoOorjckxSN6MKe799r0KJd+KtmSNLdaiAMcuyKBq9
CP1BI50Pq+oGjo3azKrZnIpOmv5oNLcIzDC1dTv26kfqXiX62XeE3KBquC73
S4NtxUyD6IDNhEsnUlhVV9eLXO5l407BxWf3nqytDvcfmjBETf4IkLq94eGb
BspMlzVG/Xx5LSm4usLh/ntxqNu+eUk/zWDC4jlKvKQuc33A2gpgXGGL+6im
Ie4GB927CI+S8QBOUzPwZosCQMDTkYFXEDhUbW/j1TnR7zgc+eMHuAdGmvdO
RPnBGl9UVHTs4Au2i1kJs0RSJ2ArqiD+xeGH1SHO27ddVXt1vPGZzawj7/Hv
krRC3foEjXMrirjb88+buy1oMeU9+hH4rn9Ns3OqgRByw07sQogwxT90BRfB
d2qE9XEaMu9qdaHSrOPmsCRrdzDBAGn1yk1njC3tYyAOD6KwxSUcmc+qxf44
SPnzlXFnEH18oA6EF5vYiUN9nOmhDKxMOsDeid+Dzm/VZuMeDlH7zKngP+4H
qbzFaO50B3yT8YxEMwlxzfyVjLBkvl1DrQHUCew/X3gqZ2xAcJtUihU9fjkW
O22o67dyM7dV/j6fJTZ8ibCSCbieDtADKBisrb66PFcKqvsRROvnbkpjtdTJ
4WJTq2y/UZ5SGe+bI4EFuYMxD8b/SK/SXSazomYNHK8sFZSre2Wa048+qPxQ
TZuQOsktkHNQHFTu0ahYtSqpYOTEw5DIFXrdS6qrZLXPDiW6HhythWJptP+k
3PtfvVZcYl3Um9pe9Ee/QM8g2e1XMRveRh8njNx7S57NpuugRRoEzhp2feVV
EH6gckK6XmMyOiOpVjWlZTqJYNpJwxJBEdlicV0yWgAC/FJyg1RGfeE5dobP
NyCO0o9kO2wu6EDrkFIDb2onj/PWh9tQS4asFha6SqrUBLDUn41OpB6d8jLN
mc66/x1y4MKL5+cpM1tt4L5MIX5/ofTzWrgUQJXSM/QQ7HNg3Tw2lEEzIoze
YcOvJSOc/jE8iSFvqg6aK+Yyf+VFpuhZl/F3VZfOePIkDo0TnEJHdJmy+TOh
0XogorbTMGOkzWAZTWRIHCaRu9Vzb86bQSDm2e+aRY98/K3JGp7D3p5HZlVL
DlZmpViisPzJLYRZbCsJvrQlQkQ/HCDAGkW44KAY6I8s4bigj4gTb/fvSf5s
HnJtsN6//b+B+CgftX/GrqvEXVtOGlmxsx9YtT0zMjMQRyupQ4PGFAwHOrMM
AwDFWxvrnozdSeuihXyXhpIDztC1NfAqvsENZ1RygF00Dr6c2SNsYNV7wOwF
M2EIB9asDdcrYlw/gx2uApdfT90r0GZhNtc3yK3W55Hzl47apme1eWgDb5ay
C/Y7HJS1xIGtpU8gDmHG8megEJoig2QTHwk8e9tH5V/glwoCRzdaAyhJf41m
7anYErNq9ONA9CYc68UBnmkGnZINLZllZpuWoPwYSB5DWp1pCB3ar9uR+d/0
HYcjbVG7yBDYa8ZNKovDgpfro08QeOafaibhV7TXm5eseaOnPvzNmRCFd3Vk
hHppyviRSIvV9GfpJ10rm4AyLNLejzUA/pAYK4d+1s3EYPnikfMAa3VZIICC
CSsp70+mga6Bf3tKJUoT+fJ6QbDZfHvPQ6gHC+vMcMjq5gpygMqNsSoyuBxD
JY5M+Odnc+vE6/l6g0IYcZZDfS/+xjEu6MRXf+UsdnZZqSvAkEVqIPbrpTVd
z4Yo/g06ECUE+QwOuRwohmEbshBbXl3TJC9OehzMsSla0XnIHtG7YbDuItwS
zqLiDAivuAiR5q7RQQU3rtWF+3+uJyIhvZyyZKcJQXcdeIILQS7UuxaMGKQo
YgQi8bv9TUo5AKZlOuRg6vExbf1h9K3AVCEpOTJ+JPBIeSmL+Dw+xlc0alF4
HHDE05oIqXhBN9MaLw1bxLer6BGU2+rdUX6EVD6zxSoJtQjX/muyqvZgVeXQ
wxbBMJl6RR8JfQHy6lhmLo/gR/4ooyyWJjw5+uSuD7lPtgzY6aKM81E5iOM6
npwvyrrI1pv9Zj2AyE0gls+PNjZmV6adwr1td7A03hyh9lv0d+hCGMgK/yzl
ynhBJujV9IBb9afGEcRHTesx+JmyMJjVo+PCWIvFZGD9XU/ef8YIFc32zcyY
R9rz4lWlHTgvKQ4lpdUL6uOJ7cii2a1cs6cWdkXnBhuHnSN+IO0OpIXl/hex
PfUuSradCcDW6Q1jNSFx0X2EU/JoVtXCqY85e2MW9cfIVZ/v7LFxiSUQajql
wqZdpgMI8yK6ErmRKoB+gfrFbphfCsqOS0+Od8JzpwYjlKFlGF72W+sd0eaZ
qToIC02Yv4bljGz4g4BxYltVQ6PvKylgLdGHMq78PXsuuNNAHXHBsiWb0s4G
1zR4syakxqv20RBRcGlm1Uf43Izdpld7m1X4JsNsgbIPOiUeUalD3SHghKAq
9DqzB11+DfsafDDqR+bBLETaxnn2CvllNtBA/2qk1MhGiREudbikZ5VMfW9b
nwZ82KONVI83lmRtC3/SA7+1TiItHnWpVd8niDPdxrwtkuzYADygFXTTnfk3
AXepEcl3KJDJHur7Dpis/tbSbCxGlW2W3r8vj4Qt9XnYH8E8Z+HxgaaWgBqa
nmgyHkS70iYvKrWHmddAAX5aqPMFeSrLHNnXhcp1g3SHkkn+v1NWo540nMsb
EcAm0lTZ9KuYjGu9+iryYnPUXsXvg0tVPKMS2WveOmWjiiliTC7ZT9kW7sjQ
oR6oP53FUqjBFuoxqPzI8nDl/Qu5D2M2EH95+3h0Fwbbozoh3VtPf+0iccy/
tUGNQMLiyLKdsVkOzmS3vglL6D1wKCs5CswOKTdJD7Cm7T/xuYGnBAqIkvM3
fdLuG3qTYLq+kE8LhqJEjb0jC8KqMeD2LPZt5Gclm6iRmMJHZGKf5qDLL+KF
Mo9IEXgmNdQmPQPRsx9IbPTAqT8oQH/m+CsRqQmpjhk51tRRtsxcNniFajYJ
Yx8J1R5DEWJMVZqeHn8lPp6g0BBgfp/RmoEozKX/s0vU31XlusWqD7EUBqB1
zzl5KP+3GC7LiEJ5w0SyAHtx8QVzRwNH5ZGs2QCAs4vAUBqg4fehv7RPCllO
VLgFs3pA5PjSYcDx1tCN58ISfoT3g8MNO5hdBDHrBdAA7aIeqpfwA92S2zh9
kReI9CeswCF1+YCqsYjc1WkwgZ4BxShlheQEJdKC6CpgrMF90LBZIGqf9yaw
WFlVyh7erGyolM/nPmIHpdmwxxqKpHEf42kSUE4hRi7vg9kAeXf55t04GVMD
e2XdJxiIQ/ijZdw33l+N2nYuDFLQ5hCYZZJpYhOPTAKJFlPiGLX6Af/RCESK
PkWZxpW21Ghsbi23Bt7ZaePRlRzDu8Rw9BLgzNbsfkYdNAxlHVUkDIRil89B
emIqsXBV8/Xod988THx1OYsECU57GK+7Qjua8V34Fd5UM8z1K08cJsTznhBH
Fxm2nF1GMe/0LQW9Ba5i1KfwqOYUV6Npq1esk/V/QxgsBysb3/HCE4ohgSA7
u6xXZIBg5o6QSnUOjQ4P62TpHlJbOzccxPYOpuXmXZcqxGHNrqKTAexQHsUi
Vk9T8/oZHiXb/WnlAMCi1YuLclDeNKbFYrdMGlmmRAIOA9zwe8cIiW+RAQIt
OmRFtg9v2+QhOCoQ1DkP40F1ajfVK2dDT2vY4FtqMecl0uk25yIAQG8oxnU5
ApwUBn0y8muZyDfU+4injySKGnii5QRFHLe1sDvFJO4uQUbAAEXk9YHaqGEF
igC0d1j6WxGJTe2X0w0Xa/7Lbz6Qli/OA9os0nPYPp6uB983lsSsRFV8sb5Y
HWfPgI4PUotX0ZysFNYK74psJ4EPYZDpj+vzUCyohFUMVUAcncKfqp93x5lf
LagToOUomIs1EgEBtdqYWEfIAgGc4k5bPJmlMiTfO1dbxX7gFEhCaTYYPToG
wkmwHI8Gkc9hH2pHDLKMIO7Q2LzV7d7U6M/VcM6q+qF1zHlURtvq1GaTA4rr
GfqD1M7pXlxdpfCd6MnW8RPsicJktZeM4pl+q8d5yzeh6E+KP6T+SdSP5yGc
65JBAgmWAb+sdd3CzWqsGfXMxEchSSJEgw18Wo59h1qEETuqO/TTjcbuJ5gR
ECr4u6I6HSLOcROxP46vZIfMe97Lt89+yghrkhS5ZZpK6czn62c/AUgEy7S4
KB9pYBMzsaJXptgUEK+uLm5YViRHh9+rHZtVxF8D/xdDZWgLYx5oW9PlK4eP
4cjFgMrAS50WO5ywWA0KjHnXys8u+8B8xnU7AY0uYAjPtEiYXNnOPKlBt7bx
NuZlBDoKJiIadMpSMhq7E0NIXSY1OgC7gwqUym4r5f9lkmYjeq3lNxe9oktd
uYCNMqYxE7CQEmVeiVLKneKfY5PGiy1GhrD1YIs2jE4SFydJQw+bZQ+h0q2W
ZV7O2lfJ44A1h8xuIW/S19/yTzf8MZzdSNUuOuk3h2s+FbPIlHSXGW6bAuq8
RXP5UDzWmRAmuLCRPGl97/h4gNlmHYOGtx56YI9U9n/RydSIuyfWGb4SC3ES
+lG+cw1j30MzCmsXIJpVzpl1bdLsT3NbQDcoQTvSBLmwfOR9DAONzc86Obct
oUEK1AUy7zzCd0HM74OKTwpMO6TBKzyus8PSi2VWJ4sTqeS1+iAX/IUAJbkV
t31uxMPFHEn8EsE+Uf4tHx2rheIVYxvnFtxpiSoEQUJmkUwJgqILPljPsHcU
4aYr/NU6aER6LiN1NzFDrPQ5b0byhz2l7/vTyCxgkLCC2RUdd6Ubib26FZsO
pmVG9WcqY1minpFG95Y5QKvl8DAkUjNYxrojUlTZCoM1+zv1H71Yosf99x3K
rHpw0Td1jJII3QfRbOqXWetq/yI+l41hIHtCYZahgdX3cOVa6Yt2sIoCt+XH
mi3yC4lcB0AnjsP5It8c8dmGEHzzedwd3J6DOcwfDvSHERMVEitflWiWQbBo
TAEdLMI64JsiqTgmqQ8UzO8hrI5/WGLr3RlZUx5vGNEkp12PGLKHJ78UJBSK
Ir/9Q0tN2ALNWSBsypu7O7xk9PaYxQT6K0sWCOOVuw5h8J8X7mvE/2hVRm7g
Z3v/FLMO9AyY9mVU9EIgs4chWgnS0kjbGEIJw7XCXfREg8BKniRVdQqp+6ko
vG6RRidJ3+oZm3itgsP0ketyAVaDpPb+Bj/xuLC/IIsv/DuLdrqU3SxjKFoi
9hxgtLfzh8bUJOFGiiz7A7ljV2n69C27mVklnlOI/f6B3NIN+gvTfIx5zdcI
X67h9opEuEjVBpJPgGNxcGwIg9aCDoAeF+SPhpCexVAtFY4YR7VAoikywrBn
Q+GE9Ivyq3fzE9GRjktBXx/cFqphfQW2Vkn7u4hfYFWS5yueFI8kyIj1AUhW
4Jn01NPoJBeNyC66h3sqRFf3pbKQc5M4lvWV4N1ked8hLCAnwysBTdKIBS5K
HzrQlH6N2Xn96RwPALWrB0LdE2U2yp0axVCfqA1g7kRU8XmwP8yseaE4gdLT
dGuzbziiZ30NHmO7kcHuKFAHVdlWzF731DUMK0hQ41+AvjcsglTYYSaLIsWt
L0Qyb3LUDqfIJ9LiN56aZkKthjItqyrsE42Gtlr+5v8dsH7jXAosftHFi9OC
nkYmEpLhD7ghtY91LA3jychtcQgCmvG9ZQwUWEL/MXNa+GjG4WZ9rPzMXgGt
UDd5mu3cNtGIKq1DgsKR5pW4m9hOToVB1uxpiQf0edvJFgtMr4+3KigRKYr8
WiSkNxwTBWAaaeP8s9hkrbMKS5lhID4Mw4DLNnysjTRezQ3GcwyzpyyhN5ZG
lAkS4v+kfuYRCqc7OH7PuHc5UM0n/CERXAK/h2blXSbWnSnhSNAX7W1Mgw63
Vn2/JwEkDeygGe2m8hEA0R07k01DGOVkLLXrT1VcoqVL+7SwLmA8VZ67z3m1
3T+oOel+NDOAP5mcX1W1tTV5uA9gyRVZupaVJOObvC5D6lPNvEevAklqrV85
HLz4d9gNjmBNywtTfz1OcAf4x1Ujf2sja5nHAXnwSKGDkC17bBch2zPeKEbe
j4vF+DdJcBXePXYd89YtUPQOzOyfKJhnVPX70Sj8Q4WeqYX5NRHzMBIhi59x
v+IgZ58/2tH0ib48RHvcH7/ThFD+Bg1NyJVKaCJ9r5EIAeu3UTGeoyzoD5N7
oy2zCfNMoCtfi3l1n+7WEK1vqAYUfKQ5BIlJnwbqTh2bqFK6SfD6iGL9Glor
PAcXU8rFLzL4ijB1QdylgVr/rWI/7GNXcWlAaDkPLYIjoI3acNIPft7LAlvZ
rnAGGT3BX7SJGeut6OIFDsjm7LILKQQe8zTE25Db5uZH1m7s4y5Z0uR9nlZS
GoeZbWqHNOzDtVhW+7+hwxnFNRy8j/aaRFrWJc9p1VkHTayYXTVaTlhL8PBn
njXY3h1xe3MKybWz76qrL8nSEZG2l4eG0Rg4e1Xc46HLxR+klHXRBLIl3VBp
veffMIbPhDHnB6xXaVr11RRi0zDzBqLj8zHcmSd/K+veNqENdcM/5ULqTYQi
pg36acg3SUwrcSeVbdLc6uo/GoLRzyrUhTzqdi7pQNPeGpXhlqGRVZ/TIMqk
w4V6H6rhu4uYDrV7mxXfI4RHSlkt84PdVOaA2RzMlV1I2GJyZ3J5DJ7ZP250
IGLptAi3YXGh3E9Dfzf826glCJNIHkn0s/BXWYZ7r4hokIlf7qD3BjS0KIlJ
Dldk8Iw8wms3odwzbej5TYLkvimVOuKWXg1xjujbqlVUqJ3KZN7JgnEwYC3D
lPm5nUGHx9LXEUBgyR8E3oKjdp++4hL1HyvHIrHkXtfT1flET9/FH1Z4vjlG
4DKexjT1i2UUt7qNPFru/x7FN1qfUhq4aiVanXLYW9Gu6PRbCqFDpuEZ68Q/
CGF8RaBN8FOYZ8t1COkZ+UANtu61fRHcS9xnCBU3zg5MUrEGytPBoT1wYfuP
Po7w11NPhWf0FAJ+rZsreYreZyL273Pjuoi4CYR2G0gxQGgRA/jqoHw2/MQs
w0ydkpjg3i4Nr91HwSkfo9vsLvj/oaoDVFCb1PdBEvSHFtKsWpfZDHyjl8Oy
14TDHWvCpGvAeq4p0mTZhtFLi6FLY+ftuxkqybHqgViAxEEsR/i7PKjOQzGy
VJxwlC+JQDAftD7UJqWRRTSOCBKL7eH2gkbzFDUCSGIf7kqtD4AHG+/IzQcH
eOkUpTtIymDx3iOOQwmpRl49sPuGLyxlNj9n0vSQAv8O2rjXa33+fEV2oAw3
3CmfQ2FLbfiJsHCVQUH7qNwI6SV5zZEVphFaNShhWP97ZGKf9prj08vs+yaj
jIlVQtu+9GKAJxUJ3yJbVA20jJ4sYg60b9Air66NX/hDN8InUfluXzD6cjyF
qBkoiVCgvl2ohGxmbLHw7PWyoFHiNMi9ufRJDHmsi3At19qTfCcSGlNw/x1y
3/hKBdntF323cjEw4VMgyjVB8JYEUE0VjVNqz9Cr17Gbep3iTUvgwLHSAYxo
7alQTrXh9aIn0/0QkTPZjUUaoIDjnDOhtKxVcuve+8PPlTKl5+3nCZqqJ0Ua
QoLuHYiB2D1GJyVEGo77gZA9zNPnvV2lYDRGVRj5GCf2wNTWEfgQTFgeiGK6
1Jnl5bzA5BC4WQ/OV3qrm7yX/4xG2SRI2nfhVAlJ7L01w/XfCYVV4ZoH250K
UqSbXhtxKWl7P0gFdIef+3/YQD2DwdueHywq4PpWxdD8jnV9QcV6v9MWmo0q
Ia7BM5VZYduRd3H83NSOVPRt7VZY3WHVU5PQWPmsGeQ2EIML8DIBzL7PV+UP
vwD6Wjv6nf5J2aH7G4CvNH3PAKPRo8vrNSZVtxrdhuwMXR8RxtdzAt/elLU6
WlLblJInNU1zoSzptucmQJV4oB4YzVFUqqkYI7bwwV4WMziOkEcZkfoW5oPt
TAhxN3j6Ms2hxVSJIO2b8QMTLJzI23QtiCNv3vtZ+JLpN8h7MzFYVFrinRSf
pLKb5obdb0BXlBzWAQAVmoZLao7PdgH0XlFXLkO10Gvp+Zwyqyn3oFb4uwGm
A8eMA38kYlrwDzpqINZ5UFKZxAETPgkVviP6gxWx7Bcddo2m16UPF+Vxw1py
OtbTVDfwHYyzUQ+KnyZ9n8noFcAXtTTFc3GbHOUoWJj9yhejWOAMeLloGK8O
isuzuq9zFm+I1SiVDMPLYR7QWAaxu5yxLOW7Kolej8QIExJZ0IyOxQN1Tghp
eHZxvwtPbXlby5IuBaK+DKD9AOGJpXaM1ThLVoTax804MeSusOvQjKO94uRV
hwXZbqYY3LMMoDitxS8eb0f+c/LihJCfbwPYIIT00Y6J/BNfJGsnwo88Kkwk
jsm0K2Mk677gzrG+ZhqowkDYF86TGDB6AYMPdj5BAqPQCxaUFA6fsqyvls+s
OWPa1jZ7/bKKGFmrkFAoJOp9FeEdslhAgMa1MpOpim6CsJPkml8q0r5S7KSW
n7p8A+seLWl4mih9duKnWva6YhKeqpRrnFNqpuIm7CoAHBlGrFhbB3bqh8gc
oSBO+kgkex9Ibz59AiVorD77KPFqstZXO9EgrVQm6sbKphWaWq+1ost/Ujya
daKmAYLs12+yURYT7z5qZ+DJoFEBTZ4ZGcKFf5iMvYl9m7sEqngpWpFY9uIG
/oOuWHu6jbIINZ4HCd3AJzF3gDBTmYRKufZS2xmtX7eUDCmDXLho4K4nZU5r
/ENEXCE3tjFYiVhHC9vXi5n+IEhmUchre+W7mtSMnEos/0Oq54X0Ffk3iHRb
ehAxqwo0nZI5FTWUdvuI7sjiZMD/fL+PYlCrV9ozkvLvcMbwaq96bwjAsPY/
I4LitmGao7Gc+AVxxhKzG4Z9fy7f8cH5VA4FDwpZwzPCHwA4cBkbls0H7R+L
9ELjkanic0IViE3DWC8hj57UqlUsfE2n3Q7QIZOWNTVbH7VUzE8tvak+m2cF
qzDOtgZqGLYNx6UJFVJpShQQeLUgVcWNRWs4jS+/c4ejFl7HrkgAQfRp0cLh
HpgB4hBQf3CCw8AI3OwAJELJ+gqsYXT3rmz2ZzmG2MmhPVigZSN7j9qyp9Vz
eo8Xzcqkyef8R2yFf/GcIwlpRKyqB5rUjMNF4iW2y4bYGs9CCaZdPkMUSocf
l/oPXyTqaZxQIfLzeQ85gWpirrr/AjTHLkmKlQJuW0WuoqHSUN7qkttnRrsK
AlW0SpicwJH0mw5m7H+FFgCWc2AyAqlJkBl9gEPZZLi2d8N35BoO3b5MsQZS
pgSeaCk7Py+DO9F+g8M9UslMmZcPyav4SIPFijbjc2YPruKBWFj+Kis5yNex
hf+Mm7FXsXgL7LiZbOnsNwUqSQstmcW8OmjkVvvV1mdrFKIIVrd4wbOlB95o
g9M8lFLHy52g0QB4UvvxpLfQZaEAc74YRbpxTuenJW6LYrOQwHqJYhytcAd3
E0kV4fv12qYdVdWLjpnjxwq+CajZdMKNSBoRe5N0pzNWDFeLD+XVAXwftLcG
q/EXewdg8inpSNbet8t063f6g9R9mfrWfpGHHW+PKOYonp118dAinzpqdOa5
BT/ZPLXqWkoQ+WrkAD5ZSIoyDTmExiJSCW5VBiZ7TtuOaTBkaYrI/foFZ7aH
/AwTze8alL+iZivOWldrXZwJ2Fy4eEH/XmUcGkUCRN631V3V1eY/Z1hHllGJ
+k4TzKEHUHtol/OuZbMNb4WFI+HixZrstS869IJzrTOnlePKknfRawFewWFv
8cFWwcDPMXtF8VGRvwT1nIaSN7tkwegGHcVEjBQQtnO9+uazZjTF76HoqW0j
Cn36sVHKQDAK28bJHfkTRKm1hiqR6ukhiXzjAzzljvc78/dSwYDtdCwNI54G
rD0a17cO8TGx6D6HWhTyyt4XO/e+SkWLARFa2IPRYxi0mtTl+6GaPraOUS1J
cNGyxq9+exgbievf7okbjEwVAVI8Zc3ELlNr0gj7AUyq2vXhPFM/hvp3LZov
dY9LiXR1+Wk3NcXUZkgooXPwW9pnyd4HQ2pfjtDvHCl3DUWeWrXb5UWIhHW2
ohjWTsWxC5rFMKdrxuep1jlf57xsBalJ+G1zhQzejqD0tCMYNS055vBwGyqN
W6tNd4IFGaJg9+rL3fgjLrs5WxwVVWVcmpFB5fBTkF266ul+BdRhFjLhMppv
qubzN9JqtuA68gr5bg97Su8ufObk21i591NjEMS0AYnBAa95T6K3kPnRhnjw
gddufLZYPACw/XA782NreYz7Dws5mlJZYJRSIJPZ8P46MDVd7rFVwgEOrUDT
57qb2CpyZYWNtsmTXCWjCet65611/vcXzOcTXwChAVgN7LZ1dYJ/U7MUeZOy
yVVQmt2bv67MGC0FRzJMj9TszkxJ259V9UOYJTmEZPnDlnpQyv9cHpnWcJT2
j7cBdc7Kvkqv+kWttfE/Vd9V7dsFwuqpqZOtGplrjUboc7Mxcc5EI6XS47I4
r0npfG1/YGVSknQRGZPUE2DozDxXOgUVgNnTFkHCWMXk9159YeAQ/Fm9DoyK
cj6KAhm55JPPFnnQ2PHDZTS+d0EoiBzBY9KWcS8Z8mYFDD2FMyOR4HgF3mw4
1shFhqEWEb6m/xIwqIYR6A/1iiGfbINlHRGQF/H84ROFWo5r/lXi8PHnRI6x
m1XuXkRUqJd2H6YGGN9Qgsm+ha/TkqmH79ljAtqimxkHCpCunih676ATsHD8
9ccfn58BeYNTrh22WG4B/Ot36TA6041fbN6dMMmQhc9tPrbcbT/3iakTuoVx
TpyQUBrUekJ5ObF/eZzV94F2NpIGuk/VWTcLMG6L++YJk6NLs3v50j0ADsDr
wPK8fQs6e47YWEztHeoApw57JDwVGMkgwLpYkUhg0vmZDIbjtI4B+gC3CCkE
Oq9ZOGAy3bA07NqSNPKAYajMpbhKKQ/igG+ntWt/EsGTqWd2bwPvuFR/s/Oc
Ffi2eZbeJ88o4CM1vHdKAJNCzh0q+gryoi9XPCLvBmrDs3cfFmD2O7LbuGgK
3NjnM1ELUQcuQoXqDiT5OFrRb5kIc4HPnSRnjoF1hFYoPBwQbiUzQLT2lXiA
wBv26JnmtwjbEed7yy2iARuUtSZLhXEZxZWwlhs/XiiO2KTSCdCfbSEYsvFs
IyFeulfKRYXu3P09+hp0q+0qMrtnBqsVBrab5AkriN6zR5ThIz3FpFEj90cw
19cFe/PcM59rXs+N38hLebWByjMdyolv2WyeaDhhDUJwH9yyewnXAnW1vj+O
cAdKH5Rackyir1nqyRJWy7Qy+8Wm6FUyyFe1tQvKtwR1qInCq+vr4sl/lbeS
hfRfnREdKH0dpjsndAqJn1oRdn5sDduxMk+KJbqKn70cnF0nou87GKgy3K+7
M3saGixgnDRQk8RFnHy7L/zWwidzsVcMMJBsoMjn0keZwxETINJponAJTCjn
uNrJ8/rwYrS+QisI2iMSR1pUCNCPop3Ew14bX7Kt5giMbsKGhBRp+wb7Mm2K
w5ajAt0KWoAWPiqx0T6IC2pTotBvWTy8G6Opg+RUY/xQCz7l2+NdFe4/Hc2D
TuDk8MGsANNFyuWkYkzjJAH5dzP9YrHxqqpbA5iKM701zf1aDcmDxLfX3RnA
HIprPlrVUJ+nsMXhb+Ju9MCTzkMEzJi23uIpbEsaze/GUGis1RI8GNrF//rr
BxmAwmaPIgaNSymW3enUtl6Bzgy8Wul5/Wr6Gb/fjCc70wsG+OIPNRU8PAcO
CkgLfnZbLWZIvQplOZi+L0BHS1KWdECjxIL0gBCc1RU/LvZFQz8Ft+Bll1xP
7d2y/rDYwODKww7ecT7JjzV44R/TTLLk10jOS0n0zLW3EexF/OC9UeKR5iSA
6bceJpiYiyXhxEdx/eO0fyJgeqOnGaLQQBm1ixkc46Y7nDuWX+vB9gvroy6D
9eutXBrPsmRDpCvY1t6a/1D9HkiBBHjuQLOO7ZjQygNqNzJHPQXoSehkqhEZ
VJoh8Zky+oj5pFe/I8r/xqZMXbG28Jj2+B5AWppWqCbHM9KilVMBZcBoXixA
20xYayH01/WKYH8Qg3dPjLLOGlhwhSjFtNnbTLUy3Q1ouayjSmqgkCGy0u5D
P2oBt1hpEuska7f6T+/fBbx1+j42kToYGzvwYx6pSSLoqxrRaNLnAkswf109
J0kf6/hsSBhUfFQXG9k5TPDBwxulEKuKB9s+LWzl4vWljqMNUyzihSkhgLCe
dfIL4OYAMsowPYV0SsxPAU7fsHYj73RsXwYr92LPAUqos2ZmE3LINbaeRz7d
n6+0RC4+71FtZyaDBwDEP//yxsHHTuTRtBsEYropnkUDd/dbzrOtCSZ0JZjY
cyGcOSOQlV+aCpCLiceOi/OWPFor3nuM6dQNL26tu0hQ4ez0zWZQ6P5L/vGd
ox8LOIDKRsOhG4MOQH2wD7l539F9n6bT/rZhB/yhr7Fss419B2oBWVrUey62
bGY/ZN2dH2c9Uw+Xqyuo0sRwM877Qgt/qEupKRIf0tC6uJu0WQq1u0EnN+ac
aZLjje1y9h84d6BghrNfT/5vqsAnPixiVVWRq7CEr5h3Zl0ika0Ylu1Y6xnO
xVGTOTASMO0x3IEKVcCxFHiW/wsXQt6oUraCLx22Rtw/61Gi+LUWVNYyYlOz
BOto6/P9HYg53M1qS3Y/9UemS/VF9kdOGXIcO1GNJef14aPg6bLykaRhBUYY
P/xIFSH73t4/sZm9xz5aVp1K8NoY6JnJp+LS7ej6x58Xq6Gb7zDFz8ReyhO6
OGUDhzGdv54ydcgY6Bvq8j0SUVv6vUAg0pSOOFbTtWF/7XI/lf/nlOgbON7g
ZYnct2qLQZfC7a8+LakHkAl31htVDGI/UwJB1himAzE2n37MVSpElnf18/Y6
j4ZDqQtaNISQf/Xd//9Lu7DCWggmTNxei8QvnhMwNlBiJA6MhZfaog8tO4/T
jylmpc2xtutGPPZIANir03ZI4GNdfNMD8vxOM9KSlfH8FVO7ZZcJ8vOLeEj+
hRi4p60+VvXpYnYAdClyBaZCHFfCiJK44C6FaocyH4q4Hw35hwS7boEd2WNQ
KJ+K/lKZ+AgWF9TrBPgSprBb5KomHYT8WRokJP2r7WIy8/r+1U20ufxtqSa8
yKCIX1cWVRgAubzuQHIxtE89BaN034TBPh8jnfL0ZQj/w54RYm0diC6CVOQ8
NToTJdOHKl99IUtowS4xqSSqb6Ukma81PXisQzSwcvrhD12EKZO2idkqWEbe
BavRP6JpAgOoUsyyD6Zw80ImgGwN1cJmcHCnT+ox6rdM+lueXBefYnFf5w99
XY06f76U2Y4ATurPpQNJ4665OMKIkSHVV2mBqO+GuqkKfuK5Y68vQ5c9TZA+
QZJn4bvLbCrh7ewtNxkBJtJ23I30huTLAd3HckWZDEnTJc7/3KKoU90NNE7Y
a9TD7nXb8uBqU03Dqal4OKesDtY52QK1hB6tpFRZQtF1jspWYJv8CJXBKNAz
tZA7v3YTRCUA4AptZt4HSZsNqdnBY3EDbbmLKHJ/S47VYQKcXwv4BjLgm69c
4uwRFTLM4cBDWj+qfFsutxNS6mJXBKBcjDveSfD4awGTIrxoRWqkcF4koXqu
TryoWuKYvbu6bX5IdoEag1Urj4LfLxHscbTUEEKzHtahn1qAsB67RBvMEaCq
5WbnL457T0/VOn3HYQ+8kKn0mmaYwEusD5bWTwSfiQd2cao4m6PsQrleeIWj
hhab7h3lDkGn8oT8kN6lcI4gm96LFQ8iYvhv9AnySoNd7LFMkET0qSCfRWA/
IPk3vcd5CvAq2eXBCCRGiAk9bEpB3IKTjzf9NI/lKkc8Kl/6pberm0Ct4rsI
s7ZK0VXwf0Ky6/u2MefR1Qhc6BK6Lwi7mBP8OadQwoIQBIKfY6v7tkbsTqZP
7ebmcI5dQgfSJjMiYMIGDVgrR0/HSVTs2IfyAgwMkmPAlIItPJhIMIVQgGRi
mmw+JTO1mgpSY2uEOVPcOTOUC8wZECIT1PM3lhPB9wLrFI9YJ3t5pu3oUgWv
1p+qy4CPNRVS2+8+zYVNPD8CsStY2oQtw1fKZSABPXOiOAOcekkPcBBt9Rq3
sVn5ahMQ86npfhXbNEL9ZlXw/oJCXNXVA6s3yHdmqSqSnPM5WDYqsw8qjdnj
HhtIJ7Tk8m+Qlmmg20LmhKlzCQgCgMtk66nBEseDskdwQtaZIEPnJLKj1goS
Tkw+DyeVM9e3A8zgmyd8AJ4/laDK5LLnUcQYwQnk9tvWSM+OOb8wxlbd4/m6
IXTOulFYJmUEwZ/5ln+cBkt3jmU2ov8s9nXjPee2iO4towefOk6p82gyJ9Zy
fQCl6RhM2/KD6NospC6eqqYd64NPUpiOpApuEOTBu21pqp5U9f/1kh8Q/G+Z
mCWTR/xZKfgVMYdh/5CIILocdrcZbBttYrO7FmEAlg5E8ZKOmC/fMZXAroSc
ii5wQA1Zw4QLXrnKXfaDcKjxF3CmjqmCeCeJNGk5VphOMle2EEKDDODRhU3I
CnOyWwePI6lAnPo8LPfPWy/yiylZdvr+aWmXK+W0rK20aeZetVCgpg3YyZ68
j5TvUh2htoiTyTr+0eXn5p/Yk08PRjkoNCKYd4W1IRZem8LjIHpsNhnU/8FK
+yPIjzcPxI9yiYoGMk8qzZi8vzt0zx7v2AlE+gKtBljZcr24iFmnHnMqmtHL
dD45hf1fZK/iCzsGleE4e5iow/kyiJpw3BH7fUCB/fv3VOY+M0TZjNGk4+LK
mNW3sw9G1PmwYxrK+g5VOd+/pOH4e2mjUcbHt+I+ifXJzh75Wkf9eJgemK9+
6adDgIjwc92U7sycukoTimLxAjx6RaZhz8doxKoi6CsIeSWhOGsLVYY0vx0+
wnopAsaI2NytZbXWFhiyxfALa9QpcIHk+WZUFe3DII0j3yLxn6ANZ1GOQ0wA
HIPjZYARGgWP3VqH4GSYOvIgw1wtM6rtzgS7MuYdNFe27O6uTz/ZDTFw6yjR
TlujAtXldtuoQeuyPBh31eynckbHkO+TG6qcXEBkJh+Ug9XLCuOlQpYhmYex
NNtXdkDBB6RTzBB996+r2jgdUUuk350vFZOOVy6DCrG9OQR6jYAs80UdFdIz
HrwAUlJGW3RI2r8QqX6wf9Dmc0DoKdhAeautKGm4jUMO+1PSks98Nyn9ApYi
aWVRq8Wh8kIDr2Jh2kblY6La3np7efEjE7kTPVGfzYnHbFXBtitE38CDET9X
n7UZDZzNB05ksRSg+4slLYcjpsw8lzJ9GvNMmQfIepfOIB+w/vlM/t4m7Pbk
qiImXbwBOKSf8tap+F8J6NFKM04waDGt9znvnHjxxTBm7mQqTi5ddH5Kb7wm
9w2v6HMwkkG3QgC3IeNUOZ3U3yXA3CnWfEzrWkddOedL8L9dB6zkFhtYMoOt
PyNwq6CNeLkA8LeyZSKiBHKQt0a2kelJ8mR8wap20hUq0IW0RBUqhv+2z9Jt
+/U6iZhgM4PM4AYnaGxXbJFyvaiLAC+0lOCPSHrrMZOtSOO1McKWQEj3aT8O
BAne6WnIJfyiebXgbMB4ODcGcg3/3OEyWOcMrZrdzEdty3uGMw72v+DcSOIJ
HhjR84/eekZJDAjMxQMQYdc5BNIArmQbQW+7N9MfFVVY72PU3hCQzXAPpfUq
AYr1TEaGkOOPPm2zl6zTvDJfMUZD7nsWmF0i4w02dQogW8YRhVfQvNi4tN9t
28d2YfGzzPIXdJG9CHADW60g2a0DMTi9I6Su0vmV5ZicKgmbtSv1t6k433YG
NX+1fhcXt+CcbBLMu4/hqscgapteZ1HNcEeiI8izrNVj/w59roIdiKw2k80g
3AbsVjCfyscjZdUMGkcOJemkb/Dp3M4rfXgWi1ET5W1+wQLYmSK7MaZEFirW
1fUXFs7K5JIIY5vF+792dMMnMZf04X5DxsSsyaAdtUvZ7XimFuZ5WOxlgPKi
0rEQ2/BHdy1BIcp+MFCPy3oQwlwH/Tf7JYuErolfssTE5jg3xtxw8tNyiL5f
9lj375AbrKuA5VKdOF3nx1/95SUCOomHIJrkFNqYtFVkHJWWlifIdvXHLIYY
U78o/LZ0Ui19Zs5YKMJNLiZbACvMuZM4fbX0tT71r8FJZdOhViv2oACZrm83
DW4+FS2LA4Og5uC1LqgL5KR6oEWOQn56raLxGb3xaTXPe/oeVjxrlfR5KcgQ
/L1oCvDFjbf+fS+OPiQedAESBgVEWLJZtT19krZVJ8/c/XEX7N/WuSL/IAw1
o9dXRywj6nl7iSzx2WTSY3qDwRZl8L/K1wJEQ3P2btwWTNByF1V2Y8FBK9CX
P34DNLOOy/5ltb/NQFTCua8YTCONYyOY0B2U2JMr7nB5+4I6xfGJkoiU6C8t
Vo+Ekkv393XzCFqAiUMnfIekxIcECFFVYSUf8Vpo6oGAoruiXTC/rRkHyGsq
Qf0Vaa+g2GgbaICySuNYJcUmU/j6GMD6rhCEri5+26yAty/2b1ib54X2ia/p
Gt6TBETvWrxBJqIr0Mu1W3DWp08n1vkEMf22uL6rnYfH/9CCZ4hz6B42avPK
KKgqDDvmUuJ3zFRqv6PECUfXpa6OvDOW6ZMugCCWHJZ3Ax+R+5DuMo+f1Xsy
jT38qoHmvT9pMPO0HRwe8iM2hbxSXnos/pxdlwAdETJIqGSvnttkJp1IZ9zK
1CoE/8fe9u6wDsAmJ2mXqNPAj6zQRLwQv0eMzJVGUkNWFvkM8LtQCxr+kKIL
obAdt+PLiS2hrQ/8/ZeRHVOiRXxZSlkXQUxqndXnlUJC7MLZUV8mk/bV2dl6
QmITWe/6qs4A634EMu7D3w266b+31ySR6b2GiINXTjpJPZknvycsYhXnWtlM
vZ1dI5qGRiM7Xx+Rb/v943+pIlLjm4tEHTRPs6l9NZTvhGlvlPXDCgUvYT11
4b1RwlGHYb1ow5LAuIM0ZCdLpubivsJGGeyXLfCi9hL6uDyfk2ytJYuVhBY9
tp8l6HRGq0D7hi+B0rXbDqvOawA1TdfN0uv19+nEpiY0pCT2Y39tWF1Kqu2W
m8B0rc7MCCcyFD6iVBlC9TO+D1cmuWgN6rWpJO51N792oVo1oyq1PYcW+RMF
bZFKX/4Y5dDAoqJzGMZ/A9InVJfLJCDaaoDM5WWJGsfeyBh/6RngDjcAu7DU
8YaOFhkruGhxeNhYDnvFUteUWSvtzXuGvUHRMrUne2UJWhlCqoixHmLMEDFd
ckPstnE4/CsirQv9jQqr12m+KX7hjMQNyrOZIjqmaR70KYIv0j47WnZO+DSN
97ezN9fOect3XJRVbFYTf788joQNjWEI7cPkEplqukn6YmFLb8ZmJ2fLAdU+
6BeDrHNAgI2Qq/PX3DwxSfw7yO7WPpA3nXy4jCcXa5Jz/snPGmY+fCZdcE2W
+iASIBK+rAnv28N0XmC6nrEaoYHFWWaj7pPZoLxbd0x9b7jPZdCbofMRHoKv
a5bjD2gmFksjBU28yJF6LB19Ye9qNsAGTQIEUJ8GSem5kVYQJr3BZ2Ie+eoN
1bVtYr51UovAElPH1poS6ZTQfFJELK0T5nvf3Y0UqlyaKZoPf8a0bZd1AjMT
huJxtzaDMBHIv9pgLQs0k572Q8HKAnWcdrAU8SJpATSkVp9M9BOYG8ZCNUmM
dv1AmRiq6aSrPIuR28LB6Zl3hwluIDgDd8ZsTPxrasISJIMbJlYZqfw0g4xe
DmDuhn25cuB4uXxRFr8+NGsDH2+LU/XAUsfD9exoPjQvnJ6RcXN3w8VRqHyy
4fYGh5kTKz0paQnwoaBkyAiYGrU+N6tm3YvyajuB4/jZ5EXk395NTJVJ9WJe
Vo9OmqQ6u2mCBku0bEjf/O6fSF4gorfw20LRjsijvBPmNisE8yOQeOj7EAni
ZNh0ezgxG/p3v/pq+CcoFGZIRXPGIzwVqX4btDibryVs3dQfi71Wd0QJ+tEZ
A5C6tlWd57DiRfy2VMbX4rW3faoXXRXwrEERaMd6DKsKpY4cCkRGzRihzzYv
lrOr1Z1sGPp9C/WTcP6hRsWWDvLMlanQPMdDciC2ZrsYvtBgFiOHVyXE+y/M
i/DJZLaHLt/tZS4kBiyKkTRQbHfQOxlEjHcLdNtoYS20KVA96F5NXNb5TuXE
5345eF7j54ayKDmCmIZLCVLSjcuvs0hrT2GmQNLYl1xgxCnTX8mY5H3AJJN9
ECM1tTaIz02atbc4thv8nYNlapAzW6TaRzeVZNTnC6C1Moj1Lskjkv5jcTOb
k/HsOclHay+D0goMmti0xLTK9up6lwugzW63Db74UiDwk85wvLTmOJL+BB8b
o+FMnKHe3Txmhp3v8Sx19vxEJUWJrKFGOf+IZBdlxei2wl/xtWjXWoxdwerJ
obff7HpNtbie5MPjDpHKCyRvWTzkFHJB44CzrPMwVQoD8ashnLiomHGyrq5b
gxp/N7E2uuiJJfsLHvmpMkZqsJmuRs7VpuX3wenBNm+GqB4I1wlO1zxoB0Tg
CUWwhHC2t4YuCrTUNjSPoViz9c9JVmy/WEyWrlzYJ7UjyXw4bAkAn0d2ILu1
1vtrTXMoNYNXECaaxrEiMfJuORB1Iva8YP8/xyLIwzAZSdeWx+N/y1O9Ec+c
ylJj6npX25AlSqhJoGqG04uA7zm6li5h7dlBa+YTem+Fecf+7KMf8r+AMptq
V8Vy5MYpa2INR9E424XqhRWJu+bcWRXEf4ya59N4zxJK2aNKEMS/otmjvwnj
6KpoeRPtZZ4oLUNSW4MjLopYE1DS5WHXp4YtEj7ku9xEdgfYL9v5/iuK1k7F
8aTfM8gAAELn3z5Uhg9+8AbAqfnNWrocvhj6DN5qYdlq2nVgAQi/u6+P+y1R
DnmtBh73NALOh4iDIRszA7urfoOHcm1gLtFtLtNac3o7PqtZtCPkLJWtHf3Z
D54hVygzrty+35xPWaXlri+DlhzD+qBZcri6qIEtmFj72aGx69Fa0GVYNw0Q
8Zv54Tl2giKVb9pIA95mLuVXtmANekwpUmhypGatvw35+VSG2u3b7F2WugqU
YHE6E7vHPEh93hAxm8PGcYMdQjiuikSFLmWzgaJzrxAzxPPb/cz2g6oTW7D+
6XxR6bKj8YX/WwuRfRLAJr6tmzA9QMb5KvAM85hu4kh6xPjNBIliFte3GkAk
rwYT9Y4cRNMoalSZ4lapMY32MxRVn06p9Vidn87RbuTtXgo3TTRtMgJGo/9l
SXv0J580QaiQTC/wIqL3VV5qK1K5DPSyZFxTeSl51jLjVgI8vXPN0ODr3WES
qzLVd12h/SNNMR3YbD8yHrGuVeKD9WjnbHIyt/3z3fi6HLAASy1HGCwfxiJr
D/MOYbUlV6q+jur4kk+Vr4Z1S97W84smfsdJwqT5cPEMVRFh4ju6Awbt3dPv
UABMg62d/HOeci7UUXq0bybDyol7XaOqUqk9A7M8PVkCygjMi0AuJfEEwoE7
twg1Obh/l3DKY7eMpjMZPqnxKXypltkkTDfm3XoTNfzh7GAkVLpUyPx5zPlb
KL6IkRx090GlD/II/y5K3yBgDWfSS8upogat5bFHSIG/QK2li9cKSusmjm95
u8WuLG+dmRZsKTreCqnAPgQG0+/3eiI2TGVuBpBfBk0IlzMVnDdpc/mlpT1r
z+8RRlTkJuJGkZfrRitojV3XWrLp2+xjNkcUT5MhCpKcDB4k90ngqhEulWUm
hnOg5z0we+J7tfAf4xZjySdTzS29XWpbRNgL31+StICQC1Sl6NJSIWNHamJx
XtsKkcz7ACQp29N6sWoATFLrYF6fqZXiulC0kIF09QzFgnskKuTSNA3/Aygh
nr+f/g7GbFXqWI0PIwCdSbl4tBJfwV4GaFxohOdTOqrcoeCn9LtTZNiHzBtQ
heKUDfm55WQPsFfpTKiVtnh646oQpiXpF61iICxEd6TjX1n3OrqhrUVKwPsA
gldDeXyCqOwU4zq1v72d4jRNxHnFXiiOaWUnwaxe2q5I3rfapZd1J0qPoVKs
/rqDB7CCB7LwxkWKx0HZrP5WrYcyWFzVpdNaQCwp/VJzZrRNS7aAg91Svciy
SDEq8IN2zZR7P0u1i0ePaTJrXUvEuyQ3/fzmxSdHD4K5/6Z/T1yxHtIWgKI7
yvwufVCbUsvV76jZ7l2NgUlu7jWBHPgmjsAR5UF+1IaDpN1RplCKrhNy1oeI
DQJvyAd1LKdyB45QvaQOyErNKdMjV+J/1+zzEOucBLh995A/8zox+OmrbD4u
k8rZ3Fx+KAFZZFawu+jJrIfxDD4+cUCzBRFXslFheKyEkKN1A2Q4WGat+2YL
rUDlR/IcLBfV27mj+Uj7WSbEIRXzBlJ43lDp9U5ToZmmOG7EdkEecXLAOYTV
2RuLIbqbT1ADoy4m1Kvs/e44FlkzdxPQGmRJd9b8XrIni9U9asvwI9kznoTC
HWr7mgA6bIel9ZjjjU5PeENXs0SZo4KOiGYvLHmqwi/Aqyrc/CAQbRvqLIwt
aUCLgQuDLWNfo7F7If+JuXOtkaxCcKrHj4aA0SH67vYxRJjzxoXWSLmjAsmo
kQQSrFBQ15PWvG9vHCE0+tIeh243Uif9SP22Hzu72AbnkQCiVu3jqNgyarRf
8q69Ymr849yGkHp0JDBlVBi4gSeGDzP6zDFupaGkhlWcSB5VKYgLVnbKRF54
cHQL3937D63yrBV9bKFm8MBK0r7g6c04IpxKL42aqkgpLXhfaIJGSCsuPl6o
msHRC4GD/BSkf18xpPyoJoUKkqT0xaHOGNDab/fAjMBkpG/EjJkfq/zfE3XD
Z299ygNsLldUZeWqrmPjiknbOKK6WkyvOQpB6DyJ9k7F20BOVWAMDR4Mw+Lg
hHeoUOR/JoHVYAXDcnRaRenIKPjHCRPwxcF+A+e0cdN3ueI6pv91F2R1xJkd
QJhhS5e9VubaxRAALXNqsLQhLROyJNjvKj+zmHCYilnOd15Suxlq9OW8HF+B
IXJG5GRN4EH8gLxL4+ftWN9XXIaUp6hLFWLzQ6y2GwaLsAbPggrI10v6Uyds
jKan9Ub/WmAXGvmuO1/fiVFkD2V9u7Nlwemq3YdOmc9Q79mfbYH0VJ6+ieDQ
6e8+DnmQo+QddAKNu16cVutTtzZYq+0DVTf3SIwIx05n4j97MclQWaKp1gvd
eFlqytgjA/qgK+ObuhXzODlm/EiKZ9ZJOBTDY7sPHb/65hMKtpODiHsmvBSF
2kG8mCOr+i399GTR2UPKSzRJ/FXFq1rouoINNLVbosu2RpRMzO+9/Te2Ryx1
iXwsGn8sjejDGmfD9U1WRe23neL7hMcpWO38H0HyEiIU4DM4aKmnD3lstPSn
8nJ5MCUaaEEuDyRqNNvAgEykEqXutdg4tdqkj/Uh4LL2SneQDZacBSRpNtdW
1vVcjINsMHU/GpNWaLGfgDDFVbuoBjJZAvVPp5b5yZcT03hBCqmgxFRxRLet
4iIJOOMhMfdgTt3RjHYV5KIAzn9COYcnuDOh0UVRXS1U883gX+EHa6W9TlUz
sXNjMXBbjtZHyOyVaa24R7XsQ7HX/RvbZrV6GgvDmOGEsp1H436iBuMLQEyq
FTOhOc7SIG9y9rhcTMX3qBDsx6Xfqafn7kzUvcNTN9I5T23c/eweUE59NOpr
OiMzdp7JZiUq/ne1U6hYM+y5cAqHSOuollQNU4suObmJtg0xTuEvWQpnFxDN
qs5+HDjRV5UHuL/gceKI6BfZZMouKbhEbI0TSeedKwIOI0XI2tQhLCbcapJr
VRNvBPPoDoM9Vh+QHh88dwonaj90Gh10Luj/LWG3FyDQqdJmIfKXxWJW2OHE
SY+w+G/ibhcji/JfuPBWauj79YyX50GYl8NxU2RfVmHvKh8fyTPf8jQRK5pP
U9e6GLlZxwXGMxFB9RaU7ZQTm7QFMr2OkVETex071oHSTi56TgL0Xut7M7wm
35qDTiFPMkRUzGrarOtH1N4hcXBS/uWRJQ6djHchtU+KbWDVoXGQicZspCVw
V8XfrCJCbeTpDWwD0m+fAUKQyggpo551gfd/EzteBzqR3ybx9p23OrzqNoSe
IeSWHwUTAABEgAWwm34muO8B4dpT0i9ipib8x29VtfFrNc1zGN7uhgaYWuN0
3wWPIr0NHwKStbc6hm3RVkY3nWyvfI6eJUbnp2CbpYUou95cu1FXtOw+fxUX
hSJfqF3tgS4Y/nQJOt7fSsBp0eS0AneYcw+ktuhz3/VATpHpZl2l+fYkYM7R
I9VtTF61rRwTxr1i6d8Tas4iGRuNg9kDAd0pf+Pj5XROkrjgb2g7/BfAOtwc
1reiht/NGkLyfHaMqq8FLaaKDX9YKVPb184i172hslvzyOYsfWijSeHkOLul
r1dBPJi9PX+yIlpQSmyFY8+tGGLnsayne2xEq+MJvmZwCsgdMiJLYcorZ/7T
SkGMrV34IjpAo6WVRszqd9BK46KK1qPG6jDjPAvDdpUcQn3XVBgT15dR4FnM
jML1fsYtdbNNYkjZYbZZwQm6AzaO2q3sS58+pwFT8XCNLooBzPwwiqjFrnzP
4FtFH5NhYYYebZ5WyhS+3J85WsQdC0sbv/j24tqYHxX9lSXaKG6F1qHXv+37
h7qaZuvpADmpPDlVhtVLJ8DLlLjcgzy5PEW7KkU5+cRXR7piwEeST4OaMN6J
/AmvRYSzcbSuQeA40X1u+K+twBU6X4A1cQ2iHGkgR3jSEx7iHq0cuscnRJjz
23E5OY5VLC6tVv2G1BDm4heKRFON+7E6irYHnWz+4Sflu55iX3eDhMYoqNrp
RkGBKm810JeJkJqETCcBJiRYbRGWZyPi56QUqZnnljvKYio4Y7ypoZvY7v98
jH3a1nWH/aHppyKv0sciy35iTtx+WfuQofC/88XNomyVvpn2rAtxuW/OpaWz
BlAqX5ai7f0gM+FR1An6xgweHRlNWQeLiLTxm1hJyWcpmQq+lVA/k0gCXwlW
xIQQymucs6QXu0N2U2+rA85ZUMw3s4R7k7A7s5N4OoLvMoVm7eh0Ra7b2IU8
Etv+E9kRIkgdR/UmHYPIIwfR7AKuHj0HIh+gXIOlbdJNd9nFSsuIVq9B+03K
pc59kQpUpA3Gp0OFFeP99wW3Qr6FXe4sFV0t6fPNlA8lE6ZKqNXpDIpT9QNY
EirysdC8jGdvK+biXOfXlJVcWEn7xVcBSVopIb0molzHwI5wYachgHKSLHZx
bZuZHAh2O8K+eWoSZhmonL4l7rdvEjK29/avRQeQovIu0xCqtj8d7dMYw7yc
vKy6Vsc15sRzdXgP7TTyoEEoZeeqis2NRK/LJu8nIk21gSW/HsFMhuwdaplj
7EQmdBd3+BkHrvAgvZEqAT1zlk1rSSC9zTgDEVoJLwqoTZHQgr9f8Ysu4GNa
pZiwoGwQUPVCW3rMeU9qROGXa3buwBoC0gZvvvoTDW2OBKvyMdKZAGqw02aQ
9VlzD5O+1OVLF5v4hgAZXSTDZ/+r8ao43jJHKBnjyhwY7GEyUSPeqIj8KNJQ
pZz1dhUgHWjlzZua8GHcnVt7aX91FsJhw1XQfRCkR6E9Wkm74YVDngVK8BIV
iuLEeZ4d1F8vttg+R8lhKgrY5Dva+rpA5iGnZg/bxvGe2GIfhSX9hBZE95RG
r6yq0zS/73vBAGamyezdKZUrl+hI1JkMrUJylPZzYfQZJu4p4p6u2v43CA7N
Cepd55pdIY2xw6cLiTJPrhNkgMxHppBtmTsEN9Jcdd/d2xI2lk9YAzDip3gI
FamLUyMnBUxpEeUabm5SSDpuIHdYrqgMj736YPhIZusciO1q+Nq/A0w7ZysY
7WrozAlt6c9qjUjodHRydLCl4c/FqnpnJTU3Mr5wIky6mnmBdmJvMmagWikC
W8NYtMIkmtXbaxfu/1P65FZEodANoToVSILQe7xeG1mpDQEPs+LvyFnkvEiq
Ycn8xO1FYxrqaDs10eDUKO7LfztRQzQlY3xVcoKsUVhwjs1pKClMY/6MyhlV
H7gdHKKPMrxSg4FyfDSkPG499D+0K0gyg/oX1G+xpzPLP4QtC/Mv1dCvXrgY
M5awMfNj3zvpm+ujIkbtwvs3xPrLMWlpzd2QRnGKTEeVYSXQyBVnNhZiixXD
l5N0YcYx4JOZOizvOCmRYrgPj0mA8ZXceYB2jDsXo3/aYkQVfO50MkIfXJ60
jvRUxcbmrIBxx7vKCxKBszDX62iM8iDvZRxwk9f+nsZTNfEexLld0pw8V7eA
wFPMgUIJrFPn6Nu5Zt3NOKl0jk4Q2sxC0bk98DXiuJftcMTlHnKdHggYxaNE
zHl4IPTICygOheNApgqvEeiYnMkXZE+rktdsHzk3z9IJbMJUJ+XEWn2+qM1q
fpgMkbPgahQRz1Ef9B99D6q0aKOXVL4LYxwFM/j3zSmoJqyes8Pq8kfNcEvu
C/FCIBPAkmqXULOSeIY5jA4tohuSkPd5Rr/FxKtA3UmvmsqGbNBAq/yu/Htr
gkAtiM4t5EOvAxd1n3Ja9FzY+Kb62U0bzAkVLi9SmSGxq5A+1Eqs4whm/rVM
j2rP2Ix37gzjvzVcJsWnOZNlcSZjcgUad3mJeQ8wYf9PKOAFXzlQObv/PRPn
xY9cmiwtIM/AofGFJa1BteWR73NrRuuRhIiHdHoI7YUc5s34JHAlNilE+bMl
8EygFAHlwpqqo6JA+tltDNQG7gcn+aJY2pkVfwuPqpjAu2imjmQWYhSOOdAx
uGJfoTSAbi7psjaUIyb1mZDY/qJE28JjRSDP+mVTmF+zZMwvWDiDL0CUdOHQ
St2ENnzCZAW+ztt9MLTx5LsJF/j23/SkM0sUDkDCmrjoZKtlf8+6jgDk5u+d
SfugQsJxZ+2PNAEqyk26+y9j0t1VTS5k+GFl2c92ckBvXzov+gwfgbbNvxbW
aZWuWFQd8zGtwZNlcX9rbZu+OUbmqQY/kA+geY1gOTIzwiawOLMPDnsTU3VY
46sxcN+9QrNp0PevQOzvGZU56VK7zfEtctmz9Nuyykcr9vGW2FI54/NgidKW
CrjKSBOKQJXS6TELXoHEC0n37+EZlubcrPsfTRey86c6mRj9oIuR+c/TRXYe
cg3k25GhC0l33gOtD9pUbO8JCQrg4Hb00dDjGGfgNdKu4ZVjeRQ5plGlvo/v
QlHVmxUSDCJOPGJ1UBKOSjaNB+NUoTdVuTixR/8fHpsVpb/TMC0MB6L3wHTp
Ps8fD7bVzQCXVlDNwm4Wfn5/+7IGParSbt0iwBcQCiEcNI6opOxTZ4YjC85k
wwnPtjFLybRtA00nSIjU6YdbhWmo7vVISspGZoVYEF3tLmSRGbOcEJ4E/Bae
vTlIdi8lr6wMahmq8YH6yXce68NMcWtks6/gcH89w+Jpl1ytO9sOSwpFEPc3
uSXWSgzE30+Cfl/jyyQDvkfgAS7ZQDIo83xk7smNmAIeee2+/DaELACEt5jZ
K3l/FG0NiY3+x8RjdTLwUH4gw358fYAiRkyHRKlFdN7daXp+4Sz5RJxNuxng
AW+uOpQMi40esis3zf2wHwapgmNFJ4I1ncBx8/MNAcREoe4S3gvf6F1LRg3I
VOsDD+px4IxnFUbbQNCXqpGG3rGVfDrdPyTynnEIhbBaex5bvaKWJA9C5Q2t
4Re3UBWXJcLFO+7QdxlQ9lt6vXI52QZHv67I9lN/1177vPfWAYoWwrTrk1Zx
4+Uz1CWAKwqredHNzyHNuarHXZYAD4qnqod1p/70LVsU/Mzd8OmLv+XhlkTX
zc7YvpvONkLrOq/OfnJxbWPf+L/2INdTKuCWR93JOcvUL0DEuvrckRz1myTh
XdtXzkU73hf28E2eFQu9oE9s41Rh8tZdhq+/GUeiishz0AIdQRFScqI9vOBM
3A3No0j9PDvPfsIJAhk3/UjtzGWnK7gqa4Jeo8w5f7bmrPCvaj/BW5j1HZ+X
v2K2y/EBbT5F+av5CLVwwffanMNJ+qqHF9+sWoVdG2UwMpE9qNO62bmzJHNo
1XYLetn/wcVSUpXqxyYmHO99YAxDyoZmxehFUwyzW3V1noGIapxpgZ6hijrx
ReAfbYbtNZGX6apw3i6dwq/DSWvZ8T/0nPZiABSzXqK1CCja+AoYqVNT8f40
dQ3uehttnq+vEwlXdvyXQ+NCePV0WOwh4GiBiqznSMsKvkTQUTK5MpTEhnFY
MTxhzMyCNimYAQ+cvt9BY11SL9F3ZJ6R54fZk0GQQstIwQaTuHFAYw2Bu+9K
CdCYt9bPRnqYbo/9yhRK1gUBSGFKDxB6UalZwxK5pJmGOP0xMpcU3SZv1Zqc
b9D9ZLGYj/M0WtO5HG8UQTLuQeWpYnE9icawq2C1PzoWPndm8sqwadj5lgrn
qiPOO/GOmqptnYwIoFiMbiXmzLfY4qK60k8u7uCejdSyUPib9BKUH3P0/5g0
2ALZQEpttk9KvEG0QCbJhyB8ISYAQIJagvjz7sZ4C/HZ/JyTw1rhjz7fJyve
iGRAC4MR6NOOehYJtOU6hq+CDaFEthRyajivWAX3v0hPhHg+T23vtwVteRYK
U74M7BTwJfSqHnHa0QFK7ZjKZWui52yKAHCEoZE7fuAwWRea8KWUeBBswKf8
Mhy4kKK5zoffzoQslvgxsbFw1ahhrjndBuWHi33nT8pvOTT0FTezwKSdbwUx
0EFwWgKRHb79qspRT7e5H8MvY36ctBPlsVJT2K7StwYVOlrd0lspNrx0ADQe
MkqQMeRxob49ODR70uWoQFMsCw8qo7n9jCDoo/M+7z91Y0paP25epFLHKoz4
x4E+JLgPKj2qwmUZ3i+EQrvbJC/PYVklg/eZZk9ZUynO2Gxc71y58D9FlqyC
bXg+7/mv6gPD721rwvRzc+0osFlAzU4GHn2eVmHyUDEFKoFMaXAw4988GsQV
eRf3KXgax6FOS5xU2YtLzxkMVdDdDMspXT0Jtsv6qMC+f+lhBeXiZW+bmUHC
F+b+SN72+LUXLldilQ9wxdc3jDNHk2Wd1QvFary/8le47osO0ZfYzsCrdZmY
NCYk95vQ3KokIe62AHqsVvaiFohahR7E294GltQlm0WCvSxaJ4/vKP7/hqhK
PR3x9gquLk6Fv2oqLKjGfbDRXouBIfuOs/YT6VFjfFzLsbjESo48tfpxQ2GX
+Pe3FJguz37PsjuwpnC6j441rtWacN/QablCBMJvjP7nVcSKsw5MP48WpNup
ihiDoMILIt/j1b7b1zc5cEdQPDIjO1GdYJwDTELaJX/Qfgqqkh+MEjCHwdcV
chIS9ZqzSzEk3YLLHNcJNpqEVtmyeWCD9TIptvJBWdumhs7lLpXZNOOKP2Sa
+R8mdjYZyowZCLv1n6W4r9Re1KquBzQT9f8Xm2Ja05xkHi7XuayRPmfrFghp
8cBUtxDtOo8JV6Do3PxwoFY+q7XhLZX5Loy1LHVlel3zrJClxpqMV6y6vusd
J5HLNjxhK0eZ4Vfw6254satevhpFkSU0avuixMeG9Z3t6VDaYq0Lu1SunD7B
ru0NXsew31kLehDJcqn3nX8vaud/ctgr0hnMM5mCpbHq7gmEaeob7SNWTQFL
gyUTIwrhcXO54Jwy5SFYW7EyjZZiZHWE2oF/CLG1U8RObgsWt1Yraxx0FxGL
jWZ9GS3Bzed8YMQ9CpYIu1NTs6EyHT5MN0LSnEnQdaSB5dP75i5BHA7Cvv1+
BFoIrEz+20IJ+HI14WxADFoFteN1YN9i2O92C7YTmn0CxgOp8FhmMuN/CNmH
+OLja7mjx3zA3vE89Og2NOY+/aS/8sfv+xtOywToGx6j7IoIdOqQP9ynYXwu
OozHne+HSziqhSuqXhC6/Y1kWVyfel6uN0vUbywOfBohCiHeGpBFRQ/piNup
fctjTEp5/9AFXkIyBnC3KkER8EFIH4LZKMyMG/Ar6hgk6iFRsKKDAZ0/LfCa
FBJOl1zwPX6Yxic13rgx3nJwdN6gOKaJdpnN+RjmuMers152LUowJYIqXSD+
6kYT5PBpcqjK/A32ESTQK9iGJy3B4eiaECaza5Cu+8lfF+Q+UHD+YYGDG6eV
4WhTtOSKxp7H/3X8VKEjD844HxlEPpkvrec0mOdJjE0iE4+I863fkZdrIZlm
cDYBWLSUPaP32vKFYpEgH9/i5xU335qjRU7Ojbip+NjpyfD8Y/oWpi83EkTm
dC4rz9NWUa9CkXGkI64AyKszBVbDJ490Z+awNCUk0CK5Bp1mWhpib33SbkAO
ZzcZ58qHHBg6TuPg3iiNe9of0fkC16ojr7EIZscP8JguHEjpkNntjRfjqC6V
e4JgjMiWqe3jhAcKLUsSHkYf88F+cHJC/LzWuCnv9OW047+IL3bRQZuPVxLv
L5hapUKzptqB9Vp39aO1DERyiOsGXeA5JVIfOSa2uwAH6MNZISzf3XzrLaER
la87La5+fo0ioj6LCd1/XfQn1eETWNmCNB+ZOiVae1ggXx2GqivNkqrEOCc4
CyHBgawSAgNyu1AI4LBmmKCBRIGYmlHq3zFxaRrBJKiL209HkY/OUoh9dmWy
0bWY+RKvykw+JbjRgkAQGcECjnOO9NMb5TdMM+ZTbYMvT1cO3oFtuwoCv+M+
5sjIV9IEQEX+sWCic5+rnkFcGBckATkmFZOjKNP/JhK0WX8UBIxDAfmddjiQ
3EpVN4qIwn4QEBKRx2NYIgQaYpJQt5JPvTNMGM7HZplJgoZsUxcIsw8gHtTb
nNfkOwnRkz1bgXhEIsbTPO2JLoh1K7hR3ZSu/jmnwKLFPZiczSLPwZaw9Hl4
KYZT7hb9bGE4EFphqXDVuNgKgSSpcdXZDZfaoLz+/mei08ENDiypbsSthKja
8ktYoag7B0e/rV74PKOJYiMnbW+9P1LLeWCaSHFbps+98w1JtAWbkV0dpFbn
lx2aUXbBeJX8DM1pGKIroetsmZ5RZ8wT7ZLe8RfSmPfov9Kx+nPIsKU9Uyh5
fNkkmclWPVJGmP+mmklTzyfqSSCuNfNBFAkP3LHKLIUjkuLD3acEqnir02s9
5VaGvg8Er0AAGSY6xhxB6WtKcKNk3gHwCysz7GAnNWZREs/14mawSB3LMtmx
6antkdJCBbC31//7MpHSp8hSjsqINLJyv5FVC7u0HdpAYKNrjBm5rbZMi/u9
XkRT5uuif9eIgE0aM73pG5ie47pi2IpZpxDR/V9bkrAQHYyuHsGAgo5AjAd6
Jy4MwUxmWkypHwR8s+iHBY94X7FIgYTUjXLeLu22qy5v0AqlH3ZgsRW5Q/uG
gIvRAipVs7zEkMTQwau9NQoVZW0RzvtIsudlhE/1LnfHkfbgtlRUvoORfXxd
bq8pbGeg/mqttMM28QerwZzV88TGHPZigpFZCoQsbuD8alw4NjuTc6QKAzMd
i15Uk1gbGQ1iPrxgEY6klx3IwfFfO+7i/yYfWY4MBG2lbR6qJbvHyy+ILYkU
+Q3pJlDGLUI7l4siE7peCVMSleuysqoxIejkfclAy4/GYg5Qeu92X1G/lc1f
5QMx695itwU4jxQiu2drQGGK0Fl4D8IDsuukdWVDGrjfE+g/yOH2aoqFZ9Rn
G73qloAaxoJtDdCCMX8+C9N0pwVIbCYJWvHVdjlbG8nQKOfP0JNaAufoTL61
ctoiRHJBGHcnAywX1RYdM35OeOj5uTpPye53oj24yt4n0/z06lGPD6eo+oTd
5EF2nIMTUmK3IJU8IwzmIWkp4qsBuGF+7FnN6ygcZmynSDzSTRcACeRv5TP/
/CcQxhJ3aXfL8ZPPWU6Q1GUwShoNYCHnCimzci7KOIL2u/hGFWoXZ0WVmRo4
0eL7r2NwORA8YI09pOAB0RYLai0L97hp2BuYvzeaArwU8QhFUXW77Ao87TS6
Yht3JKPZvcHBrXvwpXJ+5202D6l8mjjxjJvYg1pldTjQbHLp1krFDHPef9hR
LX9aeC1HQF2IQu5YPxi3CagPXAwU4USgifMupb4uwQmaEMATYg8P4kfiS33m
VmLOpABX9CAy4MKaRt87Cjx5Hnz/HCowqyANVEmugyTz2Eey0FCGwbB4H/wP
9NGIP0Drbgnmb4+12vXSY5v66JvGBSRJfBPgUob7q/uy/MbVLPJIbji/jrrr
1TNtX0Cln/eeOUBkXXudIqOclXFDnp7bR+Q1oQfaR0ol8qegfgc/gohaa6KV
23nEcuJTrf3xjeCOSDlAiMD+MTvZx/lsjCJqVGaf4yLbYDHPFyhw9HLwTuyv
qP7NTu50BzEmNDqTTuZpzwY1lpaKwvM5U3jS8TH0CH2PQP2ML1v8EszExF+z
cwlM3vbimSFn/k+Disol6/xZrR4UoswUC49tzXAQhCcCIwHRprtZieP2UL+4
PJVY1Fgw42gVigHxI5cKKuX2CpETIJW/3/bWetEe2xYSNf/3W920GwZWtOiA
Ko2auPlFbz0kvWu6A6Lr/QXeg2u0AG+Z1xVPZvJMvGD8x0B3E1PRuWJwcGQR
JXDtN+trncaYUlRDjp7aum6ZbO2MBF+sVYOzXKT2zZ0Be2kmGfg/JXvIsabE
okILx15MHhYhCJMG1dfkYfRHvigcFewxxKci65GySbAdLHrZs88YPQYUdZW7
XJlaO0sK9opMZU8fZnmnSg/Hcgv7RmC1ppyk9SlktB4I5n1pvvkEvi7LE8bn
pLqDF+wEfX4WRZBOgKYTJ1rJqM92dLv+w/7rRhPpn2s0LSl09VJ8TjgzWPOw
r+QD5SXZZyx++aFLD7aH6TZEe+Kes/xrI6tJgxheADnyGvdR4CNlbESt5D8E
Df5vnxeVGQNP0BmVsnLji6w4MbmG56uDTA92w7BO0hqdFFcgbOaj7K2f75ye
f2QoF3i1lysIL/h8xrS1uWmGztjWrWwyQmdtEMa8sF5ylEodJrlt7u+ok9l4
p+QBySMw+I+mS8U9Xcc3IR7iyiIqgXg4dblyCiFWHbJtYtUC6pIk9ltM/UuK
9bnZBAM8woi7x0yPGshGFYVYpEkyIBlm3WSmr2AQHPbIE8WUKZYK21MHrlli
73C4aD5w02pHSnvi00ZjT7SXVVTP3P3WGz8W4oifxxCi6OvQcWnONiu/Uxin
aYfxAyWAjKT6qZCt+EREyJe8GBoVHFWk84GRwyVOlSXuwb0HD5mlvi59OfGa
koVnVmDy2LOQ2f4wp/OG9QFL8lNiYkMT0mnD1QvXP7seug8w6gIHqV2XrGvA
MMcPDZ1Mf5aJKf4oHNgmo6kAFNkFc9U+dq5Ylhyrdf2DRilpWLcy8rc3d2Du
GAV+jDcazjAnTtbJBMCuoOYxgNKwpk16Bjts4kVdlnFZBrZ+FG9f4eYVR2S1
bXSvnGGY+7eRHffzqQTvGD6m9Y7E8aQxf/T8c1DHg+jxisBlu0JT9x5LV77G
1whZBCrkuF4tf8Vp9BdLp47PPAPmW1TkVoClzA2Or6RMzOS+Eh/yeHpSSB7w
KauJeQKdSW0eqhoy4B/WfvI8BFs5FJrULwp1iQdtSAomPD3SuS4j44IbPdDT
+EP2vMTMXppsMavKELnF4Y+J5PA3H2sgxoXRq0rbjg1a+NFm/XprDtILIz/p
GI2yQxkDXqQJuTyeZWwJtClwpKWu07TnfhOPJ+5lIvl53/fGD+aHX0Y9eMlZ
D5M0N2zmJd2eMLPHIzx8zrk+nBLPkC2hOxOBSKHYkCQcToaQ2j14Faqxkt4G
1OeaxLaGpGYxBfSa8VCORbO6Xo54atZm7xZYxUTj7m+LWYpKQ25QAp12iu9b
weVoLvlsSsnZjeLnhtc5GVg3esBA7tWdeVd0+KSOdTQMJefueHvNkPOlHOXD
3x0cYNgYSRs7UzmZWMHJMpM6bFJ8QGs1OOzZhHA3jlGcKL2wMyzQ7tb+D7c8
zmnWJnyl0EDrbln4qcAt+QBeQHQ6wJC+eYnB7r+AzRooUkVoSWl7YwMx2YKp
REKMklV+OtDzJB2QI/TDHJci/UKzNNHhc/443GoojgUMPHV1+Rl58mcihgKr
6nkBQSNbpAhWBOCp0KGAMR1OYhEfRKtf9un/82+0CLs0/uek5VIUcQFSigyE
342fdMXw+TO2OPJIlgOAUhoKDIQTxbw6erClf/d/MnPGZ31b+fifkU232G1i
jfmPEGTSPdnkPEvcMRSE/oisoF4gN5mUG30kDrSg0Ox9/nLxoDASP27LFi/H
NvFB5pFhRi6Vs99+KO5fJdHpg6OBGlVekmrrHDGoFuXm7NomFBABoBec+/tA
owsmAg1JGh5Rns59JULqxmlcCHMtDhMyHtClGt3K0oO4IdFh0DYgmk5ZjeIC
3gZ4o4RrnI8cHhNLrJXm2hdTLGzKliEwe043F1pD59e6kyAp/h3z5a76ur7p
T+a+KRyPG1EV9rAL24rmmSPJvkO2iQsptP/LOaNX3V8kk40keoAy7US+iE4F
1O7G39XUS9IlnHnnFo1XjZvteErYAoV/JYXZiIwXSh10SFEfasjP75o6ukE8
PO3Y/a7dR8rR1A3SpIic2K67fUBMMn2T+oXZiHAA7c3eip4lPtRQDtov3YVc
hXw2psRND2WpnJpA17RsvPYtrOrVZiOLoo9TXY1Hpop7t1a1KTQHqFBYUQTx
cd1TwH3MOH1CeR7nmHqCu2OA7CLmi8nF3s64dlSeVGAmQxEh3Zwf1dXPPnPG
E/fFYgJw0W3cMDbTAZJkNTJDiamcL5gJLHjKnWEOC54b3neSY+m9qMmmzDW9
IpltpmyB63UJDMIksvaHE9DWWzNbLtZ96zwevOs/Hgmbi2xDNIDIGJ9Ybd3J
w1Kbq+IYAfoCsc/qme7UU9MaQFTi4NRmKnGyLGsZT8KUZvN91drtUmD3JvrK
UJA9Usm4qk9xtJyCAcHgLvL2dwIYZeYjw3MrlM7vSG+vfxHzCO49XgSLM1qr
v2NRK5qG9Nw1WSIHuCiHhUlxw+mubZlh3zWNkfK/ypD6rvP/y8HzoSG96Ad5
qt2UvH22SkD0xH2zzZCe0GsqEE4MmasLE5x5TSKgPCrCvvOaYdsjE3Kcl8pe
q2VjFKGba+NtILzLbpCeKfi5dnOgnKXpz8ei1NFq2dFp4fBqgXPOVPXVYxRw
ZVgspUfdrurd4PDLZzlWyes+7dlDVy6/w8mFNZ9efTtgZr2nob0Aa0wIWCH3
vdL0NKtxDFIzfMhn+i8cC8WNSlncut9fP3MIBkjy3UJzC7I14PrPDlu8wlP5
gVxYGzr9XrIovgHctjil/ansQzvlEC8EiRocZPnPp+wKHMaP9rte8f/J1b2C
CGpmilld8mpSm/Va4cIiQWdFKN9kuaYbEWZkXspjrbRbYFFIHTaXtbi/3UOv
+m6hyE/3M4KiGTPKv1WZcNfgYGbNdpPfcqPj9FouhoLvx0ZBIbo0bP2um5tu
g0dZW5vaPyUS0vG6wL78fiSszCRKKKKu0QESR26YENK0nuCuync4y6fb1OYj
97Md9EB8dQe1PvTkYO4iv7w5JIwqrf14wb+YxTB+2i3Yj58k4ALduZRH/OXt
CUZOweqWlPfKQjx0JZj9xHPYIfmXOUA98OQtGS90SRlqTiCmBnUE9Vji+D3+
cMdK4w9LsKoJhYnBNuzANw7ZcKwYcPKfrSh+QZSz6UybliU+LexYvSvxFKZt
ui30RkTGe3IuQA0uu2PSX0gC1MQ9V1klolox9upyIexvEOHJBo7cA0wGdiOh
eNTqi1CZsqgXdAX/ndtk7TVBPIA7FHt426m+3px/u752rBrZBstY7kMIddKY
MKtJwDj3+wroc/VTds0xh7cL4wB0r2eNrmGJUTt7ZODis/PfDrch59Oq5bnG
Qf7zGKBdDTLG/01GUU2eLFaCIij/N/l6RUMWAriqcSN3K0KtowpfKlviPt0e
Ib5HJNxW1h7SJLxOB5T/kYZhiIR29w2j+4hQBlvlAtKIDsAgQ9Ipdsf4RmGY
ZD8XgYHoLXLJs6Z4gZe1ANjsSqmk4DhHUSwmnaSXFna80vnYAoNNRJcxOW5Z
VERP/FXeqag/wYga69uv+tV3CJ9AevJ5nitnYkTWxGY7fGbROiP1Xe1cc6Wk
dr3qM9Nh3qIwh5qOyp+O8KkqDSBJ5MERTtuL3yUNIS/sV7YUk0QGNwcoqFpd
OTMQ1cd6kWd9jhd7rPo9Dkb/kt3WLGb6grzz9pJtj1nnRM+2NW9UxTX0Ofjr
4kI1o8prACH/JRRAqZxJzz386pwfn/o5XGiI01wk/8rJFVS+FVYAAru/AcyS
CCDtCORcqEASPubsFr+1EpoJxSlwrmZ/64WF9/PyJSlItpAIC7oxEQNKA6Io
VjHHYME8qusFJ/JYfpGruYf9p6mN4TjDffxAAYaB4P8XDIWcVbKYhE/cFXO1
9yKaunVCjqtOdECtSbB6vICxwbcUNMOhhNWgMJ16z/Gfiu+sVZ7aAXCjcQYy
9ZS+sgYCpwx/PR6tfmINRCU+gTQCO41IDBH0U9ckaJj187syqLLGfw5JTUCp
RBaMAml7HUzqvZezL8BHbbxi9Yft2OaO4azJqri7Q7hv8e+TWVynnuT22WxP
+9WTWY+8c9gVelK+YJV84vdLEAhJzk4Gagq+n8wPfnX6sQa5g6o/XdhHbePo
tc3ZiA5rHmybRntOw0kGavNey/sdEUzOx+oPxS9igj161VY8nMG6gSCA7L+O
C1bdd3Vtlgu9NTa3Ed8BNSj7zme6snx7t3PlG2iapXqf4TzLVyn0lLs3QYdy
/yLuHEdjx1vcNtd1bAUDwQNAgznYgt4hOGt5O7i3YKuenmkVdqXTmVZnNCx5
986yt2copQe+lMYm1vOPllg8/WCBxrvKTUP05dWwN55ov/foTjNqXOE+5InX
Pka9e4SWUnrBWXNuOWd+0entcvjg20Bf/KvIyQvQhcTDuBKHZuLsrv4cpdhp
DFTKZ0IiHT1GY3Hhw8pb1gwK5gNCKzGa63P1osSxqWMZc6EoAPZmxhxdzRP9
mIlDUjNiKImkr9nFuZu8hTDOz5XqmJBddQ5tLR8uPjSaWOkAXPD1ewf+FO0c
T2NLjRE4/T0Pa+PhC6dfQCUrA/6Hq+TyfHqivAndbyM5o/QasfGkaEsSz3fp
NK+RIByLR+XUmxzAK1uB6XTlzHNGPI1Uhd134HpvLInH45Ij1jCTMrwo82bC
nLJAkEwQi3OmAjDXVda6hYxbVTSZ92CHoW8M98CVOy9xa7FEaOSN+MJr0/S9
D7Qr+1UJ9S0KvxPYXze05zEemEDnrePJJ8EUVY6p5XAFFq946Rwj9CaXeToe
C3HN1tIMwSmzvTi44+DUrTyjIOkCvF25u3ggvtdSgnr7+LruoG59a508Bi3s
czbRBZfJSnAnGSkfUXNYsbuuyTwp36RKtVFVt6WCE+5vB0GBS28AiUnWfOuz
mTcsSgVtE54DOuU6sLrljko/4UsOV49SYPVCbZCEdG0nK8ysZihe3HXjaA23
pyvB1FW5P9WCAoPJ2ZHnOvrgJ482x64uF/doDAnXsBDDuBvVUZxVfnlFUzXr
KJVz/tMMjUziqR/PYOsKjSqWVo/tEHZ6MXlSMEIBK9IKKIRaNHmyqqCaj3L4
aL5ROt0BKfY800MQYyAEbo3R9aZBmE+gCq2d9KuaFqIdJ6/QtYSMVGtoBl1h
cGcbr4xuh10SS2bLoQ4VAmaHS7AWfGQfcZd+/6+fY/+kndCv5tsEIV+0H4+V
g4sXzTQv0OerqsO41mEUjJnd6i5RoNcA7+p/3CqpSvIbv5hOe4CXcHGF+EIE
mV61JzZWfmbK0Z34kz5sGmwOiDI/eKoGk/F97UuI1CiX8+ruIGHZ7oC5RK/f
31GkRB1hNlzamujNXfNWK6/FSqt6HONb/eXrr61wJSpEa9u08fmMQTAuwx0/
diclP7LDgwwfRwMXuSdTjL9T8pkz8fzHBsLGl306k1TZk39z98WySeHLMP4C
tEjQ6koMTzcd7vb+G3z0TsEZwFx7bE3EdS8Mqk3B8Jh2emges++HNs4zOZ+C
AnzwhKgByzQgRjhFccaTCgg8577mAYRjyg+/DTTfzFPYZHncgvDSlVArxyyN
n1xu9VZ9ZaA9SiBsu7H1ZOk1Ids3J3jLmPVhLcOCR8ncBbWBiH7C2kXQCT2G
Ztm9dZcrslQrEJb79RFk7fJLVFbEGor79geOXmt/Rxi16tHzcAY4vbRooFy4
HzP3+nEaMDMEnHZuOaLVaXepWT/9nNlf34mJ7P41nppLh/2W+8ilhynvafbX
ENpMo+tjO1VZDaFxtZuOuFUZK7w4QBxNEg4vZl+EWDBY2LtMqKZOmAvpZwyV
SbQPcL9jSJF6hFgUmtLCfHpjCmK0o568SUpbY184ZvTY4cW1gQQpnzCobsxq
6G/eAe9WaRPnb0fjVcJh9/kvLPAs/Te72Zb3EXUdbOGHw29zMfRBFtO6QbwS
YsSZHjhXr68KNSJZwbNEezmU5CjoGl+KBiWAfCxgdVG70jGAx1ggDc2B7Gp2
D2/YByHxOWSIFo43qAB8+KRiD3tjzdckc6w8F55myTwJuCC/nQw7Txtf75ia
+aJag/9mlptC+z58oVn9GrocpcJ7+SL64t6leXGUUK88ZWNEdHpGo+32C2oq
BRl2Xlf5FrogXyvsDgOz444DxXOBNFyZpbSyOX6Ii/qaOwBH6TWdAI4MIbxm
ejt9jsxUBg9j7ShxCM0zciNWGXd3c8ccHTuxXR0ZXEOgYh8OsnLCRqhzlE61
qNm5Ur1gXoFbHHsJJ43wtBtrg3q2fvehjxZtIJVtZI16vRq2x1Cx2VwmZSib
qvcyGbvliQG1nlq4jol0CqTJBhK2OKn/UpvJu8WgoJot8sXoLifsYvtIEM9M
q9V3Y604sWCx0ypm2KeftB5DHkYmTnXTc6twDW+1LX0uoR2UX/jiQ38YA4rC
HKJrTxpVXRkuKisRnbRTuWlLsuglWcyoXK4zwuEiM8AnkONMFMAok6Gox55g
41tiZAqtsgykKeo2eDPx7SfTDhq3xnEwgkJYggCgztGDNbif+l4CBVTe/834
gCDB49WoLdd8wou/kmD+Y+EXJjbPJOkh+lF92sNt/VLENUf7YvNnG2jcwmTX
ykFeYODCtFOe+1U60339vbBq5EJ+K0E7o4kXPjrKdC7E7XpZKQ2EBrvQTZdJ
RW1MjhW2kkLuqXXBi7SZZtMAC8k9pNCeieSc9DICeHZsaZNVgFCmm/GSTapp
xNruRwkYrK/reMmXkmkpixqZdhd9Wg5FoQLewMe4jRjskRmaX/WreUMyAfV+
4eFmay0+u0mRw6i6gHmAd+UKg+5Vn01+Pp7fPCkqi1gIMdJ0ccGXE4MfFeS+
ruuKhhnFJdnKOxGEK1uSdZMoPMhZMYVshGxeSJonkdvxpxIU1p7neRmXk9yk
5SwJGwmN0jagPgdgHuoPHi9fmGI6jeS6lCj44YtKpaDiBsGpqac4RG1CKEhS
oTO+Zkgv9+1462ckcmmm7/4rv2+1jzcERRehKmmNVVD+JyRecQgF83joPB3h
O+Cy9aQZc0qjrLODeRsirwqWBOuxbY1ypPx2YUgF526+3w9LpWWAx2lbPD5T
56msxV8cga8gIOxpU3maYe5JaFSXPb/g3XfZlkIoqWap5yu1ovozA2XCIcNm
afgsgpOrS3LQJlmd+tLHWEADdMAC6pk5PC+Dv0o9s8ITuyn6MlQ8OuKyndxL
CrIn7AsYtYiRUhrUyojCPklRxAoz+JqZXpcMbtLNtO+uCohKuesv0lakARXF
n2d6wrkZzCjX4Rs6KNhpLuCnRTYzdC15m8Sa45dayCCrfV1JNQc5jL1czgxu
1q6uAkLlzAKf4E+ItaLxnIcYA7JbmHi2jMMrlQ59b032OFBdA1w/Cm1mOLjy
Kk7rQrBTrRZWJ8jMdDO1dUaKEqG+DOXyHE8rXDMUo2ZE6DYk6mhL1uHKKwpw
AYslC8gpQpy8FlfHL4bYLrGggEGw0jJRyH+Ko2q8F2stciRkw1EQKVCQ94y5
AxAml9LGbN911je3Wz+X5YIC4ygxi27/zGGBs6kfSH6CPIqJ+qJnqVJlFIJs
mwj0KvQPeeiBt+4TioZdczyyUqgWM2vejPUYFG7crg1WKVVDDDC2tt9aEgNh
RpPJoSqRUmlJnW9ihVQ48xwdjPDVU1n5HxlcUFvjEMMH6EpBGZWw5UmvtFRl
Rasn5MgkcTbjq6FC/Lma90DzxJRJOzw6gvhpdBTu4iHMZmp7ZQ6e6MmT/vly
2JE0yl8S8wLHrrnlyYZBrIdGazeidWLmkr+RcCHwXD9epqb3+UqFNNYTuGCY
rOubCgNEmZeE9Zv7Pw3iOJXfR0mNEtzfBjNfQbPrzDCAmf43qPyNssRS89o3
2Xyq5WtcSPnxA9ocmmmEBVa3Oatmf2AMbH/uAfTcWVIf/R2QAlO2TIMYX99F
WTBh89dq0BUIj+Jp7D4c0a0GielPhvGoESHa+NwDjcNpK2GzLj16qxKwWjOH
YV5FU8/Kmba9NFSHfJt5HiXOoNJqT5ndqF9nPvwFI1Moqkcqajz3xl35OU3F
SyAtyXTKvk3KXO7JHL0dhKJ/NvC4Tr35EBOGrng4tMEyn6WMWxSKxVMSf5CZ
aUsKcvNpKq/xa4Y/e03fC7kV9byuuxG7mOTwTclbOyoOSMrBM+b2Y04XpT4l
hJ5Fqh+z22g9nxHwJsYnec9kKjaeyJlaTjczmlPWxnGT2p3XbMuVd83IO/u/
LoGYdB+GhFrEjsTXCx6hiaQKxHMk8Mi+1xPmFO2Cdi1KTFsNX0ZRH3UCsG8W
yiLI6n9hsLkBNZ9YLYm7QdMzdvCWZmk/cJOzzzuAgIYTPfD230lfFKHaQlB/
ZgfcGycvRyZLd9EpKJiQ498JzugsC46bx+fymHoN/GOdeMIjNkN8SLkwa+gn
diSDDAaO3K6MUZEJez0c8B5QbvKtyrL+Qyt+ydpnHFXMcf3JZ0elgGlDNplL
x8FmP2AKQw0MzvuA93c1R6u1k7kdHoRcJ2YXSWl4gCC0Yo6sLnI2AQ7tCifk
qQNJmnra8mn9IqO3XmRWkl8eJQB7F42+zml5g2AGQrnUS6nUEQKJ44Cj1lwD
Mbds32z4lzcjvsf82F1NS8UZmUqDzd4xDKdZ2vZFOfY1Moe+aQf5iIrAy3Pv
vC8c0KdJr0fjiZKQl9Z8PGvaLwJZ4a4asAFe7h2OpC1rKHgwpLgsjH8vuDjs
OAO1iI1B20Ma6R9SdjfN1gmxZD6gSLGYeKtT+CFuDGHRkjQAW76HWZAx93bT
Jeb5VKVorzhF2/ebEIkWcMTGIfB5640d1gKOmdboz+FmFnrV4c5W9w+1e+uK
WGA3v0eAjPzF2DZYoUYKfRzpUKxUR1T3vyixsG6zv0erYr5K7Hz49Gfg2mIo
Ls3A1dtuIWaCZwJdeCYzBncQQwwgwAyoWX9Y1C3p2HPePkJSPhOVkLFcRZnJ
0MzkOYpIWCKOqaOHuSsFge0IsxYIGFzFcC4M7tmoXBW21far9cRtrJj6v02g
v7XfLXX8UXGD9bfnqj2PalWWu4VJdHx3ePqhENhRAc7cQcI9ZMM+/qmK7ge/
zpscersyK7PpzaCKS74fPnm846FE13PxyRBBcSCo44x1PJnQaJzfNOh8XW0R
NNPieHjtBijqpNn/O/0wzA6ianaYNXQnzU0ufuPwISvfgSmApJGxTLSD3JvP
Y6TG4rKmcIBK+C/gdzCSawk1ZY8cEcTcpl6qgUWS7czZN1y/B+VOhhHWvo6i
XdxBbdR8+qzFVeMKPz+06a5YoGTIidiVOe0n150dBBzgNAWwMUNUTFCvT7tV
bAtS/HccPUsohuzGfU+EIDtAPFq/SFDx20BW72Wchx3GXz9x23iM48FAWujV
x0zrCVv2emBaEC3+nHqJhK/z9Sxr2xHVkVTdhRUSmeJCnU7hNfwzRzkz5bzr
OcnyFdQH1gyKNMEPgrxguKgqRXC0P/NWcg8RV7THkY3hK/LyqgQspV28Mr+i
adfa3eJBkl7b6b0qHgaYMtGKBYeptPMcHfDcs1ytuEn6swzWBH0IFXhqla7u
gsnry4o6FKEEkRA/sva1J3h3Bc3zq7LHBn0wKigdD7nox8ZJ4y/CaDZQe/o0
QOZOh4S2Wq4Nsr3SZtx8qyX3k1pqVoANYTVwxzkdhuacBTgukmUul4rn/9hb
7p1ywtbxarUrzdS4Jc5sI8GNYWd0ZCptInh9PoL/ByD4omf26GbBCKs4Hyys
ZMdsLHBPBgqdtGGygviR0hrFXoLEs/ohqg62Mj8Y8XJ4+XCmAoyGIDMFnX4R
jKCo8mf0NT7wDAQGOaSVaFyD0jWnp0xunUCD/mnFhBxcQ3Ym6IDde+AUU1bX
cRxa08Yc0HFMHTqXiihtPLrP/Ht1yx4I5f4wCsQ7my/X1k6+1DVf8SPFhnlz
OsUAxTxaTxMImLPM0U2XjLjAB9aX29CEm7qTZhnodUwCQIOcG1zjiCaRraxb
wCr3db6T6yHbMbzUrFf5PeQ8NbUpqcnj+eCG3GrKXX5p9BZyi62l+D/yM3jn
ZOJM5quNh2hzsNWT0s1vJe6hLEEuYQkTpgpEunTcpeUmDVu09WxUJVqYE25s
TUfm9Vuwpeeq5+uL7ANCzSlY+s7S5bRyG+rcgHYnIwfVx/UmRErVoLYg/hsO
FiGu9XI+hTyGaI8eU3sWN0s53KutTmE98Suz3FKETIhvuhO6vTvd+e1EMawT
kIkxiXQDCfyqabuuJZDosMn4A9+tj5m6ULZEvi5/WWkgax2WIeMTXi6SL8Bs
xAalXrHUk6ozGiFCmE5Y6N8mwgsoAS+LV2LhryVR5wDC2U4g0rDRgXqFihEJ
KKmgE2MX9/fpiVwAs6VvoLrNotiZo25ZfdlFGgIMUGgDismGbdlkaYooSBSQ
soNZ6lA4A4ATnH1geUTl+KbliH9fO8VGO2hxYv8wkF5e5jI1RLaqfxIr0UMO
V+iK83f1Aw9Mxr9xB8ngcQIaheIjMwWYxVbNiF996OMOyfGPuT25JLAoIqa5
pRdAI1pQDtnOvu6Lvrte6r0DgICC//UOacI9F/wcqi43wvLs2sxdmYKDjCIe
atinFMfgvLuZh9yxryLmpqYvL+Qv0G690H43D7CZlTr3ghkOSql9VbLcGM6y
SXRPJGrwhOgmhrnDX9kOEBiGeGXL5ytY/YTGa7kTmSvwQHhp8HqNrdXNnKB8
dNrLqJwIFtK8dW1l4YBMkQrf41dQhDCs0iSmCAzp327mlj1rVtQ2ri+4tsE5
ndePuQ1uz9PufguJIlDYLQM/eP9dJvkkd9++pFn36Y/LfKWKsxLHVzhmekBF
/RExGVsyk3kfBVIaY6MBlswJx7ORJbXvY1ACjAZYJLIrARv4lrKKy34oT3cC
Q/QRSUcJc6hsKW92qCjPrBSmg9MqFfE82cVmcJdtIQuwIfz2BF231NP6RBWI
vyCxtsBo+g2bWP8fCGkEoqn/oo81IoQbiWA+MUbZcPSii2UZVy2+eQqItJrL
eI3ye7k5CSXSZOukBgFwZ1RHRNtkZ5mAKEq4vxDp0h8sjwB4MTb+gQ3P8NSh
weeOKXFqthp7UZKTTnIDI7G5WMCz75xGKm0jSNokCxH9owIDBI45lP+xAbqQ
BFfEpX4z3AvRBdtyUrOcrRDy/oKP8Hf1eWjuX2XGWWk/5pPUak6xNI7tIAY+
pf58+QCd1fg8P3YCFh7weWYrThQw6NUgQuPJJPozwGSzhisjruUiq74wZIsI
m/nRchsm0ypjq2zApBi0fy7HHN/TTEMMbZkTXi9zfRmPD0yEFiFEfsm9eP9f
XEXqlkDP7ohJyT+1lzMpB/YYGY8CWRCFapDXBtQJgUUeSkaTVe5jEVfq878q
VOZnJJs1z4ZrmBqC5CzQ84XcHvb0XmplgpzGaXMDd5JkoRn0+BP/EnkgeQMa
PgtyfpdjNtYiZpiI9JX1gT+X63w4nyXZa/QJOh5usugMdsLaYIoBCA73v/dO
DfmdDZ8D4PfPP6E0FOM0/gFTqn4U6lF1+Q+9qqSHotPXuwHmDaThjz94rx4y
skHLvdWxDytT5Xm/UWgwIgJ7ei1qjpItAcNT8LM7r4zbMBBlEbK7M1zbdAp5
CURvWZJR6hLa5+evDQ7vs+Y6MUmKwtqeib+tUx5+Q09LJPMVE5mvHm6hWCfN
oQDRHmxW9NMZ2IuBpmzP4uyPuJjJtUFIU2tyZT/T/3eCH8Mib4HeOTGxdGPM
fpTt3p6TFSemUrVwMjQh60S9cp4aVT0mB7YBnuWknmwesBruR6f3eBUBLa7I
xGM6cTcaKW7Y5mWX3HBm0LKMiuLST54IVCeoXzD3jSCPpLZcCWNfw2P9Tlsy
gKqpBKEwP+9oc2DPT+bmaa7ymyYJ8X24LcAea0lW+STlNHoShIkSnig4bIFc
+M4NSFBACsbkCE0EJTYJlyLFa2hkjXOMmRshsc/NtAb/RiXke2OLmGCC8JAa
IOqhH1fzTTrjaQIEucqn5g5jOR2ETctUQpn1lMlDHLt7Q1Ilf5adEOiOu9Xr
0jvDLVftIicUuEzgV7HJuNlfv/KweNWupy2zb7IfogJRpoKjWTFcKx1Bdn4+
A52vs9l8rAFyuOrk5vKYdHrvkYMFGnA6LUDilUwfM6Qi/xcPLsWxZkX87BC4
5r5FJkBC5ExOE35PNUfkWaw4tUV2SjD1hEWeYVNXR44LU+DgvdYSBzWPdKuK
mVglbJ5OCWtHrXwEhzx8r+KNVu43wye9UMoGLSAS/BioYDtzWtlTZWuV+ku1
czUMQmN0ZyYaPy9l2aqwdlEfHrmJSJVnhVS0HV7EW8DoSKcsFtP8m59lLKv+
StHB5g74FgiNHec+gHxdB56aSaP+IrnWB0q1yhG4GouS5ZOUZ9znVCi0zSc9
It2G5nNpr52XDzjKJEhxdriY97ZUzFg7Tatu7nuaIZUQHVA4wMcC76dboMv/
qaPXRYqDcGNukx0M0wJt2mgmE6NB2J9VvOB+9NjRyh18SDnByAR8Y8405iyI
LYUd0e+QdyoapFzIQ6NtJzaqlWPyO6hRPq6pv/76a1oOSNYGYQbV4izi1gyW
466+kEuyIkO/uqr0VqF+9aSU7/0I+m04IzAcCd/Qcs9r99eKo+nrsse12nL5
kbggA5tJRJlpA++Y5BMVFasXlsVzPas03o2n8aw3UNyLd1Gu+ZLomlg/UlLD
rtUImYex2EZcfp5dWjGn62BEPyvve+9TnsQN4zG06kHbFHyJzZPUBmKzbDZf
gF9sbVfY24jvAC314dPH/weJv67W6eul+cbYoQrJg7SFocLDdLFJxBWxPVRC
KrKuQP5qa8lj6G9pLsIWQoq5vu+ffQec4OYLhrd6fF3XlIX6yYv/uq/cEiTe
knRo7Rr1yWMzqczE4oVN0mINv3wzp4Evw1sZewjGOAv/zOO3HupuHWUXbsZS
4Sq0UWo0YyPyLNG6EMogL048R97mCFXsLvS3Te/EQBDuZGk3NpI6SkCNkSpF
NMBmvB7vtbMABVxh5OmRRjte0EItZTxpDC3B5q+xqAZwXuPiSKwcl4YzZSQW
RAPqkrwjMD/8iTSMvzPigx+wGKomZPZuTTrQczGujleUS5k1cuWCF+8At64W
DmDDMDjBQ1/e03ladWfYoEVW3ufc8h8cI22i5NdByOJMc6a8/Iyjv6AZV6Lh
0LAMnaoKHWbCPUWfWULjresFiYra6W/WazCJKj7yWFlUyfN+jTu/QSMG/fEB
HPJenr2kN1PLOb55OmGjfUx/Yf+8brx7VcVa0vpDywjXXBVDyBRZw5XXVqny
nvKIAfYl6iZ/FReJkSxpzGvJCrYVkumlp9UPYnG19S4oiNVBqEBHmI482V8h
Osc4oc5F0FC9uz0qXz67Ji0DPlf9TgwoDUEjbI77f50a/bSt8lLlOlGnDq8G
OTa2RJVxBjloW9Y2W50Zi88ozJbxB3QWiJ+rT1/lpkaUDEuOKvsGNN9NO9nI
dChJGMDxA5i2exqoZNjbpJwYZUl8ZNxWcfG2l8c+0NPhCCg7g+5h1rshcBbS
1vy3Q70vLg1DapwxtPLiUrBQP/bQcnGbUvroPWX629dCb7DTLDIgCfU4pHii
Ca/TQlCNPvSOnO2ZhpePUOcaYjwLrIZdG5hWjFhDkzIRewTxr90ryQkZeqxy
Qex69nqQgYSiIOliu2ip8J8bdoFSFCGz1nmRc3mXrtzSNk1VffZi72zmqFZC
h5nQAzsJDYEW5P4+uAy1o3ePBIzmIbsELgerkBdcg9QWBMhpyyCVaeQ33t8I
X/x/Tq8pDShZzURPmATGU8vaKZ3a/cFH1576pYKxl6vJlbHWue5d/dbjzpiD
H8UYbWfAA0htxIUQTIzyIxBRXrPhh4bb044eWkv0CQDR9kEmjaKMD3B2f/oi
E6JBMhw6ipxImuiwBfc7MOkUErB4j+Q6axH4SkZjsuKdyz0JtHJpcalKiKd/
eMndblEDwZ968DPssF0i5UwTYQ1VVoatroZmeS8liLPk2HUSAO+UVerkfHkH
vedyOmBBjPlXFtxl3Oz2jQ4W9ZeHmdIPVRJGUHulvktLruB8DK6Bp8hJmJ39
U5oTW5uSRQon6F7Ty6tpI98WqWJUoiujtreZPeI5LgcwhoRauZjd2UIvAPvU
ADGaaA/Z9P8c43qZ1pxRDAZZCSJrcy6LhAL0iQYwBh1O0lAHNQ95gvW+dOwj
OK4yEupZWtD8sVK2wKZRuJNVUT4lGvecF5kHF/uk7WBzJxRAk9bb5ldMxZVK
2MimJK+IWxF3qFkz+ynevIPKRM2GJSBnDQQ+SE61/I5yu0jgvRqZvf4Tmoi4
qVpe470yx7DZueKE2HQGrw5IfawQsHQUeNtOGSdfis8mCmE8DueNlcVmMB8v
tzlwoJRjLk0+UCDi+knO8KX0CMyC3os083PXj/5QNu4YqRqvi77cp0viYUAf
BqIPBPazxsJQj1Dbczc65kctu/2U2zmVWVqwBycZzBd423vamXeHHM9cTd7b
ZT+iQj7VSXhJIqW+7jI+f8EfW3dDNf6ZUi89d1EnCAEUL0TsnnChdsMDxRmD
1FIcKPRjEupuX3l4lrLGN/12otNGwHy1c4Mdj1OBjFX+8XY6ggxbDJDHX9By
IL3DcEJUaopRysaqbYanSBx57wMSywv8AiurhEDxhieggZ4gQaCl2yyIWF0T
Sp7qc3gsXC1+9zbGZRraiI7htry1H4gUCfcJmt2F+eq+kxCTj7QVfFu6o8FJ
L08L4+Eyl1SifkEoq0WVfcMbmya99s3wLz0vwj7cj9ew2k2f65XEp3WQrqi4
o31SBQYewxnI91HsCJJeTvYC8AbftLPZ0LUVEPMGrzonL7lDhBWIPqxDl3Ac
bKdCKpZfUXzfLYyV5JTle9ZkVw/Ak/ChmsV6WJahAti7yvcGmtOCcSIOuee9
9fiCS3CTULSqRltPRaEb5A7VYSEp/iMbvvlFAsmEUGfDHJX7JV7ogabgHmax
ui1cux8aVsngj9sFASqYmc0UvOi0uN+lRMMDDM+xw0sS02XHIw/UwSq0uwIK
yigz0PiXanMk2lbMzJl8EZ+Pbxo10atJyfir7dJ9T4Feal0fyRSheGQ1/QLd
9XaxBsgbC2TCQIOerLKFk7CSo/fxmrPLfXxcI4Dq0mWo83HFspdsSUpkN8ej
S3q6TBJ/SgA9iUxaXlZ5UfP7pkPCJboOLNE7KROZfXBFIwTs2dtPrf6UBAyg
XM43sMedqOnAUcHyJ1HbBgBH3Mdt8b7/J0Bpzwrs67CQmI56AtYSKuCgl1B6
2iJmMFMReANslQr/QIFsB3f0TlxayD8qdtoW/DsddevYDIJqoqaMP+Lz3kZl
AkuKxGcUeg/koM58L43IQ2MLaqPwkHzL0ZjNOdQQVn+wknAjqQTexi/OwH1r
LZCxG0lG5/fiBTHvASc/y6BlK6VyAj3fVtTU7Yi1QVkSzZiynFYXw8Na+NqJ
nQ23nht4aggzcFySTdBEvrVLkWD6vjpRt3MS4P10QDJ8tNpHWP1RIV4gedJq
dKYh2Y222uYZsiz44Tqiefp6fGdZucYIcaopGt0TnVwUNYsSdzRmCwXmVZup
bQ9uIXyxgIwLPPt0xHBJWouTWkJqxrPHeg1NaopK6QFhedcZTrqJ1WSRfVPq
YGiicOl76lv925yoca/w/fD3sld1a7Ji+lYtKwvod4YfuqXidodbvTZt5rMZ
Lc1yw0EXSrIwn0iIGXNnEA0db5r/EH9NYeScX3JqrvcVYdTyqG3cW6+aE0Fr
/EtHPXTmneWEqfZ/75WRzNO4Qx6TE0z6xOoO53960g+YJrOrQRjl2/fwe4l1
IL2coEfn7/BkjQdDQPrX8RzoahIyzysXwrOYeaAQ0YTVjEE7rls71Kh3uO0y
gJyeBiC4CUjS2FfGIO04VNehbfV8NA5PJ2fbcJ+3fXw6GRkpb3QBGcOLyXnz
HmIXUmsJNttOSR0y/GYFzFabS6MGtEGmq/qvntYu3t7VVyVgPpUAqPoqMyru
NfEUzfXdoBj0j5fV23/C1nojQUxmans3BvmW2jN7xmdHeyOVUlx27Ax1zyaJ
xdkixzHtfrE9LwxtHfnJ9ICa8TzRukpjrs/B3reQud6lfg34lxDrZe1lXGjQ
i+ELzd79ACbNyOhmPuQxtG4xtxam7gcj14n6XNWzQRTkvnSblyRohVCUWF0Z
Eyu/8Rmf1KFBLX7bYxpBqIEBkGGCO2PmBIg+aSEPHmetFGj9Fk3Oisew+8n+
QykaMF8REkzHZJRTFnHkV0pfits2IpRqWeIIjA1dlAhirK/zOXMV0lcU3yO6
oP91hTKXs+M6fd48Id35RD4h3HAp3OJVpyf3EvtjKJKHXKoMzI5O1QAmo3Br
+6hJfXN1utb49dzsKjuCh42pdlu17lGHAC0RFAv22Pk4Wk8L/IiINa+npdbg
C1jm4pdN7RAJoCPG+sqwNzd7ZTU90zODjugScfUKFSVx3c1zAMTGrYzrYUFV
rVRQf9jwX9cxp9cP3TbHI0UlnV012TNi2vIdPjng6CLtf2LfLeXjdm0zOb2h
QJ3VAZoPGaJF9rkzsPPcg6qWiXpjd2BD5CxObagRhogWCfZcd5TguCzPyGBj
kKDtSVC6m4vkHO524ixge6aW1CEBSY12MgCIe+X2kyaMYp3WbfMiWhb/iCzz
bUjZ8znCmkmK2+MfFNpna+eG82cyqnuPk92JM5wElS+rnytV3E8bEb0G66FK
79qaz+OghaTmahgKr1Xa8iCJainaYvu73gEN2UO2de01BHjLSbyrP6gHvnve
HwTQgM78ojD6pnXAZX9Usm/awDT0W2RM4YqKGMhkPvzoV7z2R8rUoOOiLcjU
Lzg2OTnbPAzfhF179v9tzFU/9uecBQcNb5j54FcoTewl552wgAQAt7BWnHP7
ZdpTZHrMBpp+9++PRAOS1V4bY6LM20yDsiQYh13nogW5+tW+n5K/VFki2KXp
cR4uYJVc08j+qMuUeO00aeOycwimOuSwH9bWfj+WDcrQQvGGDo6nMKxKnCVt
uVxD5NNjWhDk5Dbd2iUnSCM3i8VqyMqUPoJJw6LyECLJaGnQv+NTTpk5kCaG
FIV0wgy8STMDm5KhDCgTygdG9A3T7JnVIJdfQOwyaUbmszKUInp49yCzh4j2
h2+h9AbStce3Tghpb5yT0YAlBYI522E8fMsofSKF7KBGMQrGfzdi5WkANh6R
sqQrJuWXvgGgyKUiA69pPkm18dzIl/7coWY12StSbFnBa8ab6NjnrS63W4tR
Q1CAikwLWP8ApZcY+gkRvUM3DDRcfBSVUeIK1FDjibnFP/ehDK1vYZVuZcsn
wRy54a1+pho0ewCRxtIhf2FONdA34M3Cmxu78YZeF6AYevU6uLpx1bXn2Ftm
R1T8I1lMtphkhqUPp7jNW5nABmk0u0haIZHC2muIrtvR+WXTNqKw64Fj/Ccl
5z4nb8uv8E0poDOpFpokRdZup/WBaaBTX9y3Xz1ccLMfdzY0vNJ0X4F//FRE
n4m5EXDce697SQB4/En8JXAPOwNabrb4Moc3IIufsJT2q2io5dQtJqfIxpNG
q2TI4qFSLjERPjydH4iwCNNMUCcO9uIyuVbcWOsXpDpXu95zXKlWREntITnX
2glMs21f9r5btNYxbWHZVi9n8T2LYqdTM18SbNAX/lFoEdIe/n7+T6pWqiRa
NkGZozRaMitv0Xw+TN76Nhg1XV9LDOW2vjhRFrg841huhwtL7RnqjI8Q9CVQ
KwkfGSkL5ETawByjl62HgeJa3JAYOpXnj2PtNsWoySVfpfq/Q74tEWMAoyOc
O2UYvqmhSo9qgC7IMOvYVZss8BNuQDUaW5Nwh98TPINwbjmAWPy+k55h1uDP
nNfKjhPhJdGiykVugga5aG6+Cxtb77Rg2e/MPzLrWNcmopd46+iIg9LQyfEm
i5Xrd2jDPwVMc0h/lvybqVj6gKpQyeKbeQDftV7m3tymx34G6WcdLstODSpz
bJcw+ctWP/TuSvrWzU8KS21jgNj2yaXZDQahYdJlA8/sDvXHaezsy0e6uUcN
9T7JlN+3yaNW45ekwchDM/4zqSdbRTw8fmyq1CL09R9c8O4bsH6+FVomFVdv
kLyv/e+LteDb3Ce7XA5kuTOBEwfbG7Z0Px09c5D1DNT3SXIgI2UPMMctbkS5
QgADMbfnbZghD2y2ADCi8G6+VM6gCdM+T0rm3ZxcXeRYqKJ151ZsW9Kk8k3f
GQRbz8usrtmh3cwyZtkIV8qeiFBTVKVqFMDM1vKpBvHSKZVAqWIzKVJ7tOsU
q4mXFfmPe7FVUJ4KLvob46AEBKLt0ZWuECQpNGNN6U+4/mT2+hdWoyVIMUWl
oy77MDd60ZmrwoGGD31M/CgpB2j+9b63vAxZvsaKoCtsqdhtRDndlrGX6CLu
lnLifLYLPS+12ZaT34kf+f4ShbgpuAyMqPZX28+odPB7MucGGPel50Aq1fRy
Br6Tigt8ihRvBF5udUnJaPJq7o5dMgk5Fff5fA5omGhd9rtFhBaYhNbUGr8K
Kv6W4YRqHQSmM9l6eJMV8afa8FQ7+sTeRcvzZQn91PTeFm8o+oxbpMERmwJD
5Heerwh6jV6MJ0R75mb2HsCHyk0xgNIejdHb13Q9u+oA0A+4252uS5LA39bh
+5NA/onSCHscq9YdaV2YWMeRWD7PLK+0wBzhzUidpNono7H7ZHTpCsH4Tygl
Bs0qSUb+nfnqSqGljSVTaa6MMhxIymDsGboI6j8+ykNqE1Ex/ylWpg689DpR
IKP0yDaC4z4RK8lJeADEC76ZPcZ1t+xQSXFWIY7PYLEQmNoEK1U1YNHV2tbf
xpjZ9IRPoNbY95jsp08oog+2ZnhAt7bItbF0xW4dX8PDsx8x4jnqGGYZ2nRO
xmu+QfodpyAtGwBYAmBVgzPnN3F3HsqMPmB6JirT29kYGYCTVfg4V2gHbBkr
BW1/VRShodzVrKwAl//xFvGq5B47917Dz3xOJnFsfAmHQY1Fn0bxQfE5CRce
Jt+xUHz5FyxA39P0dYZCZkUiJXSr+PELtZ2osYEx0uYNuET2fD2hKGhTegC4
cULjU7keMzz2/5oLZ6XqtfFxxobwVW2NYQjCWbuaK4/oBKLUvzZVslStHEXA
C1UNK1Ykl62NUKD2Yh4fOk3xGuzu9w9njzVPk2T85kvxLb4gkrhAh+HEgpKf
jp0j03eD+GfVKgoVQHmwAY7c4F9b68vT2Svbu0eltEqsJ2oOrs6b9NYl8uhB
1C1jV8yL8YxdhP0Pkxe0b7ROMBRfcVfL3tx/EnsFPhE2KHnqW6khkqBczasM
Hm6uVrY5LrnkKdMe7EPeHR8+T26dlN5T30e9YZLroolqI0G6ubNdSs1Tr2nm
Vdp25mWB5I+Vz2ppDRG30k5PDzj1RVEje2e0nvPfZ5593xP//0BZrN8J8pMs
S2Kmkwp7GIw4QAkvu1Hrdcdb/2u74vfEMoN5gJVi3AcA8dbjU23u06sr4EEi
LWLaBu9OVhx1gyMMXfihfZaFQebx2gnmMC8Y6+8M8X6djxFQTDpoTTjgPdbY
IL0cGhh5QqyIdK4cwei11YQLPXw6nshkd+85E54hjC1Xc/V6lGXxmcKsYXGD
CIGBrqDPenTHZVUh9ukubFJzzTx1HH9CVeUEQ4hfDkcrq3oum7g/sd2sDWCa
i5XgPx6z3ARUvuqIew3lHQkUV8kGjHXIBxqS/JP1Z2SpwELT1uTpME36YNze
85mWlrqsMCPXvMXx2cAguXTVHwi9yzlkDAwLKRQT8kwHlWR5kfwQ3QnNPJ6i
6SZkUqeG0K38PnbL15ApVysOQdjAmvTjcHu2zTwecgFhkjaCu9xPnKUfsQqe
5Ilcv5HZ43oJwUg/AvFoGwJQhQ+6Ke/a1zaS4kE4Vp0uCOUEhbcbxLAViuTu
hqRumIkEFtF2PQ8tAlytmarZCRNkIJU9xm3V1UxIUlFOqfc80b50SURbTyRP
s0l+6Mo3o/G90l9MHzrB/XOR/0vl8wzuQksh8GcAJxHziubG3CZ7jycttHgv
PFeBSW8esekMzWVgoVtpJegcfDJWPzgI5ZMYjf2rEecBSETtICYtMOY4s2Nu
UgazuDkf+wQpQpKlP0yL1VWTHLfcRLt4cTusMoBl1E5qywLTcccwfjDw8kXj
Sg+pbZlt1C6vsh3+SyOqR5VLJlvzt8GhLNZoSLM7Jv3UNKBFUBNLFuCH4iDm
sLVeOsE45i8zpK/1j2ucAGeslHmZmGwAWwQ+ZFOHQwQcqYvkk2DWBxUWbK3/
MmPWL78MDy4yJJtfywd1DY3wM7FclNvWW1Cc4af9sohsv3W3TtWrV/n9JDqS
PhCJtlmkGeuXUOD1TkOMmJfTL8AEoyFDdbVjrGaADPh64nzb1E4vO7r8JRGT
sz8ZdBF8H5zuTs4m+jcLXVl84YaK5rOXtN+Cx4NKFbcaJ8iD0nAq5uRzIk5J
Aw+JhmsKoPHuWTe442/rfrqzK70Wptzo+h13LpIrbx2EdYpX0Sj1/75gKyIn
2oCMn/L4vGhmUHlCGpUr22aO5bxkyjn5/+bfedUhLYUu1zczGMVopohPlrg9
JcKK6x695LF+18r07IkeV2Hqg2C0dghc+xVSQqvGaNsrPgCSTcRRTjFKL2mc
aFqqlSe96MpJj5UESzXcfsRWMtQdCk+g9Bz6gDn//YcMyEcKXKirn/DSx6Yw
60mlxgro+cp5eN0hgG3RGePvonhx7+Jn6bc3BfCxFj4zpaRkHMDkKlWowakV
tHQ8XwC3fz8SCcpHgdBoRiCr3sKX+Iba3XrjcBBgWIyfC/fWhfA6dXKcIjmC
dglmSRdfd15AVvnvGQauNHd4pj+vgvycPIskgKE992VnhnodoqTA+pWPNxBf
9cHCSbDFwyfelxuYU8nTXTjpyDdJMoTODoA93v1tClGtVeO1Jk4YkMjuXKXS
beEBdqF0hLBuWpnDjR3vohf/ElFpNPe8iu76rM9Z8O9g1pciGBhV8SwN32U/
gg6RpL1ZN91Gi1b9/2BXLqLBPqAsCYsuYvGqtDn5fCUppnzion+LB+u3KDHx
VoM14BFQ1W2Bx31fLLZMPt/YksaazVBmUzRp5Ju3EOEV3R3YTsH63dLsZrD3
rS09kq+Nn0rnn6DP/Xe84Gp9QezBCe1f+LeyCF2j3NgAZHRMSezWMW8lFq2x
mUIBqeDiHuYwQBPfkljhLqej0rJZqmhM4tYpNSGAdfKmjapyoT3BzQdsYQdr
2i8FC2zOJKF7G55klpBRQnyJ66/hsuTCPS/CTP8aT5dXJGAW5gg5/NxC/gh6
ayB/twKc2opcioxR/Ha/r3ER26IiZeYtrviLR9/o3o1H75bU7QztD0tA4OoQ
JaKi9yzvT5t7yD7eXA4YB5pWRkKYPumF0VVU0oIszixDwQJQRI3NfX6q4fpk
Rt7nol83SuImO6cZSX5PBO2aofi8WYYQUJBfnORbfdcd94j5fM5A+cX9bbi1
0OVDVwAkeCbBidh62yhjSlgIs6YIWEVmJR/vXkK0L4a8jzgNupkZUvNkeIdW
ccqmIzz4f6wDy89O/8Rc8AufJWYy97AykC87KlQNS+acO5klTpGDvWARJtuZ
6aM8qNVXExRQex/fWkfOKOzu8Gfwf2QGbbMMlnkQ5lWW8p5rM7aSb7WmqOfW
cd8O4Y9zV7OsJsqwgQLywVmpYJPs6qiaL81u4kZcp8Su2PBtCd5a6/hc9uRe
s+ul4/rSwMamwlJPMPV0ukeSgeZaUsEVVkzHPhQpr6IvjADjs+AtQ1WzJsqC
+nsuuSQZWMCMRHbA3ijWIZaMw1nV943wh/AbYx506orJnY3ozqbFEVdN9M9B
/JipV9/nmRnZwYmnv5yEDpRpbxCcU+Ke5mf/x2MfEb+THIbF6+l1eNzWz/9R
NCUtJWSBZWVPaVFgIpPAo8zthInoouJ6yqtdbRAUTo7b6M6bBKQRAYoS57k/
ayQ7Q0F4sXm9gvCLwQBuHIE0cwsrY4drNQ+Kqku9lvHVjUKjk3G/effQniOR
ZC9kyfGur0UyZDNxHcpzEENP2VS4aUwlBD06XgG/3iR9neNXSiVN0zp2yzQa
83uSuBpo1N5WNmsDW43CUjGM0haRackcZ1f7ojMQQYVUf3Raz/n2e+R+sB+Q
jhpf7AI0oM6BZw35aD0ObhwCdMi7i4cbJYW5cVWs1bOl7ibs4TK8sFbb+pdq
iw+8GXiiuqxW5a431S96hhG91uFwellDScZgzWk16vyxBZ+adapd5N7hJ/oT
IHoHcdo9D+kGToGI4vlJ2GxSefnseqWvowj0ivNvP6rS5o1E4W8Y9N1xp3da
idbY88gHfb5Tef3AKNSg+XEqDE4caYnBvlHJUZH44zZ+8lD+lssDZWDMrbo7
l2R6ckSJj/3vctVr+0I+uVgdWOEmqXIK0GdUxC3yBvI/VwxGPPRfT/OIFZbR
09rFgps0nDJnHop/y7eDadz+0cjfN2DZHv47HOTN2L4fQ+gebFQuUiiC9NOI
QWwy20+daz50a78yvtGwt+HLTbjEyr9cyydUSaOPXUvR8kGnsuvMpirDcoh6
aFNVMunkaAh4vLOAYYpLIoJjjK9xKU1Ked2Y1y+gYYGZNcvUcgfPK6t4p4SH
vr4s4CtcOfhWvLRqMXwy8BCmBy0EW7G7gywscE+m2CkgpVNP5XtJosBqgXtg
ydjvgoUca9p0Mg3Vd7su8Pkzv1wB9FEqlX7JH6VW+0xR+XBPmHforUdXP3Zn
SPaDlBXkiDgX5PgdUQwUMK/r8NZA1sYftIEpPzWpMXfsLCaRbWR1RUHrIJkG
hBc4HkSr+wwnLa5aKF3iNXMGPhethpnS3bdAmEBPg9o75bD++CpzIJSGriwI
+i8DWvgOoUn1DxfnXXyceFtMArI7cro/f9pYAUrBrbkPsOHnsUtJJDH8bG3T
JwdRq1j9e7uo3M5Ky2HiMiv4ao8wE+LbSBu7B53L1ehWcG5iCmJghNymCQNv
Ic1ANXi6xvPMzmmulxDQ7up6ZjhJQMwawmJvfA3oJCJXjD78o3VsJDXCCDbK
qI5/+k3pIm7aCdU6K5X0+KC44Uxu36RkmvMKc8WA/qEEYOYsuY3ChxMkdmKu
8hHkYq3p3/pwFIoe4r+w8sm7MMtoex9Kcgge4/ITmNPPAWI0UBdpkNSbmslb
mNGIFKlza/gdGXYY1BJwSUZ6PsCnmPft6QotYiAqyLTi0bAQWvl7Mw4isRuu
xfg1LSa7lxx8Jf5aZpeHYFfkdZcVjJfjSN6iH4s/bHy8feHea/6lcUih6P9w
pewxcitX20cbK7QHFW62mq+bW2hQuKHd8vRfq/FGpoATJSrdTEicxgwHjeD/
LHYLjU/KKeHNkp3Dk485A6uSBv/m/eA76AoBRM2qehHUVmIhC7SBvVCSTwGD
zJ0NJhj+AmA6tSLAyr/21kVOTvucGBhnt0790aiptxwXn81/c6CUFj6IbOUz
DBbEoSczFQ2qbXhwefUoyVS6sl6T0lPDNeFkm8bpwAOmpGs7NjWG9PBDGLCW
fIFu6lSt3GsoVYKwNQy3YR79gdwYJOwMmhDp2iKYKgbupoNXV6lJf8HYtSbh
SxreUpGQ3vl28XReBXQoCoXKrTl2Rvy1byjO0SQkhKp4NN+nrErPi2ePNRIW
3CNPBkCeXnfzuxhtwf3dVF0Ad9v8x05JDZ4XOoDF2xehJtZrb/rJzpepp5yT
JDzqK/WTR82aIs8GjSCOVz0JI1BomLMeWmD/rv4FcXUFk8SK61zvHSIviTgj
25941j4hJVOZf8AuFU2EYNxuA/W+k/DN8HA43a0HLvtjHG+iz+Lx2fxlGKWq
qbBVbK4EQQVVIMCjzt5bBhQpvQxwf99vNYgLMVtKY1iimZCSmmFfgeBBCfdG
VTeLG7WzNgOL/RLQYr/Onq5bAiW82Db8+NJWExKHPJ9RawVVeBzTG+YVBGUU
Z6XAkoIxJfFyTDjamCgaArQgxsSxPJ+3K8XC3XTEH4c3EapSpzpbcfvFVNOB
Ap0MDJmGwwHDO2zonDNScjmbPKTIgDTjROMoRdMrl4B5lAdBJyWcQRfgawDE
GONrSr7oAMycKWPt2L7j+5dZQ3njq9/cSvyXNbrsNtrpkIVVu6iLtiyCKDX2
yNAbI8epphpdWUwu/QeR8KJX7YfbJPfew+/rfQoH/Mt7yCSBc5tloVaCmSAz
pCH4DXzCF6lyzQUm3RCX2P3S2eBmvRkyANXMP1uYuk8Ns5hfr/yNi/IWHTFj
X0n55q2qjVGrr08BA554NSEMJbTb3aEkWISmO+Fn78bmmmsQTIeEHDp2f5wK
jGws5+7foUjJMVgN9tlfMvdTckym3AviOZ2Xaxsd2o3XEoRIkwJwVSuTLcpj
F888CCkhlbJuBuvKrQ2bLOiQitlVeFFm6zKFnN66V+ZFE/NwOqFA7MIHVkNd
IlEgU1M4TnSBPzvJsso8/Cs3e4uR2wWyyyJCe+YCIMcrzktSWoZU5o9QXF75
9BgJ7iGkhVS71YyD9KF88I+AoJ6JJe4J0F+4BI7CQ81pB48UjkoMh8kGnRC/
eG+ka14TpzIO3TyA+3dTBpMvImlxHBfnp24VyqBxipvBqWkHRQ9j+3MI6Kv9
yUsKSlrhHzRyo26Nm+EaKPx6anGcBucIMdsrFHaI6ZutYsCN4cNqzcj2uRTH
obg9XkX0+GA8Xcpoz5VRY/lKvCqRf45fLKJurNkCy2Cac96TV69ObCR7CVN5
bMXw+J4icmGQCKxAsPaW2mWmUBOOV/6k3UKRqK9dZBRAwM9jyUNa4XD97I8I
fgLhXpAlKHFXoFvLIvHLINnJS4Sb/wpcrId8KQ31Xwd46H0KXC0vfb9H/COQ
IMYdHYrv2nb5Q+2MK2JMSPIyuMRNWju2smepO+s17X9224siSrakDG8xBZzJ
zMb0VHffjsqV30eBRLUP8HVfvOxd2QuLWDA6ZY0ibwJJh9c7R+d7EgpSTbHo
LfRUyPjrlonE0ZI7ahXzIEok2199a4wIDhScQvpvesZ+Ufn8t9uo5OXtO5Tu
I4PFY81wFfBNu4HbkD+1ptbcBP4NpZJRCuxl3Lh96MtSMVeg4GPzhCvITRLs
IDwpaVGuRI5Br3E5PMIAkEtqY5BIjbi6EVC64pF7e5NgvGRkq4CnSiQHL7b1
FKxBD8DTXT9sT6w7ury84mKx4ZS76sbF8+eF6g8gL9WJOmhEyuPisKrmT0qZ
h6GwYB53KI03r7cQnHS7GPE1A+a5rTlWwJjAAydGN5CgKJbgxBGEryPeWl9d
gXDYlWCDSA+ar8f20XXkSa9MJWEjz8ITM5RHe6WZ4UMBzzMa234tM8BgRPxn
HJejjdOtN/3tK1Mm8jo3z/uovZaXEfCrNq1YypTWZxAN6MlbRB/NLDU5SiCy
nIY+2Qdq4Rpl2gSyjiU/6+l/BRBvqrJ6KzqzuHBL/BvQg8yVNuwMUNJsBwFw
Jl8VL7rwSZfcibPHcrwrUgIIX71N7zY09sMn9BOERm+5hFqqFDNeXnldlfim
tZQHTPhzuNvbbfpEV+doyOKvjYAGtANEK1upmXx5IxhaFIr3JI4hv20K6FWq
pFJi0ep8N1dRAYwzZgBn01t0K5tKntDYf2T8B5OmkJJCyTJp58vKikHg22W2
YNrVtdFZKNp5/YtT0Tw1p7tuFUHqXs2fVi14sb5YmccmmdaU+jfbbcQEaNTP
spASsQyGdZi/2VOeRD0cJ8VslRJtGS/B5JdUq7AfY7tdjapsu1o53s/o+LBp
OZq0UxDUg4bp2xzGrnismmjdEvwc3wju7ZJTKY0g/doSVhUKdfSOlDHaAB6F
PuQc0AlHaD0pfB6CCGvULajPkGLyUEsCnuhVI0/FoPPsY2NLMcSvRm9RS35J
//LuihhaaxfDOaHZxxN+FTXu6tMIcp7AsufJwqTlJEk6Qdspiy+lF/56PYtK
iWLF1kn/EEeKQLD3+dxW6C2Xj43ZfATlqC3jQH2esZznR08Rbbqbh4/Z1jRI
7hpTEm/5AUm23oUmoLIUtaFZvWV2IBWBmXOamNOKnz+zBUvILcPLZ9fG9wde
jmWJobvcH9wU88lV3e3hWz4zaVCN6TW00UzuNoyFFdEKXRFw0owq9Jm0dvmM
LaDS3Rq6JvPlFXFnMcNM1gGEGg9n5q5iWajpJz9BA72TMTkI4ZMIXB36Obil
jIb4fzA2XAIhaXp9PtwWpBJMIoccP142/HSIhq2yOTb4aHMVXcmHCcJX0nOy
hqw+VMiwWwl6fBymTutnrZT4a21NX91hP2z8YNd5MnF2zTdHOUrsdj7ju6Pd
RhKwCz6b9lDK5J37zbs+X2+F9W60qi/KeyBbajUdtmVzz62w8Ybc8YP0F7k0
6hrd/tHemrgJce3+XXcAdvd3n/TD4CEymwJDKrDZ9pDMQ4H9nA1rgUs73phA
pAqoKygKuKYBvUoVfMl4dsP6kZjMtwZew+5AnQcpYEzO/R1EDLCJ9zHAdmUl
G8BBR4xEI8YBxqv8uiiUUprw8XjisEo8b5Yk8+mEmpeSOHP2tXgwzKUlGwTp
pVZk8H8vEaUArKWsxZytbdNCGUy31jc+/qmP+z+MTubU6eF1Bq9g+YH1n/xJ
poZDgfH8SO9wrhPRHOu4gK8ORN1vkZO2EW5PRTvkhZqJ8FmUVMo8Tp54wuyV
qAU35dDbgOfhhnY9Oo+AbYGHLPiMijaJzQh+m8Ll4y8ldIl0ZxYH4HuVsyWr
LYOT2lMmhS5sG5gRnDDKJlYajkncw56aTsxL78tNis5+7xXD+hoq+uwunYp0
wkFui3Vlo/J85Xtj4OTHS1cX7PN0enhRG7/G4VQu4al+CZfz4tiMkLF4qxT9
nEvsvjiONeYY0RLsFbMm4nybIO0XKD/2BX/PAhGCr7x8NY7ybfodv4WEaSij
ndqrTwlfLNUGBfJ0pLLXh/lRONprbK2n6nNBKbEEnFiFidS5LOiRW7HP6roI
7iCt7m3auu5RdjvhxuHP1cI/HQ6zGIXWb3jxUktJVaq/PppF9DA3oEsYPU+X
EBAvsNk96lHNVG5C/gnFHLG1HfQl72CHHyzZchi4xqtB0mSapfaO826+vd0a
COQ92i3PwfSXUWnDUa/B39G6OOVbCThDcNL+1JMf37Z8cJLw60u9BikCfh05
8Io2fQRBqsQmv1i+dB9JKQLzO2+csbNe6GagQgUNTHrr72W3leKwr2ztn5nq
8+g3tAT/7Ixv98r92UL+owjSRlXScrZvCVtS0mM5apSmVfDmovIheKoyhsct
cDv/Nnn3whQOLyVf4MOETR/tP6jksa6aP5nzjsXy1Zfbl3vdElOnRYguMEOr
wIu0QFB+M1g4y9mb2ekf01zrRVdjs6wiA1ChWNW0xwMEE9FBQW3UMhI7V5dK
aE03Sm8eePBfXt1vPQbfzZUUlq3Yn0laPiL2M7QJrrDT/JOlF/cQsn8g6xCN
wVZzbAPpb24MiWxWwd068v5NflzddageTuA8IC17gzEYxRnWaEW7Z2BjIK9H
j5oPiEiQ9cEOext6UF/gMKwvX7voktaak1QMPDiLNLZIkf/A9nqGU5PX/Hmc
Brhy04nfSrLyJWMpLzNIVfmlybYepJlF2pM6SpNToynYAEgB1PQWwzt0WifG
AjE2knKQprDFk5wnzzerjinH8ktqG9mbsu1hpFmiYbcJQeBEBx8ir1AApCAe
3COkW3o5GRCratxa24gW7NdceYwFJBDBStUYCjibZYbD5afrCT7BeIVLkhPx
MWgB4ABD2icEbTk1WL1f4TUZe9gL5e27WdaTJDb58xxREeSKhGvDVTjBpEde
v4tio1vR+9Fa0lK8+MF4gIs5SQl8bTQawOnC0xBfINgu5/PvxrMXlj4txAU5
Dxcaxb3eRrOWHuWcNihpHiBVbwKQQHYScbFeyXvsJNSM3xqjLVc7QlyoMERz
6fsFK3WKfyN7/mYe9sKjvFo/491GG3zjzXAJkdMupOk/GXwETDYWIuFme5iO
nT3SXRG/QpX+rj7mQGSJFKAts4e/lDL2OJcozlikIsLqFt2l0hUNSevAUCcf
Mpq2jiKlY2i9qOUTMKwAr7zM1T6HNDk9VCkC7BFLAU/tHLpi3j2qXvtoZIEj
sPdqRThvb9vJxj2xc2AR4dBeldYJO6Fv/99Zymr1XDDGUCcsXEP48K8hxT/h
AFdRy+iNeH21+lKFzABf8jY5fdb8iL+OgYNTNSBesZrhbPQffKLCfcLYLBK7
xowB5bCnqmcdIvyi95+BkHmGzPM4lWE82zgqgDdRs7MALB+ek6RYSYApZjiP
zN0u7dGlgGEirLjg2bU95x4f1O9/YeSoWs4PlIAObYsOxdp1Ym1b7qCmPQ9Y
UohFA16Nu4Ljyq7me/zcQtDHATBBa7W1pOXAJQuQ+9SFUJwZmhSWJVcKiiVH
tLNBdk2WsazehZpUc/MaaPcRrSLvoLXxeWshvksVOwepH/RwdrPdi5n5fMnw
lR9do3YtfWLwJS9i43GptcHTLSUlGhTtoAspCSceHROEUGNbCBuU5Ij4uD5i
dj0e+bm07Gr6deKDe4bRTdoDcfIiemPHXhHqrNJTR2Jg606/QsB+cA1mXgk2
kkr6p7QCDJPdPMAyEwjS3EhkrPIw+P8e45Jf+dIW1VL6MRDm3lC3AuuTKiUf
ek60+wg5GhqbfpcxrGZ5zAgFDV+MW/Jw+pEgUel5DYbI0UUg0guIzeWfdm69
RtDhIhW4AEKs1klCqfAOaZDaL7C39N7yzPf05pMZlS3EcuvLTH8VpI5tXVDI
vXwtKUXE8DdvLcsv/Jc2jrInP38Vo0Cflj+IXuyCtk6CR2dk2vywo1haD56i
b/L4g1uQc11S02reOeIjvWtvJsJghpEutxhQ05E9fxTJbef7n5WwhFaXlk5G
KMAuQ8rDF8W9PViEEjMXw7KyvMASQH+ZrECdSInpAZMHPh/5E+9mm3ZDRw5W
uZLmEKzjSUJ2F+6zKjySKCWxDBwpDoxKTD2KFRqk07BofCfQ3ijEI0/Ek37B
1XB7me/2pV9Y1BEBmZnGYT0gHkEXuVYECXRatnwRQCj7sWyBjY2IA681UJBN
W29I5hptUEVxiGgXBpku2WGEAaR1kk/X0d5iQLmU3yBDE1DzTiq1syWLwHun
GI/FOjq/4pR5Zc8ai+HE8dzjScIIw2ohddZwOX6BVxm5dJUuDHvtiDiIaOr8
qsIc/kQmGKkcQ86IoP8IcNlZAZ5t1i+Sz5INlGtrl76sBC416ic4U4vQRWP9
tfE11I7aW9rizrUVQ37BuoKATeFIqRpFHX1SOhd14p5yV1O/BA+roqjJ4hlT
FxW/MKaeD+LMhUSUJb+/+9I/DJSgtFiJ//vc6DB+9o5LWhBrCAZB9H/QvLlh
0KvNDGOeTzXFMenRyNqEsxdTb5pT7It2u5IuMXysIYw8xqNuGmT+DYmIQ8r9
PWo68AUqxHgl6ztPDMoAcFxiffjq/uTpq3bJ9PuDCLsvkTIsB/yZHtsG9qFs
Pk4THlWG+E+3OQzToSir+/8WFSxaSUxYg5L3hVhWCCzeXVIx8Fgkh9FA+/lK
JvB5Dqdy448Eq1zkxlShKpvfSJy2n1039xsXU7vHVo2gWqTAHNZAvPp6w87Y
dj7FzS/lm5K5V0QUa+kjcvaroTTUBeJGRLEgxUXODV/4Q65VwhRj14jkEULZ
LOL6roMhqR12NcU+mas4sMbmPH54rFZ2EMyGzRDjlMSXe4WP0DSPISen1Im/
yB3ofVElRzumnKp0apYgNXjL0s4f5cg1B5RIGOLFp1zqw4bZw0mccd0Tgc6p
ZZIPDEOx5ZOgJX7ebX0uFSUjcMartc6SPr0PviIg5ayddvaDsxRJMI4J54nx
PaSss3VI1QPT5ktjnpC5wIFbzeLtJNDJg9fSxBQCF6MDbx67wHgyZR5fx2Gc
ENxjD9hls1wWjfpyV2mKkV/NVO7g9Zz2dgI+pKNPFydEbknrcVDTqvxfNdGM
WyiQfhyRu8jmnbZcJkZ3Tv0sJBJ590r1hZw0njUtnbK7FZ7RwvFaU5OnujP3
0dN0kCYITRcN8oWrJ0qeFhE3j9dJTgggzfWYOE1BsgB1A9y0Qs89jPXw5W4G
LhqBjRxCWqztvmXyxAhO7pNo9wDgA/8paj8vzu9A2jJG40m9BU8Dow/N6Dck
9nh9Pm0L1TCHK1sLHcrSsBEnLmYf0aTzc4MilWyvIcfPaCN12/YzpWvm3+Yl
WdUQsvaALBqc5L0YNqjDpAoNDtf24hsVwryGyw7I1ZrOSZL6iUG6M5TNKuji
LBWCXO2uqx5PRQtOZ7JcPU+j3lHMXhT2b2612SGkkW2oHTv4AFmFLFnf1Qfi
+fp0AX+HoNTdGC8xdk3xc5NzpU5NYqgwmohNrxV/1PNb57jh63gEPqMLisUB
yDCipmyyZHaYs2aWx/aV1JRbnC+6/kStNMpzfNC56a2dJgzZbjzt21UQB3M2
zaAl16Qmue6Afh+XLWvDsD36Cpjenql8vdtbN6UJ5Nvo7gjjh1583eqCUa9x
AAmMxffUogFfBomauup187CkH1OCby5tXXWiw1uMEYmDERQFLRBe8zNFbDio
r5wYshKIOJkarAOBgcO8/ijDvZAxIKceWrIUOs1I4T90I6q9FQ2MMBzveL9Z
dVnvj0K4OADDDagaiMqvGWjrVeOyL+QLcaLQIh29BSCTREP24x42Zmf/5ztI
0n1VO9g8vqdyh4M4yKZ13UfgBwAxkdmhqhqQMGRm/zQld+Cqny50ASrR5/Mq
N/PAAuxaKAh3Ozrjtyr1uaYfEiWgyg19CRFy11Qk2saNTT9G17grnzAqMlJQ
JWtb5Aj9b6v4qdAh/NTxrYdmLSnjP/jX6TsJs8dmg5Nk4gzrS6sHySxRPQG8
p1Y/pddhHlQ642uDXkGLzTyqVbAwEab6iXe9q+OrS+5bh5lU9rbeLKQ4hIoX
YKIHOpRRMyEujyasOVYgy+0sZRmCdPTptwMmVnjnHnIGfr8OQfPgt0+ZO5PH
N0oZQTnzx+I7RRqg2f58AUVfvpQGLbK/I6F32YrMC1PaRLwy1n4GvR6XwCbH
8cifemvvSOMPCX3rMrwXWwnbbDkfVXNxK+WmZBzquBCYWuG3rg8y8hAIcxBy
w4GDOVzALkq/b6Fwb79f03IW8lSLX6CI2RMl3gH+dx76eBzHFcfy/2x9WVsP
GxK0JOitYplUxIC0YbpIYNFyHikYQjjfrFdPDCl+tRgkHaQSP4LNzUkQgn2j
/DTGIvn197cT3hpNALkeeCk5DBe65rM2OlyJQMvu92CsV0/NQdlQ7F6yjJKN
Lp0/ISe2l3D0EWhEsavyfcFxm9mVdusl84b2QxuI0ksTEvCW84kdIzwUWksO
IzZzNZW+AjuQTDaKcl0whIvHo9Tepdznmu2iIRTtZTw1/EHGy3G7LVfyXG2u
Pcrrs7ICVbahmCY+KSdqKxBiortpaczDpkjSHyQxESBLaWho2BNSnAFlyZEz
VPBZmmNYw6SQ901ml9Papt/7EWCOpKhmVmRUEQghXwv58tZMsz/nl0RVz129
1s2pD4bdc1N91MlYjmg/owF/O6DzB0x5JxvDmRG5Go8PW7r6glaIqS76t+3O
8KJVvz+FPs77I6xyEbLwGrdyOB+Jgh4zxPXZatRjW+9FQkce9b46mjKqLCyv
sp/i7GTACM6cX5ShllXcRuW+Bk6STEJvAXsbf5rqRCJCzK1isA1lkBntcmtx
v1XHhqQtCedrCUcDWXuqiv2eZIAlTbNx+J9Psa66L2gLHMPAwH6BWZhKPNbm
gE0zEgw6+fEzve+hbBv/ERurFvD5GdF4kvbtU79blIZS4FKRmqXHhuz849V4
kio0wvWv14VX0kr3/py76DmmqjV68T/1cZespeudaUi3d7FNGRws8E+mBGju
BUkiuwtli5uqYoE6/k8I374eQC17pwwHNFYeIUGqX+e5gRJBzRlvF/zwDJBT
1OoaqzeJVzULU42/ODDm4iE48V43yKZXM707c8n5X2r1LiIkhNLP0AWEuByj
wusXQdtP1Ukp9NO0A8xcO1UeReSFnIWBzQ2bg1rK+Fz/kxLEAGk0qfNdr5Tz
h/s8cO01JayazxBIVFNh3tNUm0xXRYWlwS/e4naKYgoJc8Icx6mRyk5PjaSu
jrUvXhH/pZ/Efr7FdqVg+ZBQ8alz30Ed96xyjwV+lU8+ViMEoyYA1rOCfvS6
V3k9QEdJ+YDFQe9snsFE9HcMipv17lecsNRy2WzdyjFSyWD8LhON+c2VkeaB
N4yBzBY+C1pLZ7k2OP3U9uLi5YT/VMGzzjfWrhV3Q9jUK1oFm4aT5bMzmnWi
fejP89DUV+70jET0CS8AVGk+SHogQvAAPgURTAfxVSfciWl8rHME8jVUfQyV
HLbua9eRsG+R9tUjt6108zk2Cp5xUohfs8oaW/uLgMTHaSRSaWCeJ0KTqjeH
8a1p8XuGNAAYGnNgNcNbJ8Kc90szktQrr/LvfDbbU6Eq6QZYrZPlAdMMRnAb
qvcoXnWENFbOUb3QEcdibGFRxvnvQRCIR59+NRM3ay+aqfFQOunh621WnB/U
zEksKdS3GdtSCinkyyRUVtdlHS3gtVnMTkTW/hL0uB1dtTUHUSkErCPYhP3g
XBG1dXs8IbTTR5o3Kj7n7DQqvvaj+42Ys2lOsLw02bReVEn51pAcgATj9w6U
poSJ+9nBAsZAhetJ4zChSZD5IgqgL5YiOA8buB8vRq0jC4pyGxgboPZLNEan
SlxF85Wk8Z364/RqHwGvagoTEZhDqkkUX4Yze4JJs/bEyk9Aet07c3dcgq33
PZTt5Bu3bmZi9wxiDtqaVWR/JVZREm2gzm7uaZO4hCmzhmkuWjFQw2l1Z6nR
rRGLyitbQdzEABG/b46aQm59HyL7SYDHYTSDa2GYTjQR6ccOHH/RhKFOlmy9
QCacwB9dduNmdaDXfrAZqewxTyr79M0bKt+J5XYmX8i+fvF9+STwM5HJ3orK
JfWyp/tIGBmp+Tlar7pt3Dtnga9AB0L1rbeIxn3EGYsgZMuKxDSPQRdRntjx
txnr/BFv+vQyZmiOXTRcI48AQGjYjiaXgUcuA8tPqTpYnCAQxTUcvGbDbCDI
mqmYtaE2YSRF5gcp0bTnXiGdiiI8qgscuK5EIpc3rOlST45QJ5cxDMwW/eGt
37QONM2BSAV28qjyVj93ht7m6edai4d9B52LSIAqwst+bvXnlaw38hH8Lu+Q
W6A5i8F5jIIHqeSV082ervXjHkfLQD54Ek2XvlEl4Cl3rB2v/WcKkUaf8eZN
K+EjGsDvoZ5bMSsFjy6/pwoT6ic36s6UKnvJNBp7zk67ZB8tF6SN7VJmqmqq
TmoWmSdpkg7Y+phXYuEM+iJfy20QVViUEQZ12VyhiZ5ukrqZ2kYo/Vz0o/Mr
74gFpR6vf8LzmOkA/rTIejDqdg+MqJQyoHTNO+Hm4kXWYR41NFltSAJEBfQj
nqTtBHf2UO8Z2e+zo0gCvljQ3JqsaodU1xnMYSVetDaXka4QsRdBTkW0AysD
04mp1SMi5bmrjr495fJJUJL+6AVSbgLu+AqcPNB6f7OvJ95NeqLC2EGyD+S3
YHoKSq0eE4zSyM3QPro8ayaypAnDqT3JzMxRoJaxgfb62WdVk0sjCSIF+cvE
OB2fmD0SDTEEgLYsIcLSGMizOrvRWaBGlWMT2TTq1xY++XrBdLFzNuxo5c66
Za5XbcXl1A6Cx54IJE4fYh0jdkPJbtcYqwrgidXgvdQY42kkafTtQVGgXLcC
2ARU7xyGC1T+qjncdK/T6bSg+XS1Yyb+y2hiWzxwrwSUWYPzRnBWtx6lnm+m
dUhRdiK8qwRPLFYoNJbLe3JG9Af+gYzEd74Ran62m0hSzAELACu9eJNKlYgL
+YL9G6UKXsme/2XtCYDCkFiVvyx0YKqoid8n8MuETRY98foxU4zT0C2lMtty
m8kNgAnizClVC1rr/SUT5to82wbJb+nN6v0HoN9zRq43ChxthKUC7fcLJcwv
0ItXTMib+ZNDpg9sJLTV+hUL+Y73GKvWkusHxa0qONngeaExZi4doPrRNDNb
jdDc4kVfs6FHYQ/GgDYWF4nFKSrNRWHSW1jCHPAMpA+xDDUTZelEWFIYdrZU
F8b/yPx35TRUOlfV9hDElQz52JNJDV+ukJdqsIvS9nmCK2RLW/2pLda2EgN5
yo2KHVKu/hLT5vafmJKMgKXHOlX/cgqxrAm7oPEdJ5hg3BVTdmrMCR0ioK24
A5wMJW3xEyLdtZEUxVraK9pX4RQJBZoEztwf4S0o1zQvNFwpD1nKr6y0u9YQ
xyoUaxMr3xacJGfXma++bICtBnUcSDFCrESgLBkzj4QJR1GQpMJtgzLXC7Ui
5XEmhyue8y3n2DY4dSSkOSszv7YcGduF0TL9F5cqEWMMHsCuL4uJp5dSH9Q3
K9iw2Yqxvjil5sSshYFQ80NLt90HI/FJdr9K1LFvzS288r93McoEOWnykz9P
Y6qAtt5dXQbwCPKt54dAjH2kMoGLVe7dGejQPJDknZcOAOIavjatV6MxrgZz
OJB2LOBjE6LJtV5zhvqzEZ/19DNbbWr8lhCYLVnu2Syw5HcSFFRHGXuJSawa
QMyFuR0eRXshfsaPngYrsXABiWPdVV4OEP50B6rELIOBr1DYlbNwV0HgjlUB
kfGqGBY1s3Bwfe73giDOYsl5eIrJqWnLHRk/9EYINhNjEvHWT+QKqnS8pa7x
GLWurBc9x5H1a1dPTh+DNmjp8r5PxJkOj8jkA/meuHOTJHxdXnSNRT6+hMRy
CAN689AhnxOh3fQlx2S25dOZEBHIyjZFk0rRWufkT/zhFC6gYsGruag2aXxe
4D5ASvPgL4XwgCfZADck2+oc1G4DvJr691YEX6tjFSGI90Ym0nRLp2cRrQB/
fMd4VlXOa7cqeEXVyNhYty55FshsrX/vWuNHyaeIaRwIhMPF18ZT+tyj+R5K
DEpAJKG4ZtK64UjFoLVdZi3L3oGjWVI/qnHHIJ3LVtc9oZGyCqDhQPh6gUAf
vVTGLJTG9v13XLNxF+dSPV/e13r1x00YdPOAQ1G9st+yYsTIed3t6HQBYigZ
auY5zftmHrCoZSkZg7BOflea2aNW7ZCgrGCwpJczekFlcMu4ccHRY2VATfJ4
lv6X7oyTE6B7LVZzNcqifNpuR8aLCx47rN0aXRy6gaZ+uyycwxOYrvzmaibt
NX3M7WKchKR6zsOy+G2zpAy6+jZgaabynmrfJh8DS3yjP/jze8QFDsBmtjT7
AtRLHLswCk0vfn2QsKbpurOvN0DQ97kkkZ1G2glfEiYK+8BEDIJy30uSVszf
Z0MbDHS0KkkFSABHCmKhFYPljAEyREQbdjWGuH5oe7cgVhkuR3oEfQMgdteY
wzReKrlZwF/iWWaGk7vV3hN6hdhWwziYaQOUP76CsFVW8RoZPgpguDwl16AL
ICatji+Nrd2HALT2S+xufVP9YG2uNu74UOhaTDDtfMQGm4MxiEixqYOFTW7y
wD3qiF8Yt0N+d5CDruouCF5ZW6KJ3N/em+7n8zmrc+sMNgI67ksKQdlnahAO
4CCm2NeClldQePQh9ruGgfaYSNrMpcz/UgPpS2LaE8JoXaJP1RxlYe8hkvTC
VRYzmNmLPun6pTGtlATWCkDYbPYYtLSQpfrUybQ6I3aWTSWTXoMjaGR5zGlo
D4HIGBAy7wiGyUbgx744uPsgxvy6TSzIFX+siHsQGVX39JUhrYtDWTeXS8Qm
lQQvTFT6JVK3z86uVuIq7eCRCwWjiP05xRkytDvIdDJFZ/LzR0Xwq8Oc7wHG
qb9knYx6JD8qqqUe148E/Vcw2ZMPnD0nEXfzCQrjdrOoYbnsPC1yElgHrwR7
oFNKZdWyySwnbSKauuS5+jP+6578BpeZ4RO4p2RsaefgZ1bmcI49xlM4r5YE
nFppJQaof1v/O6gxT2/kAIet1VEhqjsprOLdyOOd7Ws8vcBSvjN4L3+ypouK
RCyeZP4+XhTHGlnIBu6+Q7+2kUlYFHb1Ts9r2IxImP67F8xql+o1iDbv/FfD
QN8EfjwtHVEEwy3miSozjg2xEW4MgyQuE+O1Ag6Ff/qMKPVvdwLXN+qATgwD
zcIRDNGANfWdBd3V/p6G0j9XPRflEbIPp/+eB+hTpekDomNpa82IPazPQJEt
43jNTEFYyJh9UwzHptcARFXcmVXTLGsyipgMs3Xyb5jbhChqvS9X0dbm1Jyw
P/Wsw+gLeaE3w4tCLq+PQ3tvBjUOH57le+ach+ami+N/NYnEgljpskVveUo5
+jqQs5nzn3vvTgCLbch6rjwAzbVik80vVgXuTU4Wymx80NC+c1P0m3HWxbTu
AopIN8QQb4M711y04nyoSS1WRSiu2XSoj69O8v8H+OuN60EJqhjfBnSwAZq1
WwCZeq6b6xLZF2ci07Fk8JkXMdmCao6JFbKWCbCaVjdjG0JJhT834YAEItpf
1eRko4II9vNcvjvfhtuAKUPYoGLkPOmqGa757TNzEU/jPd3XBiI96EXbPv0S
tsv3UdlfTTgL5+/gmKEd+I7cBNnaGRAqpbZrI0fiRO2zMIO8bPw5dczzUzpb
nZ9mCaf79FuUI7pN/WuBaplx5jtdte3n/riCMJdJB0FOFAzxADQ5Dw/+d8Rl
y1OPiUCfSLTBhwhGtxlUeJegwxRQc/o29Af02yTmUTFX8pvJRcJCFTtKgF4N
HZK2L+hA6F01cT58sPJEVzdHKh39+mjk2S7fLzZbfqeAhl9ZO6jH6uVtJoTj
Km92OcvXo4oY9Z9TdkN9pW0Y/iNajdba9UK644GuyZJJzchy6uS/HujCXku0
pxGNCDOgV+sB6qYhszWB3cfq7Azfg9Mk3WIzt+ALoSNbgjGCuAd3pXFEHayH
TVy2ZN7406K5y/Jn+zb94HkMS46LXhjVJjIneY58frTujwJMtIfrzW13AmlR
iszv2Vl04f6CZPuAOusS9p8ZoUjVjhKUwYHiaFHWOIWS/qfMetl40j44hGmG
qMAzE6IaT6bijWqheV5XAKWBnra6LvrB9/RqNbW2DKmrqm3GMa2KuZj4MTPU
iZaqTgoRIAzVKSWDzwCTjy9ie4YI1K0wRA9j43tNEINdqYD2OT4DplN4mTX4
Rcv6hm3SJ8koiw84argikUIdOozqDlqxBCTlHT0zIhw5IWpDtEjADv1d1ka1
Oc7+ZPxfi/G0OtNBTY0W47+n5/Tvrv7y5ea94qxrB+v9O7lrK6V4OHYeoSlI
W9gWITLUYzyf77QH99wwqkJ0htcikV54/iw0TuAf9tPxebYdoGfKRYeBW7kY
g7+XKqCbkyLWtKv3rT7pFUJJ8HxGjKEwN2P0Yx3zsxVbNaaqX5kKP7CAjTwB
VPllPbGk3RIZ/lhk33P5y6Q6osSMx8yPdmq+RZySQCyEDhTmmn7h5ALkMPXB
VMXfjVo0DMuplgyiXKRva/D0qSIs3dSJyVFhXp1S3OxJNAoQJnAjuISPl5Sl
d1vQX7T99q1PiDXnIPmy2/tsCwRAUs694rQ5y81XwZKBBv+z3hxH6BxBWefB
vwx/toAdq0m9jNf8w10x22ApqMWSLmwKjCuknpwkv1/0IQVDVba2t5GGxX8S
3kxuiEXiCZzyy4e8GqWBasPNMTLc+qW+aP7fPC1ujD5DiRRsboNiZ2LYTgry
pziBplp6WaEkD1vOScyD6B1qFJVM/HRnO3+ytA+cggP6tZSSIT11dUNNJ4KQ
5Yg+1cdAb9YU7XxXvw7jV5gDrr1pbX8ljJUkKb8VJTmMyiVFJ6mgJXKrs/YO
OAngWtRIM4P2ZLMTjsu1FqQufmEmjFsyUoWwVEJJsBsCSyMUSl2+z8Z5c97m
5gXSGLvmiQwkRHXSgSbn/TCImsfEef1s8xVkeTEyUbS0L4bv9k+nIHeXW4Ph
LQ1WwBLCipd61ETq5XEKu2NNwWAUgznPuxA2/7QQU5Km2rk/5lsud1B5+1Ae
9yYrHzTKgm4jZgY2c6hmccvjKTN0iYJCHx/I6O11XmQvhRa59G/cuxLlbJys
/tumCMhgjsx6lg6QdXVppRF5o0/fp9j03mCRGs7juJJ5/GR7PEhuIZ+ho+cP
AcyJPt8GwLsggT0ldxm4JmpWtp1REVvGshPsVq8eks9/3mbfeo6v0t+sRt4K
+WDD6uON01PEbiGT7a8bUX+xwwo5aC6Zf/95KtYz4EMxksxITfKdHtyg9TWl
SFQhlyrTC/Y0De7EDQVxRfvG9KiUptPXmE15bWAZw9dx77yX84pjQLIFqmAk
f0oiZbOnJJx52TaaHBDyIhftFikUTgTjuy5hlm/OYmjExRdp5qhJxbXYO+3V
GRSe+WaHPOoTYn5s1y4d8Oc4njOtrrTUmcN7mDMcN8Aj1Pa5zWBfwiDRvRf0
a0NDGqNsHWVzX4TLQd6M8dOg7LELAeF+mE9RHqaT1YGZpslRJpetcjrHFL6h
AERFLzN6PAZKWSuKuq/ozzrh9q2DR0791gusgkkub65lS7AT+5fWyZ3tu6xj
s87qPy421Lvy1b4NKmP/zJ5N+EB5p2Yf0ib6riyFK6Z0343G8mlTSVi+/Fz8
8aZG0ZfujL3Ucgu/pnRVtZA4DXUT5acYptb/WVnoazAuDzX/gT5dcW+AJJMe
20ZgnDP16SRcllrrhuTOrwH52oTBBvuVUUAvdJtL0yRECy1jU0RaA0VTUpKO
FfoCTX9cXi2ydmNwIYP4tgOFW1jvUuPGEqJ8FzNeLBSWYs7N87Eh36Ar1MoG
PghA9sh4794CZBEKwUtNDSkqf9STyBK6NV/0SQTU+aHQPqkx+Xqm8LU6zZJE
TCb+pJ1OnmtDLDB7mRD2M7uE2tdhrEgzKVw6BubIsT/ouXAQpBnDJTlybYww
EpjCIeBz13Jb54YrJckhYziCco4QUnceqwum7vTcyJDA9OZKtvJpxsuftrxA
80a53uRQtuj5Ct7Ry2xsvtxRgMSynWUzxryx34Tu+aU+hJzjsDMlXZvuKk+7
FVGX52eNWz65U1FxvzzkRYD3dQ6sh5WLOUhJI02SJrUTwsXgOV7avfHkfHYU
rSoqUHC8NqF4OgsRbLdeH9K6X7F9+YfeE8ODqtVmNznRZJfw6kkY+zoi7PHM
2bsD/jcAkbwv5Il9b0mMKrkCpwOCVtKnj7Vn1Rp9YfmcwLXxhE1inFdqIWxP
vcY9Klr51tXDwRXJxkfOtCJWsW1YcWmCCIy9ZMadJVJy9OR6in0ZN+gXpSAE
FjXsPYf4lCQcZZIsRh4/WwLfZnqIgjoG0MBF5OccjPjWNV2TsWi1OxT5JhVT
2m6J6afAVLz/pVdE0MW2xahH1UbH1gyhTRi5BN8E3tSj7y9WWN+lDkNkfQoK
Q2MMWEc8N3B0kJ0OLXnvXTR+6F9WChY2ACCM+6aE9FMgpHIwTnTNtllfrr36
12wSVx26+4CNrqu25A8bVtbDwagn01EaTfwSaEtMv0TVtxZ6mNShXcMwuy8V
+38Tl39LJhnLEDpSHI3QNFtKG9H1a8hnonHIrZUZS5WEniHCONoRSf3fgrxT
pz0B6iX6wuu7wJEfZJYcjR5iuN1bZVuM47NWXGVrx/lN6b0ju26IGNC3gWad
FfdCdY8Fit7Lvu9EwdI7xEn6M4rHpdY4XcJJWZGSzp+oY7PxR06vL6F4GXKR
2kAGLZVBmtgI7VYhTbcFHB/dyLt+8opHHLC6Bu3By0wgd6bFhB3agoZ4BhCJ
EXVGQd9AyDEnWV1+rvjnrV9vOqzkUKLg1OBw3oP9umgzay7DeFk1sX67Vcdu
petsK4ZsIxJZbCYg4vsB4gw1fL7OqtdK0h1Xm25wsgEseQdFlAWgivjqeiDB
BxO6f/Z+523SjQv/3URlvXlIXcG8chEzwc46NLfmxuhtWSKmaeTtxOlLhsDP
k05TjXknzYHJZe8/u91V8qqMyQlH7e0C4OOzWzLld+Bh9OxP44UF54QxflSz
AURb1sX6imWbfk+awypWpVuS5dMQ8R2lcjuhe8SBsAzIL+BBurAcj1jje5/C
IoiE1kSffedqjVPpMfAoQlQo1ZHTg2f1/HI6Ln2pD4FGEjOuZ2zyyY0QxPcW
1T57XU8JLfkc0VS5c8vbVnpvsez/7g0WNWXGlSkxnL12kw0kqBED8zwD57eQ
FzG4r8viXdeuC8PwBWa9z/oMz5CtpawRR+IZK+XUOaFOmR0FLRkTlJXzqoHQ
92hVDsOsgItIMUXu0PIwkBXfytgyx101hiFjGPYkOKFbgdFmgBb5mA7VenlX
956cv7A3JR6gVHiMmwRUAKtvwgp/uuL0cNEOcXLLITCKjUaXGsnG2333cHWk
d/HpzWfOw/UX3XaWuojQ2S+b4whnBB6D858xefxw5OYL8l9ssk/M3tPoHWII
V2P1s8yQ3XfEBGaVn+8XasXdzCvG2iJoVtebvTJwOB0gU1aU6TGI0Wja7fqa
uWW2i5fMLRY3sKc3+6dftZvumUyH9lI=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "sTlVzHE+yhAN9Vt4a+7yJC9Gw9bfBRq6xv9kCe7Ng5psJnHruz9VrHCdetev/ZiPTJdBJQmffKsGhcT8C1xHmtnWp2phLrsA++mCi6ZvsisBHsXsEe07/2w+B8eMNZubT3xnRLX8hyEfcYoWZpsP3M1DFemdUhSKGBtblrC5P70SnbNX6tsPF3y1BZk1iC/CtfkXVJdvvd+neDISHf8HMgQ3zyVqVVLAWr5Qxk5Q0qTmCz2S11Uhb38iPyMZsNmVKcOLkqUtNn44lLSyg2Lbku5JXMC3yfQeGjWysDTWvJ9OqF5rG8q0i2n3qxyZtBXl1OMmDqRqZEM83neNPTTvFj/mJ8jY5t6/Ku1mNuJ9TFqIA1f0CcaVzZUSibQCH+yllsFme5mJHt6vWoqGt+/aIpYvaQ8aA5roPhHemoDFuwXQZQVdmFTK9+JvnaP8d88g9rYkHkh8iFqeN3dr4rMHHt3NeAbwWTcKhWB7skwU4zxi3IefrCeiqKI5aX89H4RuszfBM6itpGFQ+Nhnvr0LtnTMRB9rLOBoLI7B44oerc5yyv06++719Uggsdvm4sUrFTLbGyqcG958GWyQJ5XA2xsrr2buDtse7dTRlylaQuqWAixdujrdkdUFdAN17O6xofgrP3RsOo+1x3EHyNQt4vFIpyGJunGsx9knId5GXMxb2mMVfoD+fP/5lJeWAtDoT/fJrN32rMpqUv7s2lUIhflD0YkYmcf5t0mO0LTLWz/0fvDE4EqXlmYCrJaiXzrPyClOpgKaTdmB5Rwbjysmm4v48d6qfq1OnAxcWxkdbaJDM7bdfHhNg0pwDXm6o6vwoZpBORUFGY1LesZyvVL0dXlwQuWcH8P745z1gcFmqXIL293vrNArH1K6GRy8tJOtP+zaiBYeK68/KLbFm+sy+Y2dCO2RCmnM9VAYSqXGo5CVvBWuFPqa9KjpjbgYUNZi4oNcf9KfoCV1duPlhih0B/CY0tNW9rQS7pmAEh5b+d+ne+3zyG8LiRvmKRsnKpps"
`endif