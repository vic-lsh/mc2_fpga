// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
i9DQhjN+U8Xl8jFaCSJu/SWm/8AwwWSgmecCDoNhvhWAvPK7EWuAeGG3DeAq
5YFJFT/UxFsGLQL2S3uhHMGR/oC4I3et+PBx7Kfrgv2jSCnY0G6Iucvmga7A
OUgQN2QVIWdYN8iAPU4ZRsyIWDagpx7urEvqI9Ee2S7HNaPQXdTFFy4TPkNB
Cuy76jPMkwBZsKL1FbxK+tZI/dR1TMqW/jRe39k1tXZRDBJ/znvGX4sX4ONV
v0te+wStdddH4XYDbEzI69cjYTkJEetUgtyP67xDP7GxEh4jivZAHlesWuOn
DDdAsMkU+WW/HGIzk/C+g1yRgESapC/Aarma1PFDNA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
B2EQglonwr1RbU/g4AevdA6pZ5qNJokM1ZhLDzz7KBpKPKXRMwLCQfmhlumw
wR5XogITO8uofV5NMuUb+yiTjq7TbPtS42Vc5TKZO4DtUCbaUSGjYUk5e8zx
be9809KXSfatimynBqPLm1BmZ6gZqJaiC0iAAQjwb7UjqXiwx1I2zas6gH0n
rlD408Fpp6M5rX0fX25FtayLy8pDtIJByA6yg4g25IezaSNJ3eIB8ddgO9SG
VP4IofkvnmzQqUUQGGNRylw9AJZ+pZrmUmObiCxzzb4oYcJmsw1ZKLqvYQAH
Rv/xAypusSsunV3vjkLRh0DQhjd/VDLChRNbVASOgA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mkl21gGVE80veY5/HwtonklvpFzEYXCmAV3CohA31LSv3l+Lnnyp++IxrmBo
tpPxkf/mwpcSTfvS/0aCneydgxjx4JDnqVeftKVRQlVgPTXsvo6abRqpP/nu
9AxLDzUJU45rsZfUKY+o7k+ennqDI21YV+qWBSzKOTBTLQveRUCCoD2MH9bD
ycX5eXTPWgj1WPOnAKPwttQ8eDJfxJ7JdWBtmjGtU4MRF46KzdWnOZGIDiIy
jBH8W70TpONL1+MZB7xavq7vYmBzr7ghgei/+DaMn/qKZYuf+uzQdeImXyBO
GDLiO9gvBiPlamucxu+qxvYP+K4xzNf/1G4Byv5TDQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VU+bzxPg2SL+v+Il9u+pRXcD/L3cpN3wmef/mAjpEz/J46vwxD9JGrGhg2Xv
B9OYcDKkGNTk48VLL4+V8YhRvOqd32G02EHHDbMF47+WZyVIN4cO2Xi8PDtq
vTu396T//vw3Uz5+O0AKh8QlhrWRsR7snq+tAf0gtztiBrQcCoDRfQYDX8XQ
7DUgJ8WdmvA1V7TJTBXfQZ0K+pWgbmH6aoH8L0RLP1JdLqeGX7sR4zvFmW+l
rELOOsB6B7hm05R7xdRPFYA8/XTr7g34YBEDp1GwinV2+kbnvjzlBGKZYfb9
FdgqNZXwLydokKo9WRdKW+OrGBescvNV11/ZnjRFwA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FxU8IOHoaEEQZlHvttnMbNC5Lfv+jho7ZB1xtDWK0Cp/FrT+osIdVO+0C3/O
RzzCPO1L5KU1z1eSuMGSKw1F8SGqA9jHakG0I7G+9IyXhAkNkkyJvd7jotQt
IO3AMb0NpDP4yEzyWCGcISfFlX6JX7RoHa4HuatEID9eOhGRnVs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
fucplon3T2Dj5vXVJPFqnQxcLNmm+DJSF7j/eS5DHUadAEZKLliG15UOLXcU
CRPJnQAad4ltrqwU5JfVA1njm3PpLCSkvq+tTwAio7/85TUa6lgesL7YmNJo
ffqlzUuCg1zXq3/vW0rInJ63l703HHculhEijs9afejEb/KTRpaMS526FYBC
584xLewg/8cndni/NMWVpTyBl/wyc8WcyXcZt8xTqO4Fu0VJzXqRCzCJwl12
UEPUYuQ100kLH83qDFwFYIFHl2PaIn7YtSFCX0zel5sugtrsJU5fu3maCClj
FvSRtxuFNBVZFFnkw2p+vW2rVDDFsoTVB69tj2pSMjyfreJm1kc60S9LSSHQ
ZLv4VdTxkqVljeB57MKWn8ZLM4M1YuvC2L0U32TrWfwEqD6ynKfnWTybRAhw
sOMykgmI8sTDv3ZtkhCgTh8Lu11Lx/pocTOOuMVTwKKnegDPjGYHTZEBKLnC
hZ2VOZ2Pb3Qnz8njTNvjrZWvJjuUiz1Y


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
c7nHeJ8seBKaouj4glKO/H+GNVmEpfVCtNn7Svc09cX2bmD445qMyTTO5m/b
CPr63XIeYtAQrp/Gh+4SlTw5JAEQGLdT5ppW8UQxcvlKxNzV0Kqm/+olxDXV
Fzygmj3wcbiUYW66mequx1+7ADCES1DyoM1xllV9ypiYFwcusEc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DA1PMocUjEW9g/ipY+qd64i6zxGrwetO+XSRCjXetLbPb+w/hxUCKr2M35XL
EhqCzLlKwqxT+gNmZyOzyfJiXoKBHgrzDW3igXnmEEzcKy2bmaMdkLcsnc2F
s9A74Liko2ypgJRMNFhPLjK+pd7bpM0KUYM37oGXCLB8guA4pII=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 32464)
`pragma protect data_block
a2+dPEfcx9vb4kt969reLdFYLI6x+NeNBXmqsHabuZb68Xz9GjbLu75nfT8F
YEsFkzHjccH9WLqUc6mojlGvWcAxuYCRQE4a/uWKv4y/YGXK0OFth5eP/wtK
TnwfEzsUu+RgH12TxfE/K9oXAp1+Bv0FUAxDIcz/fecEF+2rWn8YuF1Ie16D
yZ4q0xIb9fKKTxtwnzdUP4E+3oxTUgyEAjCrI7catiAw67tavMBWz1RjlZmA
tDLYMsVdh/7IodLCBl03pzoPNT/i5p7YDucOmqescdPRISVnZYKENtA9yxFL
/ExlpOezgHJoYHmWsQhoJPuCPLFH3YxmTlAHGBfM1AUl0lD9olYSUYneGEZ7
P5vxx5PxCP2PT5GnemzJqZbJmNwEpjQk90NMCNHxhefm81fhLCH0c20/N92G
oVhkygd9vYG+cnLyErMFHenFdDc3ctNGKUMgF7KD2wmdfHsAgHO31iYVTVxf
Gh66XcZmHEHZLq+WdGhlM9aIDl29kW0OXtb36xJBX8fwzrJHqBpU0DdSDStt
PKYtCPbR5dk1imMZ9Yohgg1kUW/MV0L98mi/qB3UMFYWYApJpqiZV9L5Ahld
hSa4x2/mheAmkSE4jmAYSN+TDOFgyshDKE8fUB7mRiESKNSQZoAAgyfiosTA
hymhBQ7xaCVNB62jB/QsCiMh2sbZR67DRFDAyBNkukFfkQWc7w4gq4jhTiuV
YBgBPdOROSW0e7lrILrVLq0Qxp9zWVTLutEc+rGeBkUETXJjL9s2ylNuesPy
i7ReOzqIBPhWdh+x4RF25Oj7nmB8hQMHDQWiXTAIfYzteOQCv9CdhSgX+DcN
Ryln8KNzzK2bpqmbsV1RHtLbiUMJS6o+SLJ+WOh+Atq2qTe/I+jJKvMDDGNO
wtWmzRCn+ICBJf/n1Q31JY6yT2i93sHpbVo86VG9ODo6uZL+hYTpcFG/pgRo
1iVvgsYYX6BxLqBIY9GWv3JuNQoZ8+fWtPljB6sqm7oUAqZxaPnREFvrhoHF
+lHiQ4P9ST5EDaYSUC9vuwjiX9kFEky/yGzrHfDQ/F7Sd+YbfvmJK/tHQwp3
X1qpkSZb3V8DUSO68jpTLdVGVqxdwm6N48IMt8MVSvO5C16G/9rW4NGHVSLS
R4wJaoIkHn+eW7sHcskwktciTNGPlhCalcf1RThT06YLqpOVf6RkdIiQEo9r
gH+hSK60G2t4Nx7/DAHFtXZRfhGGuFzzxPuMhaYsJycg9lZAGU+ErCjy6U5X
zC4Ar1AYe1INjb0yj7ccXyNnljq8nd/8/YKprM2PjPM/BfaDJUy1gNRlGO7a
PXPfexEJMI94UJOdJpCfkJk63TXIWJ83Smbfe6o4XSlnYFm/jYvU/oKB9QhF
ZExgkxZkC+Zge9CzTY0FmceJuJ5ikl1EXP1khzvYWM0xfEFbSQ4Ytx5d+kX0
UadWjxxNx/4k6mxl9xe9M866E9nNVWGTft1ehtihc6xCxQHWbesZtCuk0LBk
OEq+aNxOEwSQWpaV9RTMOG5GyV3KBd7v7aL+t2jI/d9DyNfbJoU7g6EBK2Jf
zLZU6B6KhPxDtEo7yDzqUtmE65cg//FmV+1TqFnl26OCethI4IcrFoJGXbJN
Tng6DpWN+nzUrBqmRNpj9/JPKT2f/RJn+tw5hxHrrBQyLOtbNB/uWsTXlE5c
BLM9+Y6gj2WswuLMq2ij+gefpyy1aj11zHHOPuXRq6oGUEuTn7asMKiEoDZP
9CYZR2LOIq+bOVm2cXpazDSTMLBMZiipnlj+/gdpTiNYdxRHD1FbuWZHlwmO
AyMR31HYta9sgEH4c+6eBVlLQWys926lyNkBBbfqef970E5plv8TAv7hPngW
N75W8CHg5rfC4vkGGX7EbQj8fa6mw5GfH4gfSoy2a6dRHiHLofL2CDeCekrJ
MsLMsuINSIlgle48IEQuBzjCtUdeFi8ZS34K+XDnp+VGaIZKuGhb/19G2m0b
QrIyuFDXMpDBZxb6GgXtGsZ9hwYkgGcMTxuT7KzJXEpm5mUBj8ClAnI2Yok2
x+hHR+pPS8bLMg3F5tPohIDialYam3j791DC0Cn1a0M7XGtd1wCmGQKw7Xzv
AQxJ3gYL8tn8UwlcSdbupt3ffJF7P5+bVM1h0Zk0qYExjRjQVbJkLX3UaopE
ax+8AuoZlknFpsXBYlME7Nw6zmE4BkRg6gHHw+6kk6s+ZvhWSshF9SJUZ4gU
x9jJ7l1Ab/PYec5E8vva19jOEllJRElvLSZ5YwYAAGQ6hL2ccyCOH/K5rhXF
p3s15Rn0caYwSrlJT51un/ipcBI6TLp2H9I4OWKPBZznWB5wyvUs+OxyPh+x
lIY5/JfFaU0dLFJBJHzna8PiaOTOktQlG3BsTAs/38XsZp28gU3TPXwEI794
9zPMztQ73BoCAPyEsbtmSkzBbaQCEkxkInRydn/aL22/Kk5Pi3dhCwdX9uNB
wXRTVeHWiKFsdTDy9zAZVzemrwDYJjImfbKdC9tLH+I3i2132A5P2mpP3MLm
1/hYmzmoQqMO891s44u7ry2DLVt9i2VvyMwSkN/BOZBGsPSmcxurUxV0qBrS
rjRIMjDLG+9XEW4iSZp6yGMAeXhjG5vzvrpghSgSdGf78dOfZljgfnudVUKc
CroVCPlnNoqcs7v5KbVjo7d50lIsojtbrF1Ezxz/UIMDy+0P+bdChvsvJhF7
vYJ71JcQ7b1jClSpDWlIzm9js5SQLeCHAsAZ0aE9lGI9+sR5Md6lOALeqPko
B9d+VKF8xagUkPj1qgJz58PyTkxT/w0Fgy8xJlaHrwSKtcGqqwS3+1zTYWG3
oURKwUrARED7nmQ7ChP11Aa9n48vendnygee4RkRl1MIlvZ5m0IAnNeZ2hbC
tuz7uAYTNMkbMjvsJHjl77nBUf7TiFnFtktC8BkQ2xPxMAza6ZWZjVZ3wRYr
svvyGHmF94AAzPptGnX7Q3a/ao9SAgNZJwNhkBzVBs7x5EQA/ZyMxubyEhju
vj0b58O7yivj0KH213ZPeAsDmuU2MVSutBBFDmBwHuGnnYD69bgVkohAybbJ
hE5A6pYRPU1WTxEWjU861d7yYfD8C2KQBxXp8Tr/O3jAi3q+hvQimTpKra9q
FBtmeYCBTDdqTs1rveFtIOl7Ad7DUvpmT/yCvv5CtXRwj+TTiyUpVWdSWUJ/
/YRVis8PJfxkX+UcHwcpMb3pAXE8bapBuFj9WTbUxBUmhn7h1aLIiVDxTKxV
r65rmbzCkRwVEbW733V7Ukbxh6XRJdRBCb+bfxG7dgbvBleImTfQGjY7xLfN
zUrBSYqBsiGP9pClnq8tspprfmCB/VFxIBaa+NU9qlBJ0brlgBX1yp0dbT9j
J5bIldnEe90rIqwaeX2sGY6og5CDgute3dFPoMoIA6R0rx7xDyVoGZed9bTW
gDZaMHljtIf0VXhkiJ2rEM22uzSqwb6nM+Ts9QXVwYHwFHKknhnwrzMuUAeX
FeRRyY480KSGcZmTf+nur7MUSwq9TTiFlVYfM/Z/PCr+FfHJUHwf/LiBQy6b
1AFx1V3nPIkuPJ9fB2eLJvYx66/hZhJt/RH6q6nRCzqmAiIAeBCA8in+T2z+
WDUGDNNFkLPOiIe5An/78aF1bGK8nmnJpmPOsxrM9IEE/5lpu3to8IF/8RJd
gOVesRYCBeKvwHyx3coVGte+QZo53GCSUsZd2l6RVv4MlEWo6Cv0zdbiHMu7
NAmU+KhHcLmsboN7Hp0ZelWaWjr26Z17jALItgwq3qlJbkrN1Fo2z/DcoSMf
vg2vrJnccwxSxIMk6pDF0wf/vBg5KCUp6dUOQvWgVI1AARUao6IoBjw09d0C
Ez4Zk+YpWN86Kk5P2YuOwLLZhGxAexb2p0GVsh+hQv362+DhOe/Joha/eyyV
RcYXc3LEnFA875WvGiAzLjdSXPcRp0DyMuTV15iYNIX5DbLvor8gFZyK5l6b
j6XoOgSvK6N8F+au/IeLxtLab+WacVjLIn70usZ1hQz2J8KSwAxkYcNv9LrW
aKkBnvTi2I3scfiGEdI80Mtj3SXuQMNn28b9XXPsnjI+e+E0Nok/4yxMWVRY
Wz4zIpeifDeHGVsCjTkT20vtY1XqfTqNOOzH/CnDfGTPyfmkbcoQ9C6c7lnH
4+EChzGzvEaxY01wm2EgSGd0YLEbKKjXQgNFc5jaDuBRWLnN0OCSpEvBXFOB
wiMdS5VMoNzCm8WzJ9vCgU03woQdiJdZjRch695rP9THSFEBeKxbr32y+hbs
XAVXkbYAlaciUQ+RAeJDn7mORhh7+Uyhk7SBsmoeyp9uboSV2m9uWqogB56d
Tl8WazTtXdXrU4siyommGOdhlPkDPZETn9rQ+0KqYSGAmE+VYxtVBLWDiH85
TJK6tzaAnNC0Bn/uoOxU1MxcTnyqvr5pivjWqPd+k0OOgT4on9W+CNUz5i33
WwRRJ9D9K36Jnwj0Wh2n1cx3Zq8ulaHjd2/kFPtdyQrPYh5OZN2bIj7MCitt
+jM7527tMJmXaMtnyNAkCLbHjvqeeRNukFfRzTg63fIFA36UIU3miRMonJyA
qKuc2UvEYVlH1Hvh8oocNnXsUwsy0k6XCqZ4Ijloe4pSewmrWWQCM1d5oFTp
DzLHL3uAjDCIsFv4TjX2dafDXXSYCFmyuFlIJPfj5MR5woLfCep02jzz3Bsi
xepYDSrTm2/JPRKfhKZ2KYVVBoC9pl+CiN8FgueWhb4GGHOjBXI8STs4Yfxe
NDxv2Br2zFChiw8gYwmmK7brx73DrhgcGyEqRPojBBRv6xfXkDtQVyfidkfr
IAh/Qo7E5goz/sYJKmwa8iOf8GqKfAO02Bx1otO3TIVoumKljG1c40CSpFwu
rxPKEv4/cVfG3i+wG1oC8wKQEfWJETiiawzsp0UlsOLKjzx4ob0Tp6yDXMs/
mc359nZr9MJjI4h5oPVVCarh+T5oG3euiBqc5BdOuZ2ke6ECbVgGg7jMkFIc
JEVMO+HDizMhs0WXy0I8z/ybnXQe4MNd/8EBuc8CrhbqwRuyGZN2J7w/gkZC
Uz73nDf/MxjCKjIt4eF57NEMnxunwbz9nwq8PHoJqUopFVHWdSm40fVh3D3X
/K0TFHaI6w9yAOk2d79kjJMdyiIuzxSgfIfkXZy9t50gsTTiKAE+V2UJZoE4
ukb4Tnd+cmkhxQ2cBhcuO9g9BkQy9JpwDbhAxZ3hyec6Xowi3wwJTc2oSOwE
bJVHt1hGzIYQzBYOnYkUVhw7T2B3tZfg/WyyM7bTS9JeUZyL/nnj6yFQWGA2
X0I9dh2LtRNKtk0/Wy/DGpU1k2snlowyilCuBXcfK5/3ZXKcgy1gH8RY6KOD
vLHVVyUCl7WqUpabxwahSi/zeA7d5jEVtxrEBVOVnU1fMjvmwRQQ65UdE+fB
OrFnJwlufYBQ4MvdlOoU/sUUrqQJdhysMX73w8phc2mYFexaKN9jY32RCmHa
jT6LUBK4BvBHv5qG7efOUC8uaelrAdPEGOldahIWFaD8jbpCOUI+0k+1VMHm
RCnTUtDoASeK0+5/tXHvuE0wiVWSghSknoIhT+CctZRB7/jgbY73zLnHRB3W
jAKO/RsCbFC14xIiogBymrcl2+Lo0hk2C06LHelbBLkqm7UQKm/vonoIwDtF
o3BXBe+twUkqHw9GWjCZIDiY8vdmFrIs0+BI5lnZ9hWOVb9tHEZY7+wLcC67
TXvIpVqdEopBt6lpoTrLyovSebp/HpMJRlbKboCwXzqh9swNhzFqW+LLIOnA
NLMCMCVWX0s+hr2A/iZni2N2OCikcfGx+mh+iwJeIfBFK3249tnGO38UnkW8
L/3Y5zEg9HwX/UPUGk2hvZ7mot1qEEeEIF8TaQO1q4m9CxOh2l0APfAHAGF8
iRutB4MxpSKSvpi3+ReWfPlmvs0BA1kvn7M5fM+H5PJwCVI3/VMsgAxuGSMg
nk4Y5lyov9sTiFVnImUb0whzvUkIqoV3kBh8jYAkSf7c/zvSB3VIAzX6RWZu
7cpJqcdh1gcgh0tdW8YyUUbS+6kwzZTMaUIcJMlpQ8NIzvVUIKCsWtTOmhzr
TSoety+mFBgpYlNK86KOEy3Yl2jpTzRp66/g6Bq47pgZOYrbPqmoMue10UXP
UNX9iGGX2InibYdBvxFdpz1CMqzQDIZVkZqeRZ8eOqaXxl3g9n+O9prfTL0q
AiUjctqHcn8HDytF3WoMdRarvd/VspfYRAcdDgwkblsIWwRCJ817vFiNdOkR
/JkvQ3kYMOmYywVpq53gYWAikIM+ylWHyXkhnfNkV+Sm/oIMyqs1EkkdSfJS
kpZ+7OpzszuxFBYE1ghf+afXog/ymd288s9KReFXFQM8OcFDcUYQoefKJ5Xs
HtKh/n43DYCbfoS0noa6A6JG+a8kupfqfYJ8HvPog+gpY4Uucwz6/5Sq/YDg
KgblL/8AHVed8Rd03K6C5VqtpaIBqoR0xskILR6jjb3OEa52lIV54C7atSkW
vC6hceWCVT3ceCEPUQ4nlDyFkZgCG1ZY6NRPjEWHI+Be/hAwtKWUAOi8zhUy
W59UE1ZI4PqFVOgvcQxLAi3M3P4zHst8vFzWlm8QAj/TOTUobf9q0jnthzjb
6BGECZIyeJyQ0uqX41ey8WH3AuoDq15YzXrW0xsVUP5CF6KcbFSl9ZZm5CB4
XQpxK0lVD+57hQtKerl+EhZUymWVNewyEA2C0sr/h+JjxZFkAsnI92hfvwLT
MCFYOhbM5Xyimz7hZVk2LwTSb3yim8o7518ycVA+lDzteUBnecgh0FjO/hNP
S8WU6H5Xi9frvdYv9hlAwj50orCnYSZkIrPPQzqj/D25omDdEY0+gNSjytJc
Xa1AB6GZZnGwp9kKTFpr/3E4IJfFh0zyr9DghxrDJqpr/JghbmlpJRTgyvTM
8dRZWVrwMehTGdZ5BBaSBVKi7Eya6VF+KjrI0jBQYfVmwgNs977wh5PQKr2K
JPh7a/nLLUGEr2s8e3GdcU5sUhN8Z7UIK26WQVZfWhTP1HO6Fbml11l6CXmZ
PuwfId964jUCiHNCODei713p9GjQ2tZ6jH4LC+k7i+GNBqkZ/ylZ02a7us+f
e1Fx5zsCZwiLQMSwNSXyK7neUlzCSK2fiERR+k4ioMYX/a7s+D/CjJFwY8Pz
117Lgf7pKp/uE/ilOKXb9tyxOtlHBgCeoVyxCW+O3xozWQ42bxtB6VguE4VQ
gDqBEV1zkJwXuXBA6gV/hX7e1WNqw2aBQ+kv+IhL9zwyW6nDaNPybxDZeQ3W
EyM8HGvHwfinIbBTNkbad6KeOwG+qOFhuJhu3B64EHOnWA9/wD96H7JpZdYs
pl4BT+qwPrShQTTaB06zaX41JzfczURNspLDHh7PbOd8fqsXs8+kWNl615/r
6lN9mlLtXx7cmLKfDZWSCNKIhAvIWm+z299x99q4qXUp+9ZtqNYXkvuY5JZs
0TUIU1ocxshunRl1srhLaIHrXmDpfKOGHhyvy9OTUEqz/80dd6P/QCVyAQtq
eT9pc5yIfFqDttQNYxqWDghZOl3cdMutxtsTlXO78nuT8XGFVKhEo40qeq2I
gu/BxpMqj9ddY/uhU3N719y3MV7d3gq7DqUDHRKhEZoSPNvOpz53xjJidv8y
zALCcsg9hmGLGXyPaJuEZt4PmyksbbcHj43XfLqGBEpg0Fj8YjmtqA1w/Ggn
rYHPBecvZSx6v+Z3WiL7Slzk6ygP7oL602NaHzqIYV1/kLNcH/5qEuEbSiA5
7ws4Iz8WTd1by54ZAKCLg10tKD7U3/zf2uH7BP/pAhEufy8iRogcmi7/zu2s
vR1mRhVO0m3jTBPaEqEvpZXjhxhshUPW+fq0qAFxImJN5RMsNEItVwXQ2cZe
k+Kz2XptjeidAdWFxvB5LEXXC0loIOfsT8mzWG2Q5KDtRQPxXgSeKRg/Zxbu
RbLciMd+vDROyxZ/4KlYfzrDQZ0s/asVeRZfpxRNguSJ5lntFhhtszLlfepj
OCa+8PM/FfJrRGeNPkjsNS6Z+U8b6GRcnfBxwRHegS8Su3Swy0+pmq5WkiT+
v8rhiV4zU2rMjjg9RdI//Hah1BzdDWA780hJuLkSVjn9gdYBmJb4DCYerTCi
m6/doZqWNlePYV5Gsufwh/2hzUAvWmmc2zasEsYaJqGTwD4tK9NeQ2QnFUjY
pALbS4lFptKSmipzborSa2z16AapgSMJASevTAVHxcQZ1wnn5rCZnvvUtOsR
VrTKVqeqZs1bnH2CrSpL9wrBYMggQmLOtWMWAWsNB2yvJAT9jmsClnK76eXz
DPxuc90gbfVpeo3MrBfvy18J2L2WAUeXwwwiC4t0q+/XbzU14aWUN4wvkNqH
N3z8ZyAEOSqfGInkfgpNVwwhMTzrEszfwHSk7wfJ6Jfs1aqGFHWxOWCbqTE1
h9e6mrawtpFcpDMHDb2HCtNPyCS19lZ3U1AZU82PaRn2zatHROJC/GuGtBYL
lP1oQbZBRKhKYd9d4YQkgN96qY+KkfV+yzQJVplyx2CK8VJ568Hf4t1GL6YD
TvYdIfJe/hdrBnTvgroM73tsTt8EyHPQ1HKEZ1+oXGorow9FVgcPYqxhWB23
6LfKysYEM+JRLnKfiygjwliFdRzY8bc7nzRywEZ2nOBUlk6E1bqUjh6MlNPw
UIdayBKNazryVsYmk/HFOxGVk/aUGLR49YHnL2K26plTDvi39OPspFMM993U
+iJ/2e5RnZ1vOk18taOAcqCCsYbh6+NdXtjTpjCbjNKqoCzenDl9QoTNgaj1
4vSOkz82xhl5wOlCuJkCh1WZBF7Pv//afpB8QY4EK7XEkF5tTT/S+qN/hzNC
MArnWLPXXz3NrLVg9unBq9Ajh+JPZXHtto36pdZNJlMDgrkvZ4fK0/pA87dh
YTHjXT/PhqWqUipdew7xmXJa5zUWvFu1Rz/7KSg9mRRcYOZdXW/TVWUK+LfQ
w15Iu48rlZ45k83FBWhOqQhKLBel88jd/LAQNT9i9LtbC7wk44/GjswHagZ4
TmVl6z8GrtZVPM0fAYHwEk31wfDgpxTJ3dm51olDK8u2eknr2q8bq4d8unQG
/IysQrqDNJmu/FRTMc8ZoRh6oWUA8CxvkkC7jfIwDQ5NkoLERgJi8l2vaC2g
DYbjOUacs8d4Ihct674swbHiwukr5aAhmx3VsXLlYVI2XwsGb6APQEMFI98e
3iaJd28UIv1AAmPM4S7Yb0nFOQYrxqG5/nlrKIJKLZn3vQsYtLoYMGvYfwxv
5msa10FMJRhZN6yK4x/8UCthQuT0yq7toLFEfSc8DvdWo37cg4ruAJRxst/f
feeiorU4dGWcf/oEDib3s9c/N3Craoj1OTqq0fyQxz/6hBuw8XUTRf4+wuP/
0FTbv1/c/0cN7skng5zZShPGjWcFCz3iRAnb07zXM8zWS1+Gp1Ls+qhnZom2
mJClsM+4oP5wR6sATcV8Xsmf2gUjiVTi+9bAJ3ZLA0WOxVnWZSsCwH4KfekD
WvilAVGn6hXn5U5TGriFv9h/dhSawN8PxaHHZh3rJBMkcKLm0TBTlDy+1rFQ
8BFg90gBD0xCgax6IxkDrX3uv8bOrdXCOI6GjefM5VlNmnchYb4o+NLfFwxJ
4SHFazfqObgOa/xl4YlYi48vEZbnSOw9EkCrJIAjVigkKAhEasmFATn697KH
MJ5xdTq/zQT+AWUqa9a5AgIyEaWnXwo0981vNf0mwA2w4r5huRxDdxyD1W0f
zpVDALW9orjO+8NiudGXQVIfHLxqYpiklYADOr0jEQq23rdpjc+kNNE5IfLz
4Lp2pb8gTw33VsepmPwQngRkYWmECFqiST8npfOdq/JCZe4JnSYWzwv4LytX
KQgEuV5C3bNbifo3mVibMD5ec1gOZHhg5ZbR/rfgiq3IH0PO5+j4HLigaCLB
8wVB6cbSUnNCtQiarRyvg87lKZObmL7RPuG4hGyY6woyGXB4RNwui6d1WAiY
sFlcByA3K/ZhKPGn4re/DtsDm+5Y6GkZsQsg1X6aRNQB6d2eU0YuaY12MI8d
fPvhN4OIz1AcNhCLBnOGv8+xsZYKs/hI5TENja0ub6zZh0rnu720pE29GUfn
PCCZ2cm9ZhbdSYEkPUaJMdro+wd48ByUGNv07MO/Z4B8JzmRnEQv8jcm8zjs
zDnlsEzNP8XxsMOTJicGBO3PV/WAOjffYBbwbgduE56zUFD1ueG91QAN7Ul8
YV/ILW/ePQEYobUaUNXMbhTZQxTe7vXsq6Q7M57SWnMbtg/mlsDYmxH9jH2T
EAgxqEO82MP6uly6HY2MFd97Ptza7n+j2s8wGrHifpohfr8p+nevRYbr90JN
GjGFyk6oKp5RHCWWfU5WoJmo3izostFTjFtSyKEAQ3bJHxvQk1RTtYD4g9TH
aOKjJZ0m5Z81hhZgHJG62eZjvBwzWixKz2fSMbQn1oVF4SAeZhPaBe7FpplB
65lm4I1W557HBYvGnGhpBBNay4s7yYyDtNdPTWxc5p9eF1v0PvBuA1N3PzUM
jCOJeCfCm4RCwXMW68cYzFza23OtDQQdYgv2J5Gi7a30CNgmtdOlAR+HB30T
pH3zLYGLaaygsuxyRQ0zkN3W4p7WvNSmZ9l4oo2DBeeCbzaoxm5KC+cpLFKY
vuyzZQQ/SWvqUAyHoONpm22X9TfQrZ5hJrsNJ0CzVPOyjpVkxXJrXrnPCnxJ
esj675nBNxbU8hnELLq2UWORJuWadhxSWAt+3kHp5qWYq+XwDx8doq+dGtMW
748EfxIwu/FBBN8SN3I7wXBrufFQvG6tP3SP98b/x00H+0TZPJipdpPMrv1Q
inEYCaYaT1Rz8fZ1oOmU2nPUvaQYo61dV4Ls+3QkfD1L6VHxqgeRgNMMpfvd
uYulsOf3da/GDUpBWLna2/j1mSvhPrURh3XIkSH7uiiXdNGruoXbQNtYUjwY
/M9GQ4wEBXI2FDAcvLETxEymmPN/NQzZk6WHTRtOzo7CFYYI4shUP5C5+mFe
mD9iPX2PopdtGh8qASaU5l/IGUoSuyyWrBQprRx3kauyzvnb6CL+n9oZJcjT
c3gLb1UrM2ZNwyPiD4ceH7RLRGLcpHrE8cAqcDK2AC+hHvo/TyebitxaEFW8
iPuVf9Q7hIzeKJQ5yI3D+X6L4gARbxacddXSMbx3+IdTtEXiQqQT+aYlPqRk
h+jvP/UCfA6O27ffDOsq5cPFyDvZJpB8b6vMRiRbg4XWRVud+0wgmolGkSPm
+kcYUryjLKQs0E9uWRQn6zX0Lul0mW2H7SDxayAfJarWQzMTzUc3Ry1j4XLc
4IgF4XvW6WyxUJXa+ipZjtYdwE4p2mm2vLAW9hqS+WxwcOc57TlTMp4Fvrny
f2/+Nada+KZNi5XcmyBLjAJ1uXKrzwMEAhoZeJNUKoROdVWEnQD4G6CU16ds
bzbyvzyFjLV+8MENCCpcQEW/aWo5cpGitdFZScrzBEpv5m/Zw/MnEm+wyvaY
k2gfUdWk9NwkRoSmyH9jHy/jbXrBRokav41OR01UoscApD9u8QQCH/z66WDo
u8uILhSI5giZtFUzN4MkNzaY2YuZZyB+d9PBMFX8BMk+Ep5BrmoC8OJTwA0o
n3rxqMowAJXHU8aHS2Z31aV0sS6kgqLKskqK7OukIUdZolgZ2JYu+bMMKhVk
R2JT+9peFSYc+3rrC5byljDTOFv2//WmEKVjGa6h1OZSX/thiwk8zjvKXg4T
mQo1tUzke6+IiPRXM7z1JDn/3pOuEqnUl8GmAxJLHIvPWkZEeBoNFGnoANcs
pJRaL7Jsy8yIajy1NHtSwLV1axpuOpJ6CqqTn4a2akwsaWQTMAYmjAcc7UeH
/0vB7w0xZF84Dzq7D0lv5gazshmDkukN8QtrjjcsUKQdhc369gLHDIng9OT0
WyseSjGsvKKCcfg5vzcP0sMoKM2i2T5gMhI7Xt3/34jF0CqXL2tZf5dOTcCk
iBn5uFlxNJOwiYBGZW+cJCryH8M22v+GEgbm5/9UZrwBggVKWGdd57jjZSgX
J8d2lhcgwJT7iZljB1Oyd8DPLP90zoRpBCI1yYrT/PQDRAtcvSdThX2S/MKA
G6BTpawP1yUf734mAoBW/nuPz3ftel98AmSV6pg8LGN0Ok/7bp26LrUTYkPE
tWXZRtTPvpoHlwwbcFOB6OiGGrL58ugEyze9Nd1fw4KO9pHU2v+vPh7mGKbJ
tLxlNDzkPuCm/qPjFluo4ro/Yw/OVRHYy/OiMacHvecCwx5xxEsBuPfogpFp
UxPa7echbWT66WYigw1Tl0x0J/ykV3kZhudR1xonjCcRqmXvYGxYSBjTFzUc
Ua19c1fsDL0py11ZEW3tZmSewI2qpe5BLpuoIkQQi7zqpSHE9B9iAJbgbwq3
2W+l2GNagpgFaBwjSJK3qu/CIlypLcCge6d2fzz5pXrDUnUlxzD2Rws5Kowt
UlLud7bQW8hS2HoK0vnIUPYD9UIyHpnGRlWsZG/yUDPxGApguH944wlFawZz
RFBhwaR50pCVTT5QQlj3QAbJzy1OqzaP6MtViHKQrfegwhRI0JqGcdH/zUvg
j1w5KkhjIEBZL9M60UnGa7/g6Yx5ua5e0RW+ofCi7Z0iAApH6zwTWSpT5n2K
fIG8a2071E+wndRgoJn3KOsppnbYdvnt8efvdYFJVIxwB5Lh9aKQoudhSkqv
5AAHmp2UrRfM3AzmN/mInVP34B3ZONd8/p8dSkkQUyGCBUZc0kxg4o6dnx0k
1Ts7Mh42Lmoij/XtGZlHzyOLECINhE4R94DZ952sWu7Crpj/8dcGGh/eay0W
Cpl/ZVBQRA36nWD0xPru4ZGeoeZcI1yZbmWJ91DdlUylIxKllBJzSekRcNk5
smAtJRU1X6KA3AGoZRltbigkXMw6yIRGwp5omDyYqhyjGqaarmNitVxDsi3v
N45Omrpg79uIDo6kXIXHItVL6F100EQW2PQYpA53LlfpqGWbJfHCKJmxBoiN
mzu0841dOxI5pdUOajP2OmJWAH+3NINTv8Ck9R+ODF8M7YWVRLg00JP1lW0L
gIOW8gmT9pwnzzvFUvabGdDwQH2gbUeCAftfObq/ZjNJrlzmXipJ2YaQ7TdQ
6lU9zePPD3lh7+akhsGzKW83WrT/gSjRur4Rp+YbJDZJRYFsGxumEKCNJ+5d
Mupo8UJ3ro3zSfkb+MWCa50m/6djb7zKliHV3uelqiJMg/Z6DmdkkwQIWVBA
wJraaQ2chw4D2biDSO53NCagktak60zqXdVj+i6cjR8Bc3XjixtK8HOLRDpG
n7fVTXnvrTnDA7NObzKSa33ZsZzPEVqaUsUYmU98SVtxaoaO2N2Mydm5xQSN
O5QKbsMytw4kzVn4+ezhv6uVgWLLG65K/+Vagw2ftnnT8/XAV4uDIX7kevzi
qWWVKWn2HUoqgb/Q7ufav+fgFiXuTPcO46bNGIcMXuEzHSH6vVt0ppKqxTER
8jd44n2KDS1FHR3uZtbAhdGzJEBs3pPs6wSPSDh9eiJmp3hXHBtk77Wp7h/K
vVNNXl7d5/lvWlanf04p/PuMcfVsYRFtLSLXxVOVvj5F6Xaq+lafFvg++YLL
Ii9NoFH9o43qPIUdick4QAaxQKNm5wOhjsQomgBCFu1xP9QP7doyEYVUVOdf
VD8M3naaoaDHm7lZlisr3St6OjRzNSZAwRux5HD9aY+BgrYEJe6AqFDreNlV
nDKjl8iyzYvbacjCgiAoouAVSWEBbdAgtBW7zAIebJBOUoEDeYhAesJvceVZ
4TQVxMtlvCzXFdQsvG1Kh6fhZFDVpp8jRURHD69gWbuD+KXSAKQXmS4TIzye
ecZBtkdDuXrMiq0/MINpE9NhRFVjPUEbs5yDF3cWy1wxnxS3X7rhoAVHnmvI
ZLNzYEaRjokfy1W+yMJoTxtYepYa2G03ubh6RXH59nM3y2z/YQGpuZ7PNlNy
rY6a4uBcdn6RHknwbB5I/aa+2YdT/yd25GkL6WsX/eOc53rBTWIwBV3SfZhJ
lnEDuDcmOcvaPOWBPvyXx2lFh9X5puJXcac4pWK5IU7/JnCrIPmnV1IYao5j
RTZRCkIVt93Ja9OWc06QTfqw1OALD8NvJuM/vMCc04ejJhXYm3Snos86Cqju
VFL/Lh1Fhk19lzmIG5ZhX0p8ryDEQl1ccQ328ZewAFBRIj3I5i++MxvRAdNQ
fW8u0hkbYSnOQFpnD59kl5eJAD89MMH0iz7kuzWydf1H0e+TByJ10gFKMyjA
uiaLeDKbTBOIFgkeGBgsT0GCdXr/vy+yT6vGSqlkq1oBvLPRtxMXvJXlS+ty
7PKTTUBzJ6L0ADBTG+f3jguum7H11Dy8s9AOe0jpEBdQSLl7Yw6NTYEE441a
l5Bz0b8Fva35QVl8ZHewqBx7ODLmYyKxlCudAG7QB43SehWgjN+UhmbhMqMd
dkINZFSgfmb5AK0CQElBkBZFRWeN/GKWvh6mod9hNPe58DMGS32Ou7U0YuVQ
a3p++FnpSIXGHAQFbNWdQvTJQzUb3raPOt63TWtHWZDlS1XWz/yuCXRUlqeO
l3yHwtpxi4zanvYh7mxuKEgNNYLnFqLkGZdjMLYgMaKwTOz9mAtAmB2EQKiO
ZZJNMg+cOLF/utbrXqZWE3BYEcLsLPqL5DAEC24FR8g9ST6Z2yXb7ZwStW6F
uljLFue4xFFb3T+TRzw/PJtgWszJ6T8enYe6XQMwvFImF0mZN86CQhsOjlM7
3miVys/RE0Q/DiqJemtuC7I1md/7UHQeOWuv0n7F+r6hQ2znJVjYyQbdCJuV
LfOtzB+90Anc8sDHFLn5p3Q1RRdeZhb1M9MJ1M3n4BDA6S0wO7ciRVA+3JdA
xH+RaegbfK0rOqWoLxtEdah8rtBiaEhY+u4Kq6rLPnoj+D9wLeTkWGlq/gml
KSUQu8OAZlacNOKN0pOfDM6ZIjZ7VPu4xNd/zwlgNZUonGTkGeZ4Da1pMkOM
OBdeNgrmhlM5w/9ecEvUIPx4/mWuK+pWoFGcqbOvFuyscCyeA+TE6nV3JWjW
oFqlGejRzn7ZGvjSP+0FM3o3vN6VCY5p4quWX33kb0Djriy5OFGAEE5wRUdQ
HHs+TEdFR+/qTALP8hqGSeHm5p1K9IWm2aKBfhXAOJo/1RX6dpm7mZxHX/4K
1COW6RQPne9Pwt9GNo2EWD8jD5yvTryNjfdIcG/hpkmRQNnUtTbcQGd1icFM
L9mVRSn6pQ9nDHwJkCFvaNGUw9ZkfMUOKQoUMWxQmB3rGKuDQLvRVKPzCJvv
HKXaVdcoXCNA4gPwto28dMQKKrvNx5/Pab7gjTPBAsNFPJiG6gmG0hPr+Gjz
noFJwaqU1U9ft9lrS3bayBXpelKIXeYY/aAK5gH/onMt/JpcF3NUb4IFQXpU
ySJhLvEqr7DW7w5ekBuYZ0tneP6sVCH093qCY52qSlarbikPtfYbhzx2wYMy
yTLyOzGGrSYoQkcRs6I5l4mSDjzQyj+oc9dPyB+FHMeG3ZiPUuifa7+kZSvl
Xqadqs6KgBy+CpRiLFcytGpgx1YtHEQOijF+bI6W3wVw7jzGyP7VYkGDi52w
laVt7MgD16+BZx5tJMTdhQWA026vbiprNKDfSWe/uxsblfAtFOhJpH3pVCCL
92xi/3G72qjWyOPlnz3ynlbUKo8XdDf2Mn0ePBR945jeUWt+O5EViOPQwUO+
srTznAExaePASOz+J2nd1Y0ghNQmtRzWhBGlR3qfA7d+i2zdi+7QQSOjmTbo
0Pr/N1HcxMoRKTwYgj7woYp1f361sp6AbA7oQhaGrWFwT+WcZFPaSB9VScpD
M1i6vJG0LNv2+kKHvltu/8jPf++m64Rj8BO1XxeU8Q+ARLt3F0vsdheG/Pb4
BTPb5OxLmNM+KUioxcNo0YXm5rEeA8brk+GmKTG+4q2RjhAWX4ne1UVXk6HD
Hcb8y/7Ixqa725SkInaWQqGoUkyi5wX9rfY5AiXw04pWy4XnPOdZzO4ojex9
qxUQNAp7hBk07848/zt1uajlqhHLqAU1OPiRZQAzwK6qJ8ed9BoI1WW4ekYa
JIFER020omPkc1B4iEFc1kVtMFjjVtI7pcUiSPi7ecrQWGt/ljVXvU9C3WRV
1Xn7ggZt+up8ZyrOvyWC/Cq69tTvjtVsKR0JkkLaJC+XkAAUQMq0AtEagnO5
vdcQ3astF9WjNVYHTnV5ogYLXvSoWzvtaaId7PVci3zrJvevt8bstYvYyoF7
UVHyNz3sOdm4H6+tZpqUQKr+7piOCUuqkSTg+gEpv6k5O3smor75Zuy/pG/Q
F0oQ9EH3se4wYnWwaf3U3rDS9wh8wh0+usCePOdsWSNN8qV1nn2s4cZaQAmL
dryotR67SUOmuJPsoeqA5oyS4bHZrRAelPHykN97JRnZ9mqmLooH3Tn/3Mtt
RWKMJwPNpUmNJoASBJElvVGLwqZGiqEEZUu5mpNmm5cFMsGFJ3FgqwbbsQD0
0LRHmjx0ce9FQ4xTwxm0wdSKrWf4gqTCF4e6+xKfRNoWK/8GSXaHBAKhMPXL
dGIvyS6eQxxIY57+EejXDx3FJzr3AaauFrIJeE6joglr1aPZ3COxLJ94IzmS
Q6IASDSv7jJzXI1xycr9h9erFe1tqsXfCmAFuwRHAeI+BwH/eI1brjkVhZCs
x6kSaOjeZczT0loOqHAHt1Y49JsWTe/MOfc+kGXYvokt742FCy9EtxFqw8oc
/O0ZRGZxyYP7rCuwWYtkQbQg98BXP6s0eSrFvxOWqk/GJbeNQ4u/OyNvte1V
b0AxO/O7+qeZvy4+sVLqB7fx7vRN3wz0XMzVPokuEh5xCy0woaDsJ+/iJ1+3
E7BwItLNWvVkHnAb7/0XAMdvF9ELegvbhhXkraMbnBm3wsW7GQCh+tf0v1YD
FWhra5x6mgC+rTdNL59ndEKiBYhUD9o0RTZ98tKc0+0UL37KTpKsvLAsCXNs
YqqIKqDo+Pfcn3AWa87uS8IFW47D2xYiR/ezoRmgPUUoV3VCg0R9mmGTcAgF
zWhrRvnp/Bm4o5PxWie8GqryD8A0cYWVsIc3JbRFqHOxJ7BflC2YJgdbBwlN
2RFNFFXW3i+coXgqRXbUp3ZOnz/GjSkdny2t2SJoj9efD7XvkSRQGZxUIrqu
bnPZdZPktvjnLJLifsun+R7Cw4EzGuRavT/qsv7FxcIW+XwQSIXVVTwzSgqw
J1neV8/jxMTCNqh9j+7pmw6Amtjj+JFJPnoQzizIT7sgh66W30guWWdXHrQF
Kmf4ddPMK9EwrnF5S4mMXtlD0QpQ3Sb6YRioSCbWxToJOFrdLwWHa46wTVL0
53TkAsdXD1v6iHcqTkriPfnJYqinwf88zJHG4lNceFCqago1axZbm1JKNur1
xy6nlUMe3BJADiV7+4coGR7RcSWiW6GpLBmYtMMhFfZSNTloTuokbypgXixJ
znaRWRQXfjLm94ygrkYR1wtNcC7IX2biLN6PncF/v1kZFJNEcW4VWG02y0V/
RJeG2r1w1TRb/1H9rr3WQGWAeoXIL29kVrXxVmPFC2/j10giKUAyPqY6SV3B
jwxsKpSCp1m/x5kGf0xdwSA9drx8WhESRR+0eNHYSuZCAiGb5e8WwXKu9LUO
eQLg8C0Qsuqj0GJOlkGU82aU9N3usJD4tOTLHbvUl+F+w7L06bvdnh2bU8WK
l+1A9xzAd3hzPuq2oRbxURbC0h3xceRb9ubhfdO3CKMxB+kqx4+Q0SFqm8di
t9vSOb4zdPZvVvRhkSVt04g9+tfSErJm9iT4BB9rtGyec88or2WiAJ0lY8FQ
1VGLGMF18B+Dj9hwXBM+OxDaLjjMAQFmLXoLmsMQUipRsioUtGfrhZqCp8vM
Z9ucoRkDq+47UxxgWRWe4yttf6+GzNbBwENYZs0/IKt+pDhJ48sgWlxcav1U
cC67KPoGEWyVERiNbD15EKtJsPrjjhL4gDnTyG/N43XjSEeuUzDAbWgSYJs0
mCmSwgtwnSqPcPZ/IwXN97QM4o3cJZLI/6kwSYJGH/PvHQPhJfbcwMqab0JG
wyT8qnGHURQKlFIen/DqMHynxb1XzMLVT+oVGsqfsBp4G+BKR98gumm8YnAi
8KJfyeAtGtPVXjK6kqswHLrzJS2UKEtiO4i74QZcW7oKlJ+HmNnFRmkmu/ut
aFvjpYSe0pajAdMywGR8GjH074n4S5eRq3g83XQFmO9zKnE+URs3iZ0zZIJq
IRLVfmNOX0mDduIrMR8Vilom3AgU1mDKGH5ROi7JmWEoXD4pv2AOemq3zBxt
1mGcYcjT/WvP+YhbowYjShDDKMwIWeZ9Z/7uI4haeLohMd+TAGpJ3V24xiKk
umOt2Ce5jQXiaOE6s/dlKQzIyYnqoBEDidO2hxVDih9gHIwS7J2zvCjtfllG
smIr/QvgG5fM80hT4nvvTeTRRBuZQ+2dObrYGv2Ol1kTVmOxKHyMtc8qiOWx
iUd880M2Ef0aeVmwmc0kM2N3OnZnagrCLnVlhT4DPssCSfKyFdBIT/bLjQEP
guzShv7F27G6cpuecPAj9bxBAs+swMtiD5zDgO750x5X8fS8tjBtdesZn/1O
2a32pSHSCuHvLpY7mQ27NeEczM/wfV2QxbmnZUKGrciUqnNSYoFDX/GTMpM0
0PsZfuB9tz7KKDGpBqzQ03ninCUDUYZHQsVyiNhzfI7j/SeiGMHrCwat9ZvA
uz26FiC3TDLfeBMvGYu/qXI6ei0+6R/KXW+Zm6oXhYY32uwrKr3XQwmiBe2l
PFUuQuoEh8JtydVTASkAVnMK/sT7llkQzqPErj7HSBrL+oXwARZmhyaqdG8W
wX8YWiSzr0NvH2g2xPvvjApK5k4K2MG0sVT1A6/jo0GpSCftPEYgkJNlvaGc
YaiQq1owdJb8q5C8R3OD7C9FIme3VQXmwxOOMFoGAF6Orxrlj8QSKdX30z9g
/sbGir16imkpJt9Tj9t0yA5XXKsyxsXD2ejMott1As4eyn5EBgeEWOHCp2O/
ZMTrs0EcdXz6a/3eLuLDRcXmJ8Y1BEkc1XmWL8OlObVgmamXYKMii4rG/bHZ
o8l4yoBz5KkiUp80RWzuymI6QmM584IovHJ13qDWWH07oit2gUciiP2VoF1t
i4uexu1OA4q3b0tF2JGVExoB34B56VnAZymtNDHfEEijOSfRxkwnQxCxj6Qg
vVg+tZ23pukv1giyUbuvrF4GR/CwkSFyfZlgyWoQGOC8SoGp8zgmXHvONw1l
noV14lki8nlO7BbUc/G2KihfZ3rZR2ShQm8Hccxa4CRyMZpjM8an+6/DfbZG
rDDR94ulzrLSnLduXBJITXUXYQ7TL6xJQcBhREzAWF/0ixs01tjE+27LdfLQ
xy8YlnUZRUFSaEgw24H8ifnRoFuSzAU0Gvi7hd2XoDbbv5VKVQz0FQcVU6zi
YQWuC68oRw1XiT5bqmnIeqhH/7bQNLo/JMDLMl2Sfjek4w+XIthqL1svCAWv
hgxj0TypSTdZCWvAFHjoVBIMfsOgeS55Th/W52zXyLCVlW5LiPXBwZGoitY7
ZlGLIAQ8MEAFO556W46i42JY35mjggnA8bJmRJlXy2jRVl0JK3KOpuYcHX8h
mgs9ZzKNlcGlL8HKoJMAE0JQ9tthH7va1dR6iXfWm+YJp3mdYNdOXHXXgKac
iUlt74TQVmLGXj7lvNgXnziXvSdiXPmPU79b8uYCWJUtHfjEiCG8AfyyThDY
RlA3Mnyy+hNpMM502rI9VxHfFYAp9EHVizBdSrlFuBjbyPVTIFYL9hW1N6Bp
A/VbLA6oCWskw8rAmIA7BhzX1Kzc++kmQAV0NVg/Ts2CPTTwJ7tLO+TKB7/x
Bv4eYLsx7myetoHSXNk6ZjL9JXfVPLVxQrmZUjQ4rBOEFPJ/jHe68oq4q13c
EmwzgJHf2I+A3Y3jG1cd2Lr6xxmZ/NyUHvu7p3oS9J0MZCJrrQPV5UWrtD6v
EHN+4dFveq85UuWKP+fGLeRwlA8EBdkSdcbsbyqFdeVvhlnmDIbrua0xRUyF
lFnE/9fzLxuO4qp1loZop6RnlJ67VAdSfuU/SBjg2ZxYYCekgiNSrC+J7jqJ
nzd8r1I1LXhPwJCgf5q/0QQVsp6m9WesTdegBf+E1tY0H3PzVu44S9FRF4Aw
wqSGO+2zdIaqpmUEIiXKq8mj8wGpAKqcVe6QNRpzwk1+vR8rOJJAIZCJV7cy
1I67OUM+BleDkyEqJ/GX1sBFP3J5YENzrxhCTUtkwIOtCQ2j6ueBuKXoq9zx
l7sqsLRvHYSLt17/dClA5CQp1UPPMpuKUzwMJXTb0cv+XdPq4xozIul1vF7k
jEZtJG7znlAhyVMu0bXzAkaHysjkwSe64qP60N5NmjzyZysxw5q/YpZQ/qod
r47b9jqgNRgL2vPUEqgV3nHub1sYeXylYfrYUurmiENG80SB/LBnIimkDJuV
o4BG977DnwwpujvqFU5nulwY3BpHqO9pJmRNCjdvzSunhriyvaSJDj5qfbRE
Btnfr0wiBB9L9xrhB8hWfiO4YOOUlae/VcryqZNKZ1LTXVe5GXyJscHvoB0y
JBQS1hVyUJjb3IwquX4vBqN28r8dMuomuU2RvGEwrL3IqmwSBaXDAr5GOl7Z
x7Tfvg5gWzWgftmduBU/Ru+aeCLmUfJG/Hw3R5wXxbLMXQWxWJBzrY5khH9X
SOF0UT5XH8XSGQMPMYgDSU4upb8k1jiiMVJlK1VClJprhkSvghGKaC0x3IXM
xlJPIonO6Y/UP3+2G1jZbgjkJZKhYKRF60fvOlrgQVB/QT5+D6xeZCrYYYt3
5qcp6N2C26qMXMZdla0jHtUoj9C6nUZIQtA8SaVujTOioH+VniFjQCMTyjWg
HbLRI6SMGSTmNr1cTyci/i8VOO8bFAtX8oFJSF4OzS0BhEQEISVWhmhc8LSG
IW/GXcq0UVxa7QFlEpSPQvGTdA6L67BfSkK4lNy1rLvoF4S0Gbda4fqE1CiW
FW5jXcqfpwDhmZwXjxmqPR5P+VjdZdjMsYBjoB0gDfeUZwJIkMMGp4hCAhoe
L1Kzpb/EslEsNo50zbC3BfLZFLyctbxkDgW+D5NK2cA+d5lAwjLY9/RhemYF
dqtMAKyPZ9HiARstCV+i+GWbVN0vEHxXFNYc8zhdxjk0TZeFR2TjXRXOMvDC
+//GpmZVHP6r7p1P2egJFihYy4jRJShI5jbECpVqs6wpcAZugHlKaQ8TeI9l
dgY73WSQDfABLAZrc/3RZ96R6N7soNxmzOkS9Xr4xBDohB2smnIg0kAwBBPy
L97VLw7PZg9EHQP2Kj3PoUhuf1ls6CAx7YyPAizs2jZKv/V1bCvQ9fZFjpay
fuRvjd/wwr3N1SK51GV/Dsk50FZcpbIvcB8yHuA7RkIRHSDTgpL/FIUqFDoh
5QxDczTjAbZ24Gsf3FZIOCaZRZL/k5Z5W9nqI9Y9k6R2kCvHZ5y/scF3jeYL
rQsYGnOaQhfUBG1YXqg/NWHQfSLsVRO+YW06C8DL+0sWJFD+GY+4AiJkZhaj
CInBiZcfiP6euZ6SjDkCcj2uor0m3wY/xA8Hzu+vUe+NoUSVJNFtkAboEcpe
WVPP2Uf2r3OZ29SMu69jXn77phDP/zGYasHXKj/apG3Hgt2tl/R5U3A3h9YT
FE0m4FjRUD4DcXkbHJlL+diRYTOYcQfZ5BnOdKYAT1wK6FkUtBMr2P93hNZA
hcMmSmvxhO6dEQ1LqGYwAC08euBdsv2sgYdzYw6pmrpKj22mcDRJrXmFwD49
hSyohveHFqC4gN/ujXRRzEddtNtf0aQM/KRVVo0X/KeCnIaOPYgUuSxvRxUX
M7O58vw3BszPw8TtN0tnCQTWswH4J+cAx58dku/7uzwLCr8jLhJhHs9bbwyG
V10o1UPShZ2ixkiCeniDv9dJOcpzhz7x9jM7nNpTjjdGCWzdqKhWw5EqqrCE
iaDro8lB2WmzDAuyeyHIEuK/1rman5FWdAzGUpMJ/r05RacRiBpkR1BQbHTi
1Y6gY82TdRQj8Lb1qdRODTr/H0HJCkzugLFIdOPyGa2BXFKC0uF2cIdEMvmT
rrpLg2p5M4i1iAC3Aa1pfzeMfOiOgXxfmjxpcWRDrKhucIU2Y00Pw69X3+NM
dz44DYX1B2fZX3ll1/QuCI73fYHPGSdQdmfVP3xaHFzB4KYa4UxXZNmr1MwS
/bjKG5NJmo40KfCiKKopVH6PRYSLARHP5v9YD5lhShiXBZHEHLls4lMQ+nCd
NysfULQEkgG+ON2j7Ta2Gblj4CcozZozCnZvDjYb4CxW35YjwISrLDXnUno+
1COysh1EA/2Nz88SCCVlRuxPENTVQPvzAc47kqfG0LjRHznSctF4Y0aVeirD
vdvfAW4gLMx6oYSAVz1W8bs0aRM4OcjcRo+ufQfZeMx6kigUr9puk7KvVwd+
CeJMiTBJyJuf//MyROv9QW5hILlfoLYkQBSIFFI1L17OtgoDey0PzzCRGrRK
C+3ctQA8A8aGL2Qj/QdB8ZZAUFmEPrvQFU2V4cmS31zA75c7jVaF4kpQY0YW
WvA5I0atVhQNa6gM13zTkVqY50JcLxgM8jxEO533S/t3pFppM/mDr0UzRFYc
OhsZNtBxx7tXQkfNxm/UkDLf1PrweHYt4yQ7HtMLi9DcNNXRQs3liJlRBHei
5Bhd8juIYVmeEp3YDaiMDDa/jcjSK/XetMFHqw5N3prZLWy5d5N7YKO5u1vx
+1HaV4+qydD1hNGWoeThnbwVvK0ZFX2dYty8d9HE0Q6kHV4Mbmia4e+9vm80
Wlr7tdnjNzVgQNgzTUdSwDgxyTisspCAA9rutpVM2bSQVbQIr0vyefPTODgV
+FnKSAEq9t/bdmliA0+n/zxC4/NVc8L5TkATJkDwIFyYeXlOSABtxcmmLUJ1
/my6vgBYwAbmQgpGzsn1ZKrzGbfUhJZfFKucXP6XrzvNMY+FrJf5g3G/+oJs
OUQfDV5vRvvsC0oz//qne9N6eNfns109N+iLIDihBHAL2ziboV80j444UCya
JZKDKTWi2X1fMyjy+daPcLsz0rlVU5BE4KgEu+X4pw5kwvrK129lvvTcoh7g
WOmbvKDnQQrAAPj+rZ/urV/DHVExnybAMj5z5NiBe1+x3Mz3iicoa2SbZEKJ
VZWDyKTajB+4on62zcAbfJXuJ5PANAF5zKvKmzN+en7+JS9Jj5Ub7Ksco0Rk
UVraKTnOlCir261XucoVHKo797TpdMYoLuoJIXs2oPhcoWWyRx5wPfWX9daJ
4pWLmA8afk2AKn/29WzeSvcBVEAmGMbXzolTk6/yFyWoZxlz47FQCYWi9EFa
73B9mj6RKf7B9/xmM69ieTz4qolYA9AIRBGO3+7svwSxJJd9Mjw9WYw9OQsE
FXiGztfSbIthB1sTCLOke/eDhWVhdyoGQFYHQcYdPX9Yjd/oBJ5+1JT/T0Nk
WvKacNPvu7t9q2J2ABzGBLBe97wvVOGIth9BijPmWqVZUXX27P3RD5a5+3+N
m85BHRdeZINx3oGLgWds2g57wF+Te+4giom52/17nwVJbDIHaREkV63ZtVU7
kpAdn8mpcjRa3iLuLmBpbkWEc5Kca6DQ8KPtiI/vBFmyoqiKiuewrSV4uVFt
JlFOTTZLP0NikYo44wbHDzS5+epT551P9qvG2W/w4MniRHxqEs4+sDgzlf2K
L7XOvQuhw3iPoqKB9QmHqJJgBxPq2x+FPNhGXDmDdhxKsJbFE/dOjRvo4TYQ
RCxFwNtyhHWCHGUDkV9j0AMCNLLUxFq5bPPluNVxLbHjDjg6QSH7qNfZJPiK
d23OMSx0+zTxwtrsNh/gs8z6ZF5sTSBoWLkgXLx0C1jEm/fzhOTdzbCnjY28
jXcVSXD5/QSMkBKc6v84lXjCgB/x1rRfeF1CF+WAzrO/j64WIwfR3G9Cgpbo
AfI9SHy9PoM2kJNCClwBuk2PSSGWn4lPbz0sj94bZQQ7Uqig9ShthS+tp5Fq
mg0vm3LxFJwGv5LZuIs5ZqcBn/e63MQ+9JQ559z0BS8Brdr8G/2RVfQf7IDj
VuzulUD8cmpOPEyCaLYz8ehUM2U/x0/+nDjLQ8MYCN4PZflO55jat36nKORL
PkyAkle2Mq0O9zxKo6Ezft9HHszMCJZ+EFSxHfoaYoUmIK6Wx8VZ5trM8UT9
yAuo7kSlQKvxUoVQdWJxDCZEEznLw300yIo+yWUXFQ5FvyjFDKNekEtTeE/N
Br5A5PR7blhvBBi/moeelkMnwk5DZLj/xiD9bh6X9VHQK9lu2bFV+O2IjpUZ
qZxc3+2KkuAp3n5dvs1wYS8Cjkowi3s28D7iYe0mWoiw0vdPyu5pBwwqXjxJ
DWtREFaKK5vYy4BxnVWJ4pLizoac88dlCJ9zxr/d0FFRNi64TIRal8ldZ1z7
GiXTyg0xsb5WZtGqzGiOaYwhZGmWzaM3oAyZmaUnxF+ixRrBQRZ8mCYbdHsq
SlEOcbt7uHIcYRwt+5DW1IUtXJj8d4FNsJgL9LtyKnb6jCteIFdYNNxgkQ+U
Sf61zL/hBU3vg1KltkWxNhmAPVP4I4tjcdhCyzw03ewmlqGENdQbSts5soIY
7g3jilHbYgjHjnR141XpuQ7KsGCYXLdX6bnH7ULY+SK7DLDK0nS/rtTilI/x
k7DqZy0dAk20c7WUPnZYmOi64uCoItlW+OljKFKAj3vr/1iFWdhOLggB0d5y
KKciLc0QSyIrgPj0Q2HYBrDCqBq6IVnHmXT8bwOihWpQMppRxtGt7+bIFeuD
LwiyUfw+eOIArQV7B8amBMnspdGTZYJJkwfIg94wP6Xdgic51w0phA/5GMDp
Qi7J6/5kFBmbNCALnJTpLIjqMaRcHDUdup76E8i1pX5i3QKiF7Jszml3n76d
mKFl8AIq66pcJnMgbrWVwk+VX9P4e9JBXa6aH26T34qWPMMQnjF6gkdz62jh
IUnHNkOGJzCidFJa3ULpcZeRE+r+mnwkii2MbwVD71Rx9kst8oC+kQNe+26h
OSXyxHyF5HKhyJp8ne+WjbZ9yxN4mdj+/GLg7nHE+uo75am0yF3N7u7JfGEj
FXezA2Z1AEPAcI5IpY/0e/fYxGKHy8+M+QhHuXA+atg51Vd5BDfcTjT4Vo4s
Ap8H19wJ3N2CWAPUS74pQSQ0+Hs6oiKtj/17tNjONQdrmVJGmZP05A4MZVdn
9hmdrJApXAdL3Y+1Lex3ZD2CWadDKkgOm3R6GitvZKjJJLUlPGKoFMi3CM/s
PzuVv6q8sXTyXxM/1ynDYn7pocj7VecdvS8JSBWMpOMM/d2JPnq9+WpahGMY
5NR9MaIo0iyZIRIZQllYPLIy3rwQdwMTsa74Xd7z8K7IZ9DuRYHEanGvYZKz
UxB4UjMOCTX8eoHTITdFTntrArdMtVhMwz0hYxgFKXyGGhyUt+a2xse3ROTS
6sWSqDrsJxnqkR1/s5fC3SapAVI7MngqSJWfvHhabbEjsA3YqdOfrT7Hw0U6
xArmishmleBmrv4g1d8TKuzkl0iC7skuGFDWh2iZZiPTRo16kBLwUT7A7LLD
CcWOPJs2TBPzulhyDY8ijaM5NrAPMyVNungs42u3Z9/LQ1ty7KC9J8AW4+Vb
VpTJjzc3+pHwQLmjpWgVMEB34Vq56qgShq54UZ0tXfjtrwHhc0JGFzWS7fOf
r5gSOg1NaF4QLlyqM4AAKzlmaENwbz2QE9vF/VOTpf/o8bGEp5CQLDsAgJtF
YZXhmziGOgsNhm6VBXH1/ZpjH+npjc4WxTUjS3wLPgEb8NlwzDECN79luO3M
JAFuNoES3ZDW93sKCmyfbqrJlGrQWzxwXy4ui/0BvQAb49mphuYUl94byAI/
4uBXhy/C1ygyJQ5wp+I8rVaY+Lv86sXNn11Z1wTyowRQ/76nBmN4pEM1R26H
JKWX+GhXPgLv2FmoWjuTcok4NZsd0Jj8yGt7xsMROzCheCDBqRZUc/aT2MDK
6ontuRzA8TdWswD41lH9Xzj25HMHDpK+CBMmMEPdaKjkXGkoN3ruwYqgx1re
3VA+9R4VURWQymSJ5YNLEFR2hSWofLdMsl0j3B38XOQuMZV0Q9FTT70cHykz
DU7kP5XxSlVPmtybufPQAiNmSMxXypRVsOepc1qNmtQmrf2aWPn7odBxvt31
u13CEwjotH07i3Gn9EFtR+iA5bqovWWknuKVvgy0bm2OYpfRKUslkkMdU1AR
YfgwuiAc4Wh3VLSTc0aj4ahRrIcKHPZ+h0Obx7SXv6rMvZSDvuKrIyligujE
aIWjFjO1oNSuCSjOyMqByAmM7EtMqtAvzOVMtQaWP5AvRjv981tJ0whYNO3J
hrR8aiivq5+UFdOuwSRmdbX8SyEjWp2EM9wxz7nswm1gZCx7rP58Zg63DKGX
4UiVbvsNE5Ft0jkPEBLime0Fkn+Q4Q7zFJmfndP2SP5LT9WAQpBYIEcB6YR6
8oVwCYmNKgiBhG2ObgY/1mYQOrT3yVSUkJS6PUb1mN+92jcbZz6DulbuEUsI
wUXmhRs/Z5kC8OHfLEXAouaUV8aRirdv6KdJ2dghE0Lfj3DZdVBV3w92gGq3
9d6vS0LCzSPiNQIDvbOKjY/XsxTONau0cbdgH7tMjyhNaLWgqwCpWCyX4ae7
RgNef4kJ5lt/zQyCsv0TLA5KQ47QAF4wTDVe2TZ7coZ37NdiENQcL3E89CCZ
RAai7utcALaZNBuD5+UDrTCBACJrO3VQ+aTsGTLsZaps2pEcFi1IvgWYKAeR
a8a2eBmN4HoiRjL/TFINWvaVVFWDDF7y61lovl7Ihxdi7Oz+4D3T/IdZn2B5
VPsg1fcoqXHIGykFdTrUXt8yQuzdMGC5bCzZG+JxpNJ80poyHn0cWude7fX3
B3L3DIYJVZ0Bd7PBnBXF+YwMrmzeNkDv9NGSSNpc4ru9DtK8tk+Os+q4NgYB
+qyuhk1ilGovynxleYB+BFbRUHJpuEb2R3zd+TRuXwvi4k1dh6odP61zyPKf
MLwWrryMlndQsnQUmDMLkaLurd+CnMoeBd+lcqchv8Ds+1mz0qINxZBCcKuD
a26Ntc24rXUH6pFXJz6H5wKIcuE3aKuBJhfMCFxp0CiE+CmuKRWqiUT+h8fw
3oWjJAvqiVz5rRVtbF8c0aH5p3zKFHiDFaBCEVaFBEa6seJw99XmkSAtiit3
XGtCwhdoy0g+TLxdKQctzOcaxTs7j475ZETqrBmz2HndwMgeFw1Obh1k2Bkf
OIrA7IwLiami5Ex/ud2EG7QkHeIwMSuX/nFgoz2M081xDC8dOF7zypd526yh
+fP4mbILxes6T0AHwO+ouECiLjQOb4e/9UuWzhLLB6IpKyGwYuiTZO2KpNW6
e6UPaYPgIe9a8ngRdoUGY+pvbjNNiDFkKLFEhdNWhkIwvGgM97X7MOS03cdW
6z6JpLTTq112arKWSX8pVxB4hCV2u3dDQ5h+z3yz5VIU1gpwLoDDaipUSeOW
hQG5r2y4BOt1n59Cv7eXVixyct+NapAvOb4eHNBqOktCmDpEfk6bNQB4uYNq
7GqI+RPmFXrSyc37QG+/2Z0nJjY/cKJj9AVItiypAcwvCaTVLkYcTpQnWnQ8
um4cfxd8kodZjYig7ups17A+z0RHGwi2wGXAAXWskk94uhlEbvgxDY7IS5Q/
CdcQ6G+UVorjMWdc/fcW8iPUTjDuVBZlLDlPgqS/NONGlbGE8ZUn5fzfT+jR
YgaHrfnUUXB1hbbqDgO1PLdrfjtT9s6u0WcZu9io1QcZvvgOe/8+Zd7cGaF3
/g8m1XAbTVQnJdyg3lZRg6Qb3uBLCYxspbKDt7ySKzgIaoR07HLLl77d6Ywq
mZE0a9llmJLWQjLWwU92z3TILAUQpKAeg/jb7JbsNKSUbVAdwEFD9CGrqPSM
AryUZ8pwPEpSbg7GKIh4N8QeoF1OPGNfBn9EXuIQh5CCfZliWKK8/tV2SIsj
vze6l63zjec8BKj05ik2dZDxb7r4TXaMcI9PdRBi77BGChwO7t2AqLn6Mxhm
dM6jTtsCC1NWzyoTFYh+ogXNdZhmGCfEpq+w0j0BazESdVO/j5lN6q1+5U36
7+d6ecMEnxAGm4zNc9aa7xGfd3HHWCx6sQVXLFOjP1b4UH7ZoRs+Cvqmy5DU
xbtFkysRKSY6+hwEneUMMkjmhxiYdNkZ5IQ1LSD4P1kIlEkeFEV9BiyCKYGe
pTBZyB27ec2iRMGGKel9UCr0Q1s1Be5rYx71OyeF4vVjUpcveYRoJ6SqdGh0
a8HOQlqY2hrZ3F/VBzl8KTmOtaffAlSMYd5PBJTpJZ/yzN9eTyqgtOZy7JOG
kAQhMD0mxexfD8BBvOAGcRERV7q3V/BTXplGhYv/p9MejqUypBe93p4O5ceS
7P2ZaOzXzFiP7pDqTuWfK1P1hHwEsmv9HFkVFKWFYetk6pBESZLwur5DTY6C
MF3phmftk+89dpg6yiCZEkZ+w8vhKtfepoxzHYgK0LiBSwe8xYJrAAb2uCsZ
qwDzEUQh7RJ+vy95zjiKudMJvXIKUsI/941mRlYc74P+t/TVkf/z4wv3bchA
cb+dL9YX61mjBrcJL/uAAFmI95pZx16CKbXt2DoJKHEkKRDVJuj6YhrLOR+Y
GncDni/ouSL0QyQKUyMLFUqlYm3uqvB8Cf13NUez5R8qqadVetKps2sCW7uJ
vDIFw5fGeAhd6B2CHLulrzjpItLdD++cTMDbh7WOiCFOQIEm1a01XgjvpzPD
Ho6L3nkhmlcG655IHj52UrVALUq0tVahsl1XBQ27W+mQKJTpRG4djlij6yN+
DfnajsfWkSQ08BLHYh8w0PZ7+RHLP233xW73l1HWbow1EuFwTXBWM2TwzSeh
1ydNFRdrGDx/iktfEBCyqUU0ym8BBWopJDgpLrFmLWe+fF0EF94dyPXaLA63
D7ms/I97/SYZRDwC06Sk96p7FeDqwc1RmGe4YeAPb1EQi8/0j9qtGYQGDl1v
Dczns0Up8JNFZIGLqzt+c30NL98I9LM6Xw4tj3hLwn7Ep0MHUClQTgEz3+uk
VkmNyG/ZSY5SkKAoxULtLYnFSYawRP6SJTGnw86pEZnQpa4O0CrvLjIkBEy1
35RCwaKoebkKZK9FBg3sPv6/VZyL0pQkJQfgqeE9ZhhGRJrGcAZkWeuaxKR+
KdCau3Hx71dkE2h37S/l1IxFLo9EZYD0fixW01dH4IxW0/BwebI1YsUpTkvO
Y1EYMOYGRPVWblGNVbsH9i/oHATY5cJjG5sODwMqgK/0sbLDTWHur8NALnAK
C/dC5JJw2KY+HJk9wnuvzdAQ0BH6PVaMoufnNngf59+cMlhvXrHwfplVvwwB
d9qpaxSfF55N3R7d7egxgZmAOgP4i1957vgE+d+V0sTr6TblvMVuheBs7REa
El9i8jmQNdI/+mo+RRx1tUxo9UfIxjuzTvtXDA45XjF3Zu34WQwP5uZo/r0i
6WfRwiwSpe8xMiHsjAB5WZKEc5JJA907xtiLiCvWRpRjV7lbQMgskUlNcJ5D
Q7L635NNULrMdfmwQErrZEK8Dzj4l+RwC+BhCRhvk6lc29UHhJ/1vFuIIsCR
pGzcv0UGTIyfZetVN0pSO20WE2jFqiDuh0pxo3GXfnLTtLX5Kzhl86d9b/0x
guxXuecNnqBHi5BgVKVe8YHbat8XDia/73jb+sp4UmWyRfl7bMJ12HPm3/7L
r6ceWf2LU/5CqwEpdPWDlWUYMGwNCPKRvC/xJkZ8rKbc5+f7BJHMBw+0NjPZ
6Duk3eeFVp6VP+deBCugUaWZdQW2D6Dkwl4dyntX/nNIMlWz72hdH97ar9pf
ZWKm5zu8P/vEIUwOav7on/3V3fIWP0IjMG+qs6D//FT84qL2C0ZJdER2fWQp
O99nWrQVqrkCF44HQnHrUuDU7zFmr1ip30YgB9GstkeFrmjAZbm6zt0G/smy
mXpKUZ5vThp6HqdGcvWlk8cHHZuoPsiJIITTE+vyKPSLBjUb9IwnxpQvBqb6
9gJRWzSEImH4qVj1RbntrGt4Eb1Sud4KFSql4H69BvxfduTgOQFV4XlZlC0g
xTgWDT819s1/6chvwFLVxKHopfa0DDhJ+voDdUj2EXFs/CReDm9N/0wLGj/m
7Q49r6k9exksAS8LmygYZ08j6bhqiOa+SgYZSlr7TLMlcKGv7QxLDcgd59O2
IZg+6OYmGtFWPKubDXKPXGSTtd0yCZtan7VwL21Cc5ekd9R1uL6aluoRKKoY
rRC7t9OHF0TcMIXNSk5iKYkJtBBmKFcNSAJ9y162AmPuyD2bIxWu10LjtUfq
ahgyBc8qcGrdA9JiFHiQaQOXuW3hneHOobF+n4kQUqp760VQSTKeZOirgkVF
e20iHKmA6tWi5HzN4rPFYrEnGGrsd5n0BN4UbafAKPE5BByf48kI7nvAcz8H
vmvysMm1qry3nTneGRWvPcgYnG09wsSF+6WjO5nuKQxAwyl87w4MGDmoOaq/
3lNva9zCFVhWK5w44MlitV+z1SWhUjJfeMSDwI7mURg60BRt8X3Q24oerg0f
5fQQB6T/mVjme1akU0w3WYxq6uMMvTQnM3h7GsofAuzUHZrR9kwdqeK+OB4/
xag9qr2f+T4RqR0KclWSAbGnVGoW/1Pn9ZT8s4e2QP3x9bPTwl2mJmWd1Be4
+N4WYIk6az1epCSo8JDE9TwAo5FGX4jhgz8PNs5AAdIDFVzbMA8Y5yrGbWrv
47SvjwYShFAsBU6Pn5CtPYG9iCdt8cR/UbsCDD6qhz5EHDM9mdWeogaLkQSe
YhTIH3dy6GqUW/uFm9f/P2FulbMzafhPN6mwvfzDi6FFYtb3SGEYY8xmz13/
TXF1EkJPR8k4wiec6xPFQnTiQpuhxTohwmc6L0a0MXGflqUK3ighZQ/y5d2o
bUCDYnMuw7ILFEaad+amBkHt756DdVQg8XRDdWawRg2Z7MkQdE45lQJsEVKb
tYEJoS/5m52jjahvCKqxERaZDemIJRsxLXiTvG3xuo/9PauChwbCymocxRYB
s+EmbypU8IS5pwLEkPwCGnG3UkrDJ5uRnpBah524GwpOW9tKqSe+Yd8TUHlp
RZ57cZSaUAIjqpDBTp8VCg13carREgqW18LBZmbRQtHFsECp2WWi+Ir0wj1w
osl8c04BO/IdU7h8KCtIu+5I2GXmuBWOYmxoNH47uCQ67mSwQrMBkrUiEDw0
fucVj2Md7be7IBi0ASj+rSryL0SWwG4R4V9Y7f/dbKI/mmFs5V+DmOIMAaWA
rDDAJ7VZm4npQRTyGSq2d4zSHogN1zIXp79H0maDxAZsAk/9s8s81mvXxfWa
TJhhWDVcsOmdOmN3oASfqa+kTZuUlxCoIgBiyRXT3JIrsomzbtsqM/55iEjb
5wcXkUX//T3zZKB2wUJvDde97u0x7AUOaHLu5Tqi6pjWHEcKrhWKNp8Imy1q
m2t8ASjBz7pWDJXegVg62ghqVfweV50ZHUpIqXoiC/KqtcgE2SclsjyK5UOu
isxvJGjVGTRpxIJfveMOr+GJYnXYET/yY0zvZA845uOmxmLvuIspJO2fLsCV
XQXxeNqhMnYHiSUEKAqeITj97PzcAlOPFT4hVuCx8Sw9kjFlUEAtwYCUP7Gp
ioxbWLs/P1UnpzLx8WeAwoMVLUNTbDffqbvSfPRqIq1OD313MvF1v6U1KyRi
adcAYOSULp1BecZtz8CKrGETHGRd9WzvtmO3r+zzt4jox6qOJv5gcd/1WxzJ
7owN5BtHnIzsHi3nalLFwoNrbhNnmV8yCDOEKn4OXhZjHIs9l300CwEIhbrj
Iwi2i3YqYM4S3w+d6pccqqaxREJp7XMPnhmt65MxUJiDvjDumfiZScrcx5nr
LRlsHrRqIxxhe/GwZgVzOaXGkypJnc7I7obkMTc1Hy4/pSpZYApe4qVPuaz8
YlnLXR/JGYO8+WXX4wCTpyxsH5GI5WzDIaX2xNqUEUtMuUNsJisHdYMsdg7c
vfGiIqcGUTuVKk5vTEIMoCxH9WmJA4HnOBWBy4J0d1zhKi49Kbaco2OW/gQa
32im2lb6KeWYOEwq/8liFxx+QWatnussoW4KbSmNKH3ObZHCN0lMNGZ4lrEY
DoOi6517rBZIY+q0hTlSt5Ka9cR2MOw4eEnCAStGeAat2dzpgjSfXJuNsRTl
XgM2/KvBytq/SjPsJxffJ0fEcf9/2PAmTOkbRrdAl3h4hLASZyBcP4jlUvAr
/O6ikU1gmBD7yDNO272aNlwoFGU704byFKRuqOVQmZhzX3wk9oZsiea2UOV2
2U2n4eyln/G+K6HomBo6lRbSchpUWhaf/hScjFaeyodyw3ZzPN+xMCsF68C1
EAcWJwN/tlTOpmHgDD1b2qlmhK6qaZnaOSnS45F0yNZ1h3C3/FdGvw7L6bOO
kfArBo1wmU/gSaaazjL+/u2lfjqwJDUJLBl8cBNh/H/mPPdm6P34ObpjJhF6
NR19aNcoajr3fJ6s5OzmKmncLim2G/mG6YTahd9/P8q2MvLRwyPWMNwyXLro
4g6qeUKds9sDPcDJtBnSWpxiZw4x7c1fpDDsptVFCco0zUk6wCo4bW07TpH1
HbG21He0pvv1KFeKPda87hvnjcrTeKqT7jK4UgcK1CU8kF3Lfk1ElDGPH4dP
7Y6zIhIlGzl7y7kTVjsAIzyzS7lh1h/gRQHqV76u7xrh4dNUqrJNNRWtvX8G
nCe7vLJD5dELtCZq28Moop8gfKaGrrmD7td4tL+Ju988aCrk1h9px2mhLJSt
ZKuSfrrBnzkhjdtwy38+1DSD+FlvpjQKTF8OE76UTi06gh6fLiGvl+3YTCfE
yTEBUzz+H7sNdeTxZTDFpGf9ssXxpvl7baF9AGneOlW5p/dROOqmNR7v3Zqu
OcAQLGJNOGjH8J0ffQXcnKDDGs5IY3sfYnZg0VVlm4Hesu7QLxFYbv6g/idE
0JIcRlLi/LUyDLwu8vY5KPjyaWamrUyRJhX2EAwiFlDpwEjOwzZg/95b74Sz
xf6tKeY2W78EPeU83Tmn7ZmX4V5JvEYFZXd5ySkmXC07kPjzLzCAu74z44od
i+BZuuFAOhwxDGhJXCEqgyNRXMgQrsYVXpzKksXNxrOz2h34h12A9vztRe8V
sK+3LBXf9N8uRyuY21G7wkOkGmA+LLxCEThK+Ybgv39fQk30pG870oaAxvVq
KuWhkvQrtsVdz5tUznM+h9ZfhDvq0KfoC2Ln8fqscOWK+vMG9gGOVEXq9HEd
2ffJ4+p4+dzuDqmgOZ5nWFPL3PKUgccA0zLqwZURKoD4I1arQEo74e+kyWsq
Bwy6hnnebLpADcmDu9Fo/Xevekv9O/p2ubkODxmFzm7216UjvU41gYQkWpIP
+ca/xW8vTwYDaQ8sfySZ0bQK1kFaReGx4RqpEcW00fLrPrVpyh8Iry278uea
VtUSKTjYgwdSrRbQqyl9grg0eHMo7tDI6tkKxOPo6MHLtSgoMXeW75l8kzbD
AGHOw012HV7E7v/wfLKcWvW5YxRvv+0in784NwVSSJSOaoAfek67gp+YhX6u
nnrVkZvw8gHbh5TGjKvGULnSF5w59UZ6uU3I+splewrVU7KII5Ehv2+O+Sx0
NnJzZbDO8RG1NPQTXZgmV9rjIIUcQhG8hT/sBSVGjBBSeyx3bYhIaPJke2z+
pv8duRf8e1DIH2p/vyJJVLAhTKkx6lL2jP+7W2pqaWPG/UgQJZZeQh0Y+6Uy
PGSOIhs4VeVq/Z6MxMAH+P4Tis90Bv7HDDnngmg8z+NmpReL5xPPJzmYBoqc
wbgIlLGw/w6tdKCZLgrgZEQIcwgfNGZ45RTuh+mZmAy+zK7Q6/CzZBNgX0p+
KDG+3fQaIwdCBjJnd46QQRqcUnRzd1G9Wg2iMENRPu9214ajgk6iZ+Y6GW1F
fvgCP8B5EtzFEp5ytUCmbozCHwVOaNPLGhoVPKOivSluyxINwl7Wo48sAZFC
G9hRcuYXMDZMOjzOuB+InupFmxMApjEjywGnCpotF0Uce5K1UNjzge2Iqfis
SoYdaM7IKaorZ2ac/ikyT8X6TR+iulCt9+y/8khar2vO0GsjNekr7tAYEOLS
WfuDVCqTbLTPntdnfOQYDaPN51F2Nem9DWcP/xZMy44mnc2jKDgYV9EyKB88
zRo6qiTH9iIP0/BdUKVWtDwrY4TNGOQ9xrsYdK7VdlWbzYQPC2z8dbUhlfDR
W9wUNULIGugH3PNCywFZuM1TUboRUVs6H214GoDt+VCe4KW7Wvo4NNW0/83/
90h6BZ9KEWZSA3Rkn/QU9tRXAXG48F8fz4AOS304km5qcm66XAPEogIvz7qC
gyyC468WZewPnAyLbnZ8ItnABYaKU41EWw0KPOdpj7e/wCbnnSB0Y1eoXr2K
u7mMyFw7gbwYW2dw7VQYnP7X3+Mq1xHyiB/1p00d7sJLTlZWVNkt7f2bSd6Z
JAw2oxjzDPaKanK5PzjFDzNEX9KP+OUhruHaik2XhZ0wxiZ7ks9um9VPyc/f
rxvlCDmkLpJORyzbyk4HHCeo95UqJ+bPYKZ08DhJIJBaRcWlEjOEqsvgW0Wr
xng73bMTRilcZkB2QNOaaQqP8ihdQpDfMMMyc5AopRT599F8gB8rJJAGD4Uv
jDSUCJbR/FbQn58paCS6+8aKKTuIBTCfYFkEoCt1GXG5TG5lZ/vfDCorNaOQ
3+3kQi6bq1XuEIJx6sjF6Qrm8F4hZJO/gJY6jCuJfvoo2ctuADSk4jl4amMU
bUVkyl9fECKkfzezcm7E/WZYXgyP8c4FNung90SohV28WHPM75yCXU+tBw0j
kv9eef6KXeiTAY4wt2kl+ZFH/+AWuvwAbVZwVkPHNWW+wSxCO9aprfyBnQJm
+iIoTTF/QH4VtYDBdHatrjaDtz/FBsJW0KniAEm2DQNFDWFbw124F+dBUmHX
4PnENNqz3/5LKYXRc9r6amkhO3LStS0WuhYOc8bIhiXjR7BL+EfM4iQ98PGE
xAUpWwuwtNvzfV+cqxjRzcOcwKye0GDmbSQMzMO3qrcm7cF7P17scm7IqXOk
8Dl6mx5UV6AlcnS1lvFMMoz8GY4UXOaqVTdj/SlAYUR7XyLQGIpIzv4+2yhu
5igcmMHP7pMTKkNVhigbAOSwATpiTMyzguDECeq8K8x9DCeWrHyapbqFQTxX
9EthtI5trSUnRw5GNv2f2XZ0bXi+oKEEGXmQ7CY1LshecGVbPNzHGPED9L9B
StBL2d528uP3xnzIiG5TLFfioC0loddIcMQQeAWcql7Wlc7arlb4qUCdPG64
weul+X2JV68UiE8+YBgRllpIHGgbKvC0E+KaDtP5g6VYcWqIEzmZ6qF7JPfL
6hzpq0i0YphoF3LzJSeSueUlRTa3ZUmoS4hIWxn5fwZc8LgEg6Vz1krgRWnJ
6Yjk1JViICsiNxDwstzlEqBzwtTlDn74y0bS6EzBBBq43r6rZ6AAgXW+WZWU
NpQhPvBpYIemU9uV/sjymXK6oGAxN/2DEoeXvwpYPjrn+Z7HvMl7EG+dWFr+
s9Jua3o+Tbu8tF9YKRo2gmDexphGR3AEMX4X8neI1wgqYAwMZOAB6dud8MVb
6UkYVKINMnBok4QPsIiPK4uHS3+dmIBaU7Dy6YkGvjz+BLv65Pfa+vRZyIW2
iIvxiAv7zV4IF53lnUZ6Oe4sMm9BgfRN9fKaH8xmxnlzemkWYXkii7b2jxxp
1qgAouiHLiqHus10+S9TtRpp0xvfYRvjN5hfgjd5d+BxQGAip6OOVkos2SZ5
IdKV48Wz9tTwuKJtdgKaYU8BYyFATWt3ZmpGmzSy9PwUiPePvUOJy4p0AKa2
YM6zsak3j6F+ZSYPRN22Lnl4zGIgLzB1PY6HF9FtBsysWDvnAU4COO4Ll2UT
ej3Jyy0xukMBYe5fIC9YfHI3O90bvsbSZhq1stS8ULVo9dLkp2wxqeGCq31F
0znsm0ye7GyulG3Irt0HEkrRMfH18qEy4W5ioEAMzYrKbpudnyao1zcgN1vF
8Np8r7zDgEnVR3Om49KR6lJ5TSaUEi27NqMqvoIiw6Coz0rZXtCM8RNRpKAZ
v/QAgzv7yvEafyTMzoLHgJgm2QnreY2teBOFWwYqhevsDjjYJq4NqVEehguE
RTvAyMt1i4GTVbOIAQhRLCFuGin+Dx9AS9hsA9rhiu2Q6XhKyIh56cS0liip
ErNbI4jgrOjmtS7s9roiJ1XxOPEPtxcWX6fJws/e8mDd7wHpSdNjPqrWjck8
psM2aBxW+RgI9d9Pa+UkqPrjgrbmC+3pRGbC2Nq3ULF2FZTwq9ayuGrfJiM5
NyDU5tF0dPrraZDHDxPVFaSBkZfrZwSQIoz+46vKsbzcUATgvoT1wlGJn2nJ
daZ1X9+62WYat3E8NzhwY/lxzhktF4qFR24tsu77MylyKwRUtH30E3XSH6Mk
uC+FNlbmPRhU/RfMy3MELY+LahMmNBcMg7Y4H2yK7nRXhM0KQ8ptE+k7ojpA
qWbnM2be9O54RUU9N92ykaawnAxlqyrNwxCpxmgJlu//3+LwPfZvhkoml+Bc
dIUDvmhmUjwwIkeGepGi1nEANsb2EVwPqU4R10CV3VzZVW72gLHMHUIliSrY
lj3tyIL0b8UWVU0a3q87mrXdJQS470c3T6Eevpib0YuROJTshQF+aCtp9fch
koilLDlBqkLWAu9NJ2EJtXTx9qLXAzRsBCUyTUXBroE1XhTTvRXKWy9NmHLa
JLxNhFZrEoskVHYHgcEjSh1IdwJmdx8AKTu0aPtoBHMXFV+9KBOYKCRO3cFN
mKVK5kY/7UHF804O4bOiAM5TlNWf3zFWGGONtWkRNwgwIrDj2cZ19L5Nqb4p
LUChs9y5SRxp/++zCEL87Tv45ii5nYFAtQSU/z126IGdNO2z9ZiW2+jIx6hw
IQnMmayOgc5HiGCdKSFbxCVUxHgOpRE1D7n/EfwYQtRt0UEDvGPTBkq/wLNK
26XqRQdJ2MLlJ5ueGWuK3nS7Whld/HT3CWgcFGznEK2s2BkV6qaxJdY9QJ8J
LIvmnAC4nYD4jE63SyrBBIbAq+zMofpODCmDdVMMKz8w/1AYVCTKMu7ZmeYr
jXsCHUfRCCCTADCGhjyGa0zf2SFXq1rziwscxWc7DXKkfEiHaFfPCzQFQ/fQ
x+L6z/oWUTb1SEsoLoBd0subDA7Vk+k59s11IAJzQmnfjkfabNXUxEnh0MeA
LC6Mt+rBEInfVGMsNmvgf7HCEndT/KF4NxB/v1JYZhQSjLmEb9z4gDzv+PYK
Qyf+MhbxvICbskgef9QICTifQjHhgxU7kOlWw6v6VpifjR5m45eOsfY0sULY
SvKxFmAYx6gPcwa/t4G1aVsKvWvAvPSzoxDvqp+XYVPcJx9VOkbsAHmHmK5N
HKPvq7QzFHhIlOX30DixeZ68EjODFPPOT63TnW9N4I45rYrIpCjMZbCPKta7
4StC7go8sYs/9uOBgZn4wx9MexjLsVjWELUULqYYjq2hH2dqheeQkEvVSN3M
BDScK4ZFQZr+FTzaJFsvGbXwoy/jkKo5PHO7mGw+k0RwiYEeSdHyB24rN7zf
CfOfGa7SdkD6cy9x34qeDvXFgAGDFievCfUMB1SzNfvJ+m5A7sQnN3ZzDPWy
A4vsL0YGxaSCFUYDqRaGfHcUnUoY82xW1jpwbBx6pkoEqqf6UHvWSDZEqbmm
nAnRjxCAKYTT31HVy0+jhHVV9Htj0wimlLMJg+1OgQZ8vJC01fKT/51ZWIDp
CUWwBT0gV+YpS/dEK1Z9yLnHkLcO3iedJGH58AJoDM1KgRP0aL/X4MDfymy2
aWAga3SKuwdbYMJeOkp+m2jqCK/W7YF4lOZsw6k2qwyY5B6EphqNdHP2GPCX
FsRk7844rBJlsYYt0R0kurV3CDX0uz1j7ZMURvDSeEt0YIacIgmCnzoFhDE9
ouHJ1ByHjS1k1ljOiZOWB7M6aloSh7yKrC71UByjJyDDszbjpaZBE5Sb7Gdh
YMQPUcJLhbFeRcVYI0tyYvzLyJSLkQtWbwi/76hElI/ICrAZSvrkFsGQUj++
s+4Qy8vcqYRAiBketCI9A/6guZZbHO8Ghsm14bZ8pUyVsU72t/fd/uqys4Ns
ZTJ5s2ORc9Ki1ugq5G9UIRV47aCALoRee9lghPG4Po0XexVCcnQhRPluzHtc
3uLdvNCJieTpzCvoeMjRbFl8E0GD7KSOZNdTlFP7cTt8Btr+rHuHAnXwxaK4
ZiFP2g0V5ZI1wFygXMLxoWonslkUzUImbsFntLhPrdtjboF8vNV4fwR2Mxjf
Mwdb94QBE029jps91Bl2OsDW7oNJCsD+4u/4KSpf69bJQeYA7M5929m6VNYg
jmftIrBL2Emh6GshqzYEp6MBC5R5iiCQtRTB62i9auP4qXZldurZCYFt8i8S
9zIkVmsk4LMpCT++UqkcE4zPOIQPGeMBuZjbZ/f72IZORiYbaoduFTvp7nIw
I8P3g1dIj6RzLFXxRa7b2+qDJz4CRllgal7ZeBN7ikxQNe/6sWiEib1GQ9l7
DK7SaAG2ZB1HHD1Ku2u++e1tDHPZIdt4VFXXEolUaSs0PV6FXCLnAAQ13/3a
SOFEiBKSruArXGizoORy6muOPblQUfMdQjr1SmY2O7w6gdS67slhaY/CkwbG
Wvw6xjKCbqU5fwfZIVGBX4bYmpoiLmtJlA4hwwIPJ6eYjm0qLxYD6FxgqDyR
LkB7krH22+m+Q+uhvWTKVq57zwzmDOBHyfaTspj3fNftUXl9W6WuhVKKjqNq
uc9y746Re8KSuex/9o+pXjWqgmM18wNsSF93T++vWbMyCsjVjSCaONsbzDm5
o3i3xPXpHxE9I1tj30+jZ4zVVkFnvNSBprwPWUPC6o16J/pwDtuJSoTWjMtk
Bjk791yxK3AA16RW/yYeBS3lhc3rghkCyoaN81mizO3lc6gbTCZZChpxkYYr
T0ilBoORuDaqnc6UF39FKFUnpSgjSJSy2WnEGv8C6ZlmOEAkFE9wn3Xu2aVL
cufcyR+RjbNNqCDP5HEYfh/5O1sjpSL4SR3yiy8sMPEwmnVsqFtqXujyZvgP
M30n2bFuyq0OvsdWknBsIohFSmuDyMLg8nE6p8FvpZV+mVImBPuXKF5csqkY
mbe+WHt304cpoU2CEB6GLHDc+cA8nQEOkeBsiKYtGESRfKoo9ndvuYgzqIoo
2IkVVZ0B/0laSBQGaekvVCDxgJyTnC3Oo7j6oplGqmhcw1+hwoqd2qEzjEcR
n8TyoC4PE7bFPMZ1WwcCjNUaXs4LpJgiS7oT7c7RxUSV2BRJ5befYO4Mc+Ff
1sRo8VStBF9hdxQ0BBgOlLI1L8cdNdG/Qka13ssKBGirpdD1TIqGPZz4r1Eb
bKRjYAZoweSfJj1v9mg0fU1/hS2PU1JVA+1JZZvG5U6K7QW7RRrw82KdHgzs
5m8zy99LH5UF6ChKQwd/y5N+o+w61Jxi561eEzE54Sn/8J2euJ4UmrJrw+7k
szyAx809n/pXCmDuFzmRj+Mfi6QXKqPEb/79wxrJzvr8jHQ0I397E7tY2jkT
LzKPj6fdm4OLqiIcoVWmm0ywjPOtuQJqAntc+5VrvGcCp7J15g+tVgkFgV4I
Hyz6wM1t0UsWv2vDl3rRssUmi4nguBy7D/N+ttg+7LMvLSG6mahlCA+hcnGg
c9E/bBjBXg/ziI+xLD8Yl9r0no4pbthzHxa16Sp+sOzcPswSAfY3fIGkXOX0
OxF7Gbn/4r8PQA8RGO9zHaOV4SSsL3/2IB3dGioWWHLaCi27EYCD/OSJKPOi
DShPiWhOV3JXCTWTO/+RqbNttRVUJKCOifx+2y66X7/rO1YgmW04WRiiu2EF
uQSUbzvYUYs/Dx0p9OzRN7UX9Aid9wbHQ2jyVAzW3U0s1dUEhWNL84H46hMy
5OIbSyIMEdCmfHyS7yYnxeMigOB9+m4WdS53crg61H92gI9X3YWY911KCVVV
t6Yr8kPnRVN+GMjefuCGKoM24jG/ZDKe1RKgC9QPBDx2zJRW4UJvANaSO281
py7d8hToo/JxNSYq0fb/Cl2JWkjtsR2a302yT647McPwPXnslC+SKt7+BIFV
MZGHLzWEU7UTlED2zf/PO7QK1krQcTSt4v3EBDOsYvAfgq9nTKBXJrxyR4++
sv8NF6iXwS88o4SCwv9YCOtsPcKGKWTjz+V20g2GGIOful1Q68j9PlbVtF9B
WIwbAxpUN1GprXE3wTQhqMCRg7RcEFoh5/hkmQyQGK9q1OuUYMexWtECO0Kq
TObVeXexZ2AR/xfG3BWnHg5qES1AN1lcplHGAP5lESVhsg/Ikm01MBzIVi1o
LLaplwMewP3NozrWxcXFBucs308Cjo3edoP/R+FkqJ4pRi1sLNBtQdgb+g9T
awyY6Fa3t662xS4SLWDH4Sq2JWEwOOFckA5jf0IqB70DU1030ZQlmFjtH5Sx
8KZ8a4PHzOraQGrJx5sifsgiHdMje3XEQnmVURsUeTtrjJngOW8uvQurhf3p
7X+hVJ7k74AFUjJP8qxnQl0WLimDH5B2mRw1/wnqRoydvzum9sq33xXII/Mq
RW5HTE2j1owG9ivhnzxd5LffnikFbNoIys2xajjw9LUMCba1RUicXMATBRVq
t3WOoZwXbkb+Hhut98FgZR0OCQqg5BpyiPeWvuzNFRCWRm8Mqum9asryA1GX
CEj4ov+eo/+0TYKEwmUOL/xfn+RU0Ax27wYPigzkHjJN751z5kAw5GLVVgT2
qX7AscKixO4iLlHcRudFAgRtzyfiOIjw7qYVWgEBwKuTKc3sKdL5ede2mUb6
YzAilPjpDSftHjJdfug1fC/iFFXunjQCagFYNqo7PpwRGBdMXC5liYk05wUe
mIdsmBAHZblE2hFJNlyqNKLOHRt6BL4RkIQP3qBOl23/0mBLDyTvA05wOXtw
UwiQxKpTj8VdBZWpJnyT8nb9vmTxNkRgKObDlhTTCB/ABPSu1DPcMQ5duNd+
ZK9gCDOQTU5FFCuUX51o9jt0tocH4RvKOTcA6ARs6rgoIXplwwwjIhejju0j
Yl3eoOBA3RVWO38JYdNWP1YRnxxJB+C9rZ36KxL3VLhebtBXMqh7k/Ey35vO
ar6PIi66fd36Ycws2XXJd9NJEl5Rv9eFeV87tXZtQc8LLBm9TNcj3ZzCmJSs
bTak6b3VG4yqZcg8dtFdJbmABLvc1Ecc7APhrrpIUDuOT+CAtjyV5pCjVw1G
xnaWPkhNC+cEzvFTpf912jbDAXGUKIWQCIpuR4Lp6Akfi3/WmVTyyCQtU9MO
0o80o9ywZFs2S7DOKe2Sb2W22eutnBQM9o9CokMn/u2gOQ9pibj8oe0ilLGq
VJWKpJhDZnHpfL3tQT8QKsSFJqM2kq4MzdpZToDRLuxRQSD+RoaaX7Ii26Qm
mOAieMm2YYMT48HZDdT31JVbSgUl0MuBN3qd8Ikmd4VNW0yWfBpK89KtRKq8
X1uwqRir43z5VNudBaSQBK0ZahLZi3t1E7NXSh+1p2VSCul9xYEu1dC+ZzJQ
Li1dI6jXkDLfZUvBEJu1WEdeAvSaTmH/YBd7zFD2c9POtYB9oDmCcltg8z6n
zQETVG2/iDlSuB2HCYBvZUWEJz9YfcfTSiw6cR6Ru2CRairIiScpn9IWu6My
qM/FnRUwrvHR1ZGNH6tPJAbGqtPBAgv5m8vVRo4Ud9m2nwMcCfB511mNZk5p
QqS/utUhw8v8yuwnM23TD/1XDAjbCk8eAdgniVxo1GkJj83yuRcAsfpEXJ4K
Z2deWxJlBVHmaBJZdVnT1uz6VWcH3juzIOSSrTeXLL/2xCURl9D0K9xIyTSp
hW90hbwMERi+2BzH7EyVeoKhG5LJS0DOPorXlQfcmc/dj+VO1Dr0/AFDAxfq
kws/LisGe6Zln/cNJHhU2I3vK9sKtJ8f6HqBlv6Bud801idttr64NujBXifU
fiMkEzJvnvL3CxByd7s3ZsMPaC8SIp0xD1lMQ1XexkMcHjdE1mbgglQHDbDN
ZZzey4zJUBnCXU5mmOv8/Jk1vnid5ZyufxZbHuoiYBjm1btzgrVxrGNS1dT1
TXdP+GgjR6L5C042wQrwDW0yaT8uT2cAOgpPoqO5RuOZ7FCdsuSkQ24YCT9Z
EDvEMwe9QLrCSKpzy2g7n596KV47F2KCgG30aoENB0n6/4QlvqtQzSWp1uFX
WnG+tYiSDEoin6yd4ZVvNfNjDOK1KceHmNfDBqML4BoA9Wj5MCTMwG+rYomb
MlgKm3gl55S2iNhKUhLIsOPbh4LM5cZSCPkJHYSWgohzjeYiKxZe3yAhbMgs
dyWJLsomeQhWQaEv/WejX6khIbrWh44E9b3en0mRSvOowgqtCRDCYfY+dAQl
HskbAJ6p+EtmE7x8dDrS/Mw3OvNk5PoOLDt5ME5FP8rdqUAFRzql9nW3tqcW
V5wx0H6d+9G/PTy/u5xWgWZNnsoUIE7Ebi1ftABQtbHfX5lCt80YItGtWKS6
jqkj6CTgRHrSZSqTiEmsXQE/dfTcBXjYcFLFnsX6O66EQC/yNp1r8w6Tgk+d
aItZbHjOknOoiG9iXgOYzfBDqoGAF5VYn0sBEJfQoBvv8lJS9JibUyTpas0x
MWPtB1OnOq+JcsQ0L/kCvMauHL4zqFRatEl2dnNYC0wm3PixOAvigHFV6a7R
TRK9MAdvtk9FxLcNj3fHufe5CwkEgTCDI35YSSHFdowSJQbDWoXcCj5ePs4I
nww6rGPidDkYitRUC0G9hUiNZY+N0ZZoanFBqpmJ4MxkipP0mThvby/IGjUT
FOJzrwUxm6mxPGfXGUgBc/baXYLXau7XzbIJS7SMC1yNXmn3dV577R5jCa8x
E5Xptte1XxPhpBwWou/bt5ONWO7gzRxlm0CORjD0/Bp6EPImfeBn3EagFE01
gnPK8GLhCX+39e/4Jd54GRLBdB6XIPJ2ERlSVHY3ackrxdyBpYrn5qIqqBw7
CkSdEpXGh5Wk9jK2YznFjSi1BRMPFYFYSh9s+6tchU2/+a7rP4Aigvphl2gR
XCW8JFuw38XiG2BZhGQ0oYPucdrY3QTLPy9POSLCZQSsEKcbaKgY1Ahe1l/C
uXkrRamNsKpKQrAdDdp943tpoXWTNLAdqRTyeBopXIRWZ6mzvvMFUpC8BlNJ
KS2ajXU4jAjAhPkm73UaE2pB84rF1QicSIZq1TthpyZjHE9ENUP3rmwtMzFN
tMnmC5jwKutHtkTeNKWa4Li5U/n9HRQkJGVlxnjNkdoPqi3JJZwLDPiTJIxE
gSxGPrHZhpuqZlQvhlBkvFXwLCxnDpabp8ucxe0Zx8OcX0zXeYOwAUlblaDi
8aY6a2Rz05gBGsQ+mBbMGRm0fw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1KuWGBbRkN76o/Ia+vqAsS1fMv6zQx7mSbPbid34oxpBqyl/Y9Ht7NU9rKxiNIqC3ewoBT1TlIomt4sTqtzSQlk6YqPgmoesYI8hJJu8KK1wK9ZYCR7VWy7V04ozwB4uA1zy8Cxv85xncvldF57iystRIuUgD0z9WPjS6h93P7FLlhzQ5fg91v7oGKuR5GWwkiCsYJdb+neYRjSUINuiNr/0wWajSeSX2MrkmwfzTqQO6Nk4r5J3htdmFmX6W+93nRudA7N5dIwOd+hRPD+CmoRqjd8CH2MKVLP8sykFwd7marSzEcb8y2gSQfA7ctMBNS64h7j+Eq/AAC0v2D0kDGny1zSw1hwidrTFATcrtmiIU3gp/9vEsMvCoc3f6sPIbyN0IZj86XUeu0X/gHpa+3345UNy43GLvStNWjcaPCzkhy1eGywk3PNO1MZLYfeJDL4lPh3YW4pWlFV7MnUHzeeGSon6M97swN44nKCQqsLLmecIJON1lgIAhCRFsmxQwibXC3updnhU/379nBYuVnDYSbw6OQkb5BOyx1H2KSqJPwE8/aoMPODOA2o4D5DgzaG1+HS7b80s11lDgmWRXQtnQxSftJ71Bm5WPgdbe32JKgHSRH7SU+VcZy2s+b5l9ekFq7ey/hR867k/85xGH7U9abigRrWGXuXFgiYvJnrgSctd4pOdW93VD1R2cV3vEhbAYk03A8YJ0iNNwE+YdkPaGaa0bUpOWNHOuX5cS39JArNoAUTjpc8sEbRtxEJD26SSIpyTa/pGR+NMWCPVZ5n"
`endif