// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iquwU6XhStpARghj8UWxX1bSFSASjWpzQhHpUuSFkiJ1vZYEd/IAYWf4rKRQ
KIWUApC+BQ1IpnY/v7BH6b/5MOb2JvkPE1n9bUC09E/bj3Tmf1xmRCulWnvu
2SaruClddeuXmrtuv4uqS3KblPQlqjgTrA8HMLscnRoDdpcV75CwGrJGuZSn
NHGiJCmcR3Ui3b9BuVdHLD9uuCQAyyFMlqjKe4vg71HLL4MF0P8aRQ92FegX
34JiVhDG6blHXolEuPQ6gHhmdZ+MaoLVlfEbS5tw8unCVCiFQnOdkTFCzy7s
C/PLifisBZLQvlkZJcU63EBgPAuSeljD1mPmEgUyAw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qqd/rceit87w44P7fD8ops6Si0tNMosQFWMzRpqB35UsfiT4NFLnR0yzvSIg
6n7swQDBHOhfW3IBFJj/P/8vVL3qEpllP4UxVe9xcsE4njKHIjthMnGM8MU3
q44BHPsBegtwu+v3kKMMosaZqfJROwJns+viJ9BJnlOmkfhUuMh7EtCRJrRY
NB6xDL5PKqfdkIFUB3dk2pphT4fkZBEOaWn5JbM1GZtCQIFK59kZMpQyalRd
g5ztzBitB0UvXWPjWoXfV7EUK16R7mqOd7PxhhpJrNDKf7YKuMGcS9OmpsoX
pSQMhBnliiNh5SUDT2oRNJ+5MzVr/o9kHKPUIxlRHQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tJDEMqsTgbzg7Vv4lq4tUWoRHwwxigKZZOqQauOajITqnYPpsNLJdekjNm5G
MudVQ4g7bCc/4na5dVeO2C0QFRpCzrw/h1k3SCl5T3rAmRVOOEOAaGLQCYyD
UJsBrD1Mo8LKWJxrC9lxETFfcVAWuMiGDt8g6e2qapFhQOnJ16hMy8WRnlcX
w8euWsO5Y/nNPBGBN/mbLPznOd79S35o3mgkwYsyENkhNeCIrMWyjyt7WVwG
JmPfFFHwGJa1u+uRFLkA4Cu+IouFbIz7Sg3r5TQq53ylbRf0Kl///2f4vAwI
VyDy3xd/LVdOq8hej2EUhFqisCIaZ6ADdXOEpfePQw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Lu9MpOG6XydARczeak+CIGwZwwXdGaKsCV6WGz2XHVO9laiTA626NJHgXoyp
bKd2iG7Z242x00M8MmTUsR1kur816qtIpTn+kiFpGgObZsTcC76+GizQhUca
A/rYqaXiTgM5Rws7gfllzBe+xdboI6mPcdj83cEENx72/6AnTGmDvwMfAH37
bOshqbQiALkKbyk61lOXRyHJ0LoGTF1j0x2POwCGnOBQYli6zYwweKAZJKYW
tgmrWEGvdR5qwOP4d/Rzep6gq6qhleJRN4p6v/8WDl0L89oEU1kdrRBCv8Mp
IAAYMfG1XIO/Ir25lI3TeDV0gIPJ7kizt7O+0i6qEQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JpmKKYSIMp/4/cbT76Na3kQCeiGrB+7dLJZuucEpaX61aObluYcWRL1zLaRO
I0/ZYotnGBO2JvhVFM3wbVPVu52bL/KR+Im1EysofxGD4wnEHEE5jugg5KKZ
nbnKIufBYic+OwAMUoI2FUGs8cXZ8OjRuXbl0hL9z4h+cOrJxBc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
rTuZ2UPcmIFNgzFTq77bzTH1cVkmHv9N/kdpXaTqydsHO+UbAVl6clZxQ+Bh
jI/r9lcYoRXgXU9kPzrZXqhgMWexuRhEXm6/8bRhAGsJLYcz8rZ8FCTe/wAv
fS+iKSENKBLAF9fCTxza1HNzsC9XYGElkQwux3XptLCoiN+IpIrSchR8wPqQ
Q3D8qjZ5q382DRShKBaEscI8TLpJu86xrHE+sHebk+K5J7NzBrUQppjLJqbz
ARPdjONyAOcHcIJ3JathPbDwAOkesFCAf7MFynzwz4YtZOWMKo4I1L26xlFI
Twl/0ptsEltqvSZWAFuUEY3shaAa8/aA0of6QY7XG8CD2FlhaVzNs/TPugCK
3Y2gIn292T+1TiE6jx+k1Rmr9+mA3mMPgYSL1DxJo753Tx6J7G3Viq7Ny15E
pL3gP35FfLvRmr4y3XshimFreMICPV+KHYBMik/K5NGKZTIYiuPcw6Vyif3d
lmzqGoYFD1frkaVnSnzDA3FDFIAR76Gk


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fqTIrKYh7GkvDN8hSoHvkeLmh4QRuXZZko0oNpNefpw4vZsU9rNAg3GzDZQ1
APAJXFBhtNeITOFu5FjPY32A709szUDx3tOCoToKybUdmvqQCSdy6xQFlNKm
GRwIXPM6CkzSKvJfX29Yx3fhLPpjy1v7tdOVzO3eplcAqez2zjg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YpivqwM7gyoLZVmsESwjl8qnYlG2I4DHJ5JrpXEvh6RmDqDtiGmx0iiA3gHa
V71co93wiZhkM9BJ84V9vtL9qB23gWN34ostVfewsm5ZlUkS9AJxCa5gGgVK
0hoiCVklkhvmYYUDFZ8ZmQ+LqPOlgKOFPYbqJ/qAsmEgVIe5Zqo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 91632)
`pragma protect data_block
lnowiY5KyGV63HoV9UKgz3b72rYTvExSvcGGp4sVZ+n9Rk1fE8WpR+nqSVi0
tUUh+7758fv1x3jULv78XrRJgYT4wt4eQCXEjHq3nxZLxGjjklhex3ATA2m4
aM6k/3+wUDjfYe4jrw2+TvAuBjwzSurMrn50TJzs3VVCU7YK/Z6Ozf/f11TL
/NLbLfWr/ncHdd6qm7jqds7bD2phk3ALsB6qlUSDXplWaYDbAEkPgxhbE4Fe
xqqc1xOfPaM70Y9i3W8pArKLpNQ5LVMU4F6FHb5jsyFRRqxPz1DMXqX81d11
EYXQTIKh/2YnlOUw2rDmN7T7rQZjO0OyqgLGQ2EME3JMb/5vQMkzVeS2oopQ
APkhUT6LdNE+wRlhISl2o3m5mSykfvuqFJiMw5+N30ynGWd1nrDK1DVUwAOP
mx8Kn3m5GC/5Miqt0sFaotCjuFbn96H0EwYVBVGmOAog3RL6EsyrQ0KrYcID
mCfZD0kyviNoLwjmhxW9ibrafqOZ8dyj/Zzreznm2GrUEuP2uI5JgDmsKeDI
8M9a7HmiGu2wGdwOWHrAnDAmWW8wRM7KEG/LL4zTLF50K5ycI+dqHmO2RCKb
tn07TNdixxazu2jnqu4wsvMMmu18BGAsPbUtRJ9FVel9MtfzI4MdLcvSIwBJ
C8YOMw7lHmCczLRPQKtE2RYdIOQRqpI3YGQ8BWNdzh4Zql7iWgwNnKsPFxjn
IAYoKCSvd/a7DV2M5TYYZV58VaBpb7/+c2rpaZN3+SlGszUpoW29NYQnHWZq
z3CFejhze5/z6DGfPKgZhnxV7SKjqzdvYVRt9N7W7LpAQ6YoP06Qjd4kj3Dq
jmPpAJSFM9z1roYXnrvHIprkX/0jxguRAM5K7tltyf2zrIMeaNCgQcIO1NCb
79X+mZrtquRjNV+yZwE9CYuy1MYaRDWzv75KSnVHlE2QbiYW+EuN/zkjxa6f
C9sCX4v1XlOzyYTU7QDdJZAOJKTOJnRDXfX38BNorIhJnvLbyVdEIEBKUe9M
8oPPvvKcYO+hTGkQm83iG0DnNu4K4iSK/6cRtKGg902iX37UjU9ZcvVwPKlW
J6mSxRM5MtSWllcH1nuJJcCDrO8EMGHuDEXhHB6nCzutgsQk09a4lsJfKIfq
jHduOW6Swp1uoPdtJNUEt1AGOoCAtbd8TbimdCHAs+3CFZykZrbnp233d8he
hlsfzwHjs5CGAEXUqaodY7YlpoqOPwNlt50KCva8Usd84WBQdSFdxyxA9tmw
V9BW8lAfzO9VLN1Qha/o4JommB3TvPkBiXKkdVJMswAiQC1G/aq4V5+lWheI
d0DMgxzGqyL65ya7afMMadRMU+UPMQvha49dU2k7CPzS0MYnLASShZD0RBTM
nyW678ekDtSoutPYB4tlLkJPEN50BWUQjKw5GvZcO6vhD84SoXJPl9s4NVr0
LvPcgAsF98IxfZBN+inWQsIoPKmkLL+yCmKzN2vesei8YJciIayAuCgzdhLw
h6+2BPgXlp84y6/6ihS+5cRcIaLpXm9NCK0+ZZXrnzGjlYxIxaFiVk3bT3ox
83yDvgsRYWIYQW2XKFsE3Oeb4ghX4pfh5aYVbUdGAXbP+I5Hcgp/xXxFTDBx
L9Bh8dfnktgacJ8Uclosm125gQFKcOvqTb5LR8jJeAS2MXXT5slIvpqhvFaj
Yv8XJRdC/4GZPHFh13m5c29pfF5oibTwBKJrf/WsuLAayEYQKb6FPRnSHVZp
mZQA1dtrPfCJB7pDYn/19yfpEemLueQQ6wi4Uz8rS01guP4ds5SKRT93iSEv
5JrEW6A94GVC8eUNNvskfzT5Nuu9oGvHDGJcHDNVQC/B/FSltR7lV5Xbnok2
2F1U+JcwC8U2+ZNglS5P8OL8i9ARSq38FaaeI6HJg1bTPZ13WtyuIyoAkYz2
vdng3KkLUUuxCgw2NjwHmO/g959yF+Rro+oYeSuOjqgFaLibtMdgE0Pi2akQ
EIoHyxxtCScDwdWqOFRdFVPHiqgYZ+c+55ZHsMcfrh32vP5T04vWqqlyOggg
3WMqfpT2r86vcoHBinkGptE4Q85hoZoKFqBUQI8kZs8qIOK0RoHUWRzwipc1
rFIviY1jrNqsh5XlXuaBO7e+w67LV8msFgz6kFz048BwGAOKEe5e5FpONKS/
f4h06ohuIbc7BQ3LNDyepzY46aRuWybvb9tyKExAWnhAzGMiBKqb9/I7BVHd
z1IgQ4wV/kqbeLHN9WuHPJF+xMsIK/8OMaDGkkK6Y6XkOtoXBQPUS1FJBoqB
Pid/MWV4SPVW8x/BrJ/9kWxs3kM+Vsb5zziWXvs7ZQxiVLVP9NwdKLBJ/Xcx
ORzWEzy6jcTairaG/OoX+uFtbVTAxZUzgz+NwGqzlzGerLQvH1RqbaDHyMa0
+pZeJDLimgk/z4TAwow3Efg8NWSOKUxOkv0jzCB5Ib8ABYHgwIoZSLtgXY6j
DD/FJmEmk4QSKAGF10ykhrMk137vS3M9gNiXfTuJw0auVeCraPK6xaFCfT/h
aLXOVFRWTCKrvmVOpKRlNuGQx7peRdJFWHWqUzAQgBMflDFX5ngNzX6YaR2L
tQ1BIXGjDbBGUHJXxSeYvYDZKoS1tKwRPcMA50rjFEX1xy91BzRvxV+MdCJA
sQ2RupAj9CyX0AEsljQkDx8SSifC+VT0cIefGcvMuG1o2YEbpLfUigA/R0Up
2kNSbmdr6lLNw5OwmJlojsWwp6e7YedjILmoiN4otZL3uML6QBLHQyKUZrQS
YK17U7oDIhDce9MowMnXTa0yBmfufGTVvjEbrpiPStZAvC50rOQZtgwI7X92
ROfwOPuFUn8naI37JF1e8BAcW7l2JBaef0liotQVifsSyavsjOtFlzmPfffP
TSswWigomsVQPtC8V+UgR0MzrZz+DUe2Gf96k+IM2eC8lUEXXwE+exzvYuJi
LBIRziJG0Uh99GPSNmg9iKbtsgtS33fgKwdrIFeJI4o3tJo/dR12eieEQsUu
pHSSVQorwcYBO57XhsnUymDKIVx4qR1hTFLP2RXoP8Znoa5RPj3YBc1sQBzu
oP7fs7Qgpc6zzVy07LGk/kE0joWwk6QEj2NnOr3QQmO1oXjbOjqpfe0Ygpx9
C0U80Bq1YmjAWX9nxg5NNIjeBKkr0aHpYoAhT0E8MLwXvpNMoDJd6UoM19g9
atdva0nxr1Y9gAwa3pYvJZ9nqHXcFOjZO67co+97O5nTgX3Lc25bo2Gh43sS
L8EgJI7ZmAAuPNVO3UQRclYrktSjqkLzaupWs5vONjC5faNSdstYwC6qUon8
Rnp20XeTaN7ZlO6Q8O/6rqGyydIoYXWTuVWqF9baqcHOEGGzZkeGzlHd+xl7
W34f9oEce7Yrwt/6pTttc1LZd+s9JGH11keyNkS/OJCoLqfqxeKB/TTZbzBL
9ABqRkPW+VHMDBXTjcNzn0C84+RB1YOuGvSMA+Au1wW8+29GytN8RWSyNso4
0ZNAnKRY9seRG7BpAbMwlY6b9eJkziSibTrdqROJy5YSSCw9NJNRa5jXJFI7
EAfa6OLCpJrfbaOiAB6SRmCT4MLWuXRU/OBAPsf8uAQzlBTjrE140eZO4UpK
mYkUHRdFyYU4pdB6ObiMFaA///gyDYb2Dr4KBJJEUHwqilq6uCTsLOE5PGol
+Q9vQ7IeY2LVJbphypAxD3fih6t2pX2ugvc5/FeLANqvjWk0vu2aYmWiDIUP
xzTbb6JSYNtM3EUySEKEJxRzF7cdHmuM4Gw454b5djLvsCfKNHGpoJlg54MR
fjTCbkgyyROmO7+IgvdaR7YZqjFFtFamXJlTsQk1fIWy75gEFt8mUpsbZJhx
nX0Mp3thuBz6qHSfnqZYDqMaIvarpvl/JqTx5HTw/mG2tEmtcdiwqs/FD1ke
vW74kRqIwgCoU5SKVk7BQqOepl4PaIpsA56hzsnxDxetGlml8Do+l8wrz/ob
t8FAic0c1Qrr27yR3SQsCjme89NVbK/JGnUmuOyfWqzBba2OM0Y95EdLTmuz
dZ0Cmwf7QfU4PDZAWM7o/IIhEQgKq878stNZlJEBKBIj70W4LALDTmo49Ryz
rOAEEokEwU8mQJEfHk8T/CH4WdrRZLTLbH1ikNbJdkxDc4dAQ+yiSxYA7LCp
3+ni71gY62Pcu4hMhnbjGVGng3U9jPeRGnbWFszQTcFSPDqLD5ItMhc6p4mJ
F8CYTNxvX2hnNRqmn/zGfnLIHQWRt+Fhk0vX0Q6mDZj8ij+md0eNniq9u7AJ
myM8M+Ijf9zG/jCtjmbEsllgSqOH93FzCpiOdY5+q9hf5omL7+hYOzcsDyF3
fh4pyFZFoaXFfJNj5geR/LyfIJU9YxaFkwdpZQS+1Vf7uaHejFMAXLo6M8E9
9GVzKsw2RJmgCWRUm3gz49B3y2Gp+KqNbZCgukwTVDvaQBrdZiuN0BUzDD0u
CJBI7VJpuIUgYUv4Yu24t9y3kRyaBhPtWPiwsPiYAs+S5ekYQXoxIIHzkOxw
FIAAhO0vkobxnUePepyEwSSFC4F3FVDyf7AIvtnKlWf3XZs/yvMc1I9bfFyW
qAh6vGQkXHdxaJVoANv4hTadH7oWkE8ZAE/FRsoBB8OLwnaMy9VfpnRQR9+s
keqo4dMfCHqJ3wB8d8N87BxA3/YU1Ty14oGKfbWnwsqgv7uvcWDIBXkU5fY3
rZp99uzQhVEAz7au/gzKNIBq4brXJ7R67IQWzvGN4r9KYvw1zWZvlq8yHdv3
oZiBvm1HOJ2XW8e7ElUtL8gVxI+CGLcoWd1YnZhAXf3ycrtRtZvfXswlv6aV
hGUB6oYg6Z9trOLp6Ytb1nygtVax04EyH1oKV4mxbnf7JPr0mwaNAz9K6z62
QPSkB8VcN6QUXPwpLIqfHoqTsP2meMLFWgxFqAFF4M7r8wu9+S+rxeGehHRZ
/NrwObU9SD0InR8L5RZxp7MmerHscNemhW8CcP32BgaaLem4xzbyZh+QrJfD
OXjLbnZaKFqCoR5PyOqY6kje9U8BjuLhCuSGSRICf85gdtOlE1IroKhV21nZ
lVaGOUMRxw492cSyKlQh7p0dY/nxc34XGT2+jBOkHzIG/syTzC7LyLZgW5r0
jg2qwgM++KlBmZPf/4XF3b+iPgROPqr3eH/xQc2QmsLd+8RoipNCWLqh9wtj
doBUYhUvr1jfMo82M/MWwUpb6FAQ16ioeihUJA0EPvjQHr/QgbVKYX9FIrOB
fT0YTGyMofB2IOtXnUGZ1GUCnKNCSHqpHqD4ilkIESWf8K0IstvFneRFyuPm
v5Ti5ua315/qz4RGNHMBc5hvU4LnuNfqmRd697HHcUE4eZLbMEuBRVp14QMH
3t9xW5NdPYG7ju27PhFhWAExJQy6Xwe6OKrRZm2QZykNNRY1FImfr1H2j3m6
8c2hcHCPB2kNwfrdqIunsLZI35aEL8vXdqTmOLWpuaF40+wsnjS1NKt3xBBO
mez1qB9R6/6vDFYiiNc+BwwzN+JAeF5F0eIJT4/ZL8PzxP7jPNU9VW8IRVNA
IGlGQZmNeHBbtLClPiFc3QrcQAfCdzo8d9YCVcEsUGwVF/eQvcPSKGol2kTV
luij78pj+vqeNvsYdQTaCLIS+uQws5x49HgkF8UKgt8aAJwK8St3/dlQmA6Y
G0Cqv5HFYyGuucFbEtVzuBzlPtC9Z6ZqHAFtMr6pg7x72HjuMMK0VvftMmQD
EU+adMSgpZr6E7iGfGp4NIQmSZoADIjFqswirA0EZZ9s9oNpUwfCEdn6e1ua
KPnAXcOdD1OylLJhaPE9zAeCpxoDszgeuBnQ9RV+Lf0WpJ3GKFRwHJHZTej2
Wmt9YiMvGlDd0PsM12/VvW0+eLD+vaKR/7I3n3x/31+NuRnHWX3pQqbpWman
cpxOW4mipGhsffMMiBRuG0vDfOv3yWWTni+bh8HcXdHU1Vu85lXXhTBRs+Xr
iCmeTt1P0dd9+mKwRvBu/CLZda+EASBAZ2UIZa7x1qX3vJjlFUW+I7BKB7R/
RUex+i2G8EqifvP+kxyqIer7tBKG+98ieifzQorMVSa7qBkY+Pv+ZK88fh2p
+ztut5W6Cljk4gQWMHg8+SQ07MHeN/k0zadPFraaH+cJZxrpV7a1MNDJ5b1Q
TKJoYuDdEWN38QHBcSva+e4e1F4xcighfglhNJTiN2i9ggYz6H0QxdWn48lS
P6MdIuXu6VYxyE80gyEgiuQ9SX4r8ckeL3GJ2SkcsiN+YMs3z38qtbnc0NMt
jt1QHgqVXLkjVxln6Q9pJk+Beinuj5S/5H32zUFxz46xZlDceF5IGhMHtz7f
n2Jbh+qzonB0dy+Oo6xL18Fu4GEhPRh2WDvUREZCv1GE/YIyODybtNM+9Rri
TA/3Th+Wde2tuVT8rboqYLGcILtJl0KaeFz0T1yrRrFlwJv0ZuQCWF+ThEKo
G6HXLZbcHj8bX/1O/i6EiwN0L/qwSs1zb3ww5DevmcAjGMzOIQM3hnyCWrlA
fvDLgswAFmZqD0JrIvTQl69inoVBBI+3m/0Pou/VZitHg79fQKZAkAnbUY59
Mjw5y0sd7s8yF3M1M3o0VX3KdgzfAcYKBHm6IUHS4b0/SMqqoP6pUHZLtp+T
RhpNSNegNncA0cRHXs3Um6gFf7+1VmV4hkI6cqrL8FfKs5Xu/FCGHSPs+35P
CGI7K04ZxUFQY/PQ2a2qpg5o9nzdXTg6jTEfaXA9xCxHhGWkP5O4/OfwczvU
Azl54YY1gJBBxudZBij72rw1YTnxLK6ONZF35BrAc7gxqh1o+G2n+EeAlg5z
Ix++LdWU0WBgx9tBOWuAmhUnn34zDtU7YSqIKwH6L5Ymwq5m6o1rmmt8jua8
igyYFW1rxrTem3PmmrxjYHSfe7S7M1xiQ9IAMadSeZVeLtSCPmYIGXzWGz3C
iRbrhzdf4mY6+CbSzcxfimmdlV4dnk6uIC8oYtMAkCpyYCvXPT0U5salG9ov
GWBeDnvjNtOlo1EoxbhUWz2GC+30zU9wshrNfou3Yf8B8BcmyRKKGTB37r6D
+/Q8b8lbA4t8wNkG7hjGCaER6Vt0r8838dcvezA5rQfTEEm8ikaFvrZzno54
RZmveQ8ER5ef2VoCMefP3wdxP7bR6tElzszCHOVnYc01Y/pAxQxO2O7sC3Zm
kYTie4DzPgbRWW4GjPb3AbCfcquP7C34S9FEw99YlptrktnMB7zEvsvA2fba
kmTCmlwT3O3MiUEQq/w/sMrJNG9U2t+Ln5FOv5KsTzX9vAbHP6aVwrtdzKwk
OfZqO85wnxVleIO33OhpMSAxe4u3bagRB+J3ZdZQMXZfBBoTliEHS1YJroGJ
FRqBsiIoAOy/qjIFDt9wRRuXGjzoRal5ctF8R9eedvGj8Suxf5DLbyYbHtIT
fb0nWaCA3/G3ppubGf4ioPM4jwxk0DNjpfAz0ul7Ha+e/Ea+v1hSOElbGStp
qULCer5vX2yW52/zz9kHb6sZHSdlP0BjLZuv1aIVCG41O6pmrVRFfmheUfDT
qZUSQx28M+sYb5b+ACxRlinTsWCdx/GAqNmNeZEsejzpqQAjCJgc+POlEXGB
7ypYeEe7RIq8GT5KyfoAAG07LTvcEpiqD44TVGfP60ZSXmF7UtXvEQPQJMOW
hrnAtrxUH3oTGpe5/rgZa0RWYwRlKnhwbmbipsrd0/Rxq6dcAIoplktD+syi
T95RXVyWZl99WUvdFmUjz6UC8+5fmxfazrJN37oW61MMoTOvK9xSMV0GUf4L
pgAtqz6mp8WX36BaJITbgisFWcLih1p0ohcPpeOzUxoKum8DNPxo1oplrhTF
rfNGsTokM1nqyyNnHspoubu6GGvpot9FwP7dZXiXHjsx/lpFZqc40npalXV1
8YQxFqJYOBZcsmNk4Cq6QJnc6yKiPz6T2Z0tWPmva9p/JiPZ87VWg01p5iJK
kCskBhCfXJNTFkWCeBSE9GxzjQQMdSrsN5eGFHEe7jUNl1fO3CoHIHI5AoPw
L98S7ERRJKyAswNUO5/4J5QcgzeMUGU/3WmOGJEuiXbYkAuNbCDd56cG2Z6s
Ccd/7Nal3HcMPKymLvzV281iAIxsCalSWZBJ2S2tPLcdDMfbtYO7gm67YgWn
21wmEAMQjZ9oVJTeUPixggoiicr4XGjZ4E5AtEtFfVKcJhvGS0Ihorbufogt
M/Exj+75VsSYorLwnRA/7H1nfR1wqyhWSKJu5kSnrbVvRrgwV8NXLzU6vwGq
rEwoM3yxTY9zmn7ltiM2L/XJZJdUIpLvmBcF6JZbHVZNfCyPJOudOpz5taLd
W9uzgwluDxHS0NcAWuwpjKq8xOSrIZGKAmtfIAV6PMEh2cicG/PG5DJih1t/
4j0KU9nf2SeaQqET9pyLIUve3yMd1c8NLp+ZTMHaftI6/wekLUdqaoBMbw1c
BqrKavg2WDg1nOLjS8Sdz7TLL/vyvMQImmcd3QU0XQ7plfqYa6jIH4Z8angg
NUmMuL9cjkgELTpyWTo7M9lv3FeMcvpYWJMN3dZ7l73CSxNbQLOpP9eZACMX
1TaPhOguQBtTJyAd40RP2xMw8uwD8XE0kolvLPutbYfEIZC70aH5R56UjhPu
gUmwSh5ozeNimzaSAfC8eYiKRbesoSHiNJeOE+0wh+GepCMF82mKLxf6Wpl+
IGxAQ9jhleA/PqqRgYpNrWUZsFOx2cj56HHqunZ2nfSJuWPx9IZO3cnpxL4o
XfkKpKunw1GdOx0LXGZhuGXlhkXpKqTQN4FhycOwMaerj6gEPgk/mUwAP7R/
23EwGyOnI2NE8Ql6P6ByH5sB0hkotW8RE8RAxQD3gXzIFZVhfSEE7qdhW/BP
ekgyN7WbE1O8MhvcVojsx3j4iPdw7U6xwj0EkXl5yruefVueKsww6u0qw/RD
9hYRY48kLcIgTi60PN6WPlOvXr/mfVLIGYb4Fvs9w9r3TB1/m2W8c9NXSpYQ
jhEm2L0Q+kxiHYynfpnVQJZm1VAEdqffVvjEBPqNg5u+4eXECg4Gk7e9NC/l
hqkTWZKxuDf4mfYXYj/oXt1LKdQmoCQuidvhiFPo+AKH4A66RmE3lcYzFzjM
7pP7MkmHA3iVMRBomA9D9D3LK+22JFLPAF4sxXRoRAKRsGLpbkpnoFScqojN
u6gUmpArd+NvcaeNd7uE5LDx0rOOlSqBdam6bvE4H5MIEVMN3taNECpvRTgn
L+944vSSwV/44boMApACI+wFS6WfoxopZEJKH20q8OE28vVpqzxeR1fS/Hdb
wAvDnHZnQh77YS7F0PrWi+Nd01YBqea8VE3Fr/9sJgAUqGz6KOi0OlZvzrl7
lMYOKeB5jMzgfTVIKK5/zHKjZ0l/J8GmO86iJ3sOWV36lDsCkkQx7dhbrzuL
3UPIy+5DI7gDgmZwgsyDn71P6vPjS+ad0DVM+3fyGXlrKWuA4K4k1/LZe3WG
z0ocOGY0/7be6iGum2OygCdVbX6IdLbxhvfO8wFlg30d7tG5njKJNGveuVe6
SkDHK8CBYKLTBw8Ase4OBn3kYkTOUTtXYxxfZ0SEwAGZa3FrhlOw+jdn4L/K
7HT5CB2yyDGgTiQuOLTHGRAHjsLrjYpArwcmAojDQzJWpwa4lwNcTM6XuOaS
4N8xvWufqHp+IbwhHdF/y5JOzN6hvYi86i0SCamXHDoBYNJgyDvC4u2fdxth
0v0a4xl07rwgBOuJZIqfQjqGx0bEmHAbm90SAGIh0Vw4UJa4e47KlmckaOge
4LAWezUmVQDNE0ol778LyIP1PTTqItVTXuOTn25W3nl54ZqbB2S9RWWskVKU
As1L/CM8lMHXIuZr0neP+YsKtTaY7YIz6M5fh0jNLdgutWAXpUEHhghCTnEB
wO7wAI5OEDvjdHV9PvdqyRQXAmPJskyan31olaKfZPB967LzBWQfLdzl3RPS
mSdh5h8GePJ9W5Or3Xh8QrZCr56KXe23VCjRV1xdsmifgdf46biXKG2Cd6Fq
A2iPK/KF5LCCeMycMUUxYhPa7erkw84zl/vySItMa4+3s5f+fJ10BsMrmwvc
Wu0EOrpu4WIqb6qKSq2cUxhbUHnoTKU2lpIoHbtjJAhthWIvKp0P6ZLaBQz3
08gSRLvKAnPWlk1IEA9vRyphHBP3wHFkaU4/kxwukESlFMAefXld9i4n9E5S
yq0sjIzuy0TPnHUyLrGy6IctPu1+edfE0Qmb1Vqq3BMzkQi0waGMHk2lOBMD
+wn4jGPGu9UayTppCEDw5/AOg3ZiYqSQShKWjJPBsYvxqX5xseQKENjhRUAH
IW2OuIcETAjmSzVLlBGpaicVfDd/Vhe77krXlLRw9746xrVEy/T4m5o+HDw2
+4TSZwyigiyqOgcUW5L45EB/E76Gr7HtRFTJMM1QSq9Gta7xinFpVrBvx0BJ
2YcRtZml6yH0tNeTREhzDsomnYN/ce2N1IECNpbKwbl/afufbFYxbOtWOb4i
vl5stzetXD40vhIRjI/jp6ysHZJjs1jr0bLcVcjZzarwjwTadF+PeZ0oC6Ji
X1nvd39LqHXLvvH/dquXJd38g7VjYt8/gnuThI1+laXbtsfebn1s4Ufawb+n
FXDsbxpbeTM90nA46yQcJZM3yVEsr29cDSZh47HzrfBDovP9ryKX20Bxi6Sc
Z5NukHxtxTpoLKu50doEhk30EVYxsP/pLyD2zNq7ufss2kib+vamVdUhzX7Z
acCD3bqJ3msXOhF9QR8h1q2vCyMYtHm1/hAGZwbxYV8fX2wLmogJjOPIM0rx
dQ/EPvhGLSJXq+2eDlCufKZEaEunE3RR13t1CDEsYZOxgHCdAND7Rt6oGtpA
lWicyR5eS0fYJKbVIsTNyzAeh7/vNKBO4DQjBjFSNVNztfQmFhemWnkuQgrP
XJJArqHx1hjRKtmUhyrdF6UeGZEG9ZWD+fJxiAajXvMJzDJHaSvfGWre7/zG
beiVbIO6HgYQsJDU8rJEQqOKRbbt6R+yI92+3qCMZC0Rnvc+gamY6zj9MHCM
DrG/crUjrXLxrxPwF9YrDkTubmPNeXBq7ypXfS93xQ4o7yX25qwpHgQAdDGp
pMgPt3qiT2Gi5khwT9mB9xV2i0RKFbFmv8Pfr5KUE8MzThRT/0DyKO10fpn9
+rsz1K5n+l3q9fGeMrd2TsPK21oNq6ahwKy8rXSVa21tONubCvpRBwwLqcqD
46YmU608J6lTVtrwz17zrdTr6+QXSpm6WBjwUkGvQiPjNmGhQN1PUTbdog1Z
TLtRobmV1tAOEYEqtXKbKL0TTuyQ74VdNtj0N/UZQcAh66cZzhFGJEi6EL+A
dxDSAh4LjaH7fRD0OjzlR2uDYjAcd90ioF+lWKyrQcgwdIAZGICDO+AEl4kh
dWOnqpX2nS9WQVuYTUo9izUdQIfkctSxgFDddxr5/BYpiuT2byeFxNjnds3K
7K9twrASVyKtfW1u1WlSZW2lN/bn9uygW2IpTMghFtxuj+W1Hyaj3ttz567a
TMdwthR0FrtpZqRiVHxSMyG1m0Zsgpxv30UTpKt+nx6xwICJBlAPvP42wGaL
UMuSRMyUuMU2w8NuNgYHSi4S8vn4aSyI6hX9NWU1Pj4qY3HXANx5UWdD73Ra
AW5MLayOWIAyLVxn6lRMdlEfdVnrMqSc+aXw3wE86b0SLN8QRxeoLdfB3lSL
Rkv6F8jhbejs1MkhbyC94pVdUFjRbcWO0rOFxLE4IK5i1+FyBkfDB6/GII2E
gikcRgVTAipr2VoaJV8L58vuuU0j7eAXtPkGUzyxZ4/dbXt6v2PmJ0CvCNhX
DKDDXEK4sIgWQNGFFNXHGif0KazqPCsIYupKvAVAG+JYhD00Eo6ct79OicHC
PNS2ohBcrhTB3J4Sfpyde+W7EuUr2xpMowb7dpKPYqIfaWVYX/o7t7x3JWwE
246cfoPlzR/ATNObiKDOv2EbZ0cmw1GmyQNvLVlUjCFq2x45T+Aufcq7u7YO
0M37opLJR7wt8wli7PVpgdkwkLnazlDP3raElPx8kyskZnueVDAi2H4FwDh3
aCkutVfSEVQp2CeKrwyacsye+coEcLwG4FOpFb1dFbISgLsO7N1ROxGMyCVV
rOewIYRen3NUDkYQIQ10SBHCc6tC6qE8GeqNLjYBim9saePaW1oOKn72Nkad
pOAUztxXMrq63UkLNsI5zmRcX1Z/dbHUxGNVMNlYRLhXZFdQPTBuezBhCzm/
AMfxPNqHxds0K1cycF1QlAneF3cuaix314K13ctthGy8Jia5T2NKsMkBFOEW
8Lh5aqRpYs/e5uqytyrHPsSKt0kI1rohcTJ6KfmjwC/z4J0q60itqxWu+cHQ
6Zk37cAlTcODHgYgb+TJ8Li8+C/dt/WaD4TVvvJwxthS2MnX28LOPNYpqPr0
RIy6NPkdmbVICS38YAsET9pHZEtE7I57y17cf0Gku5UdcdKUEPY1i+zTnpFI
DNalHxIUFCLD6tZKIT+Jln/QNPqt7nBPvhXZiiKKob1GS2Mh1a1CEAZCfU4H
9bXTthowtgMB1dXJhE7f1JfQileBLdkaYvnUMZbm6vyFzmLFi4vAXUQeCArc
VOga2K7U+Izg5GqCGqrS+aTuPdxKJIOvdgtaBU1xXYgjaZnxGNI2N5Fjd5cI
3tHg0LCcmQ2QLfC2yIp6x42Fzl7GF7qtZRFFzZkn3LWdasAX40AIKAPe2/Le
XL2vsU9IYDBNVEZS6y4IgOPk+WAY3jgfnDYJ7uW7uMDuToE9BbFvz+bCa7mN
7cKKacKPuJrPKSPRtxlbH9z2xsv4XUceKzCQ0A7PCLE7E1Q6dG3RI9XLBdrT
+KGSPAGXOWsTdye/a/+7Ip+d+FhHBmUNjqqTH1FSWgbQ0qKk1GXJYnBYlDhK
FHalKV7jqKZxRJ4CKxURAcTx7LXj/c+Vzdvtcj7wFHG8JMUCCS6ABKEgEJQv
wBZr1ChPtsPziWXzYCLdDUmjKfbjbZtjP3BD2VGa90fZXqqub6KLHbvGWZrE
+ScqY+2sD4iYC752hVCqyb/LPnJMacNIEZyIYIFt2m2pXaGCxZZgjOT4Y7sm
33RLl0htTxBYXqMMsplzttnif+rtQv6aerXRk4TaRG9/ETXxrKuflw7UOpCV
Vjo4kOXKNH2Bsq82K6KrmuQ7EcHju6o5Qj09bK4O36IKo9j0iK68lnn5lLre
Jdvqxb1X6X1b1SNPrt91GGGyXkfCX08404cf/3F2dtMoFL9xiQW/G0HGfXZ8
UH+Ztc7zO76OgJxNfCARV0X9hmlAp+riDr7o7oASBJs4dzyXDZ//jJ17oQB1
adsQtHAXgNUir9iLo/okoio0Wyl8sLShpauZ6ADrSsXfzsoQ2ZntefUOYPfZ
wccQisJ4ZSoL5kJybdzNiIjtD4YBw+xxWSuqiLxj3+4a7hW1yWjGzxdm6Ocf
DM5ZI56t5OR5kv1i2x4YRluG/8skGCVCZoL1VhRsOTYXxjXhlj+Nw3xjphof
U/6XCeZJtpN1FZvcyB/unsOZa9nQ9fDeKfcRmWAhZwCYo93yS+eIsaKsIgrD
zu5OaQyPA+ufcRvgWE5iu8VNFnvMUm8RzKzup6izCnkjwzguoA8zcv2bDJkW
nlE9jAKE8TQII1TRAvj3AkaiwdW0Vc1JbqfkvAiaOYjLsYE1k+QW5tM5PcOB
YWgUsmdW4WYqBbzXG6KRvodzGEPpMKKBmwcukwCjtLofsKGfbamRUOVC0Gbz
4KYspxGlsh2SugwKaFh9Re7KvXq5N9H+qhS5DQNrRY1YhIUGjBg2RhLLv5kN
PxsYTQ6/t89OboGP7S2EPUkNT3N91uFjmqhMDiPqZ1D7dTj0psCYZuA6hTjW
lf9LnrsoDoKEiN0S7KYi95DoXNkjqSKpOPNvpA2fyS7bYX9G7sZsIjgaS7OH
1l0zHkHusCkoxO/VJlJTBjuqqpkZ6jM87X0wvMiRig8K79xynraEb/xFr68W
8MUUAx1ashcikAMZ5KZ3mNxGlaNcD6Ewztvchz/8wJoMkNmyWT7OdSehtHgn
kuN/XwITSs62k++pe4A0mDAuF+WTGwy+JOUqE66Stw4qJnK6vDdF+X39yRDV
KAxgCADaHya9J4RH4Eolz4hkCCe8Y6/pqaZKMfiGBazS9ZEBDOZdRvf9MKxY
ElykFSqMbnF7Rhwuf+3b1WyZkBGTWQbL2yn5vySBGjf0HqpDrlfKoTei5WlU
SWXWxxRZ632uCvGEdvL79N7qbMlwe1EpB+n2yqvMLDZcEdSH99ghPs7Oe6TH
akkjkMwPEVHRO8AfFucDREgyBQ2hT2NK6yYhT9kRrr/qL3juADJLRIWgV2Wc
JHLVeuCytDssyBwJRrbDL6+ZMSAzl2U4Q3liEAMJq+uvDUfnlJhqk4va14Md
9BM2oEy60KQItizOHO/ZlL12trwXg16CB6ebbUSk+gwZjef3M5egFIrXT3rG
D/SGtUODu7kVMuH2gOPVt6l8tvl5CZ8ifLbgZIJjqXly77K1LUrGYkyF8+fM
Cuusk2zPx6C+3HcAayNhik0eVJbCqQbTT4hYFOF122VaciZNmDJbJq+HuzZ6
MmR75P5HNJwrAbrSWOJjGQBkSDzM4l8dLSHdB5T8SHuwxE36qhMy6XpvJx/U
7PEH8GhllpprUW/19wWzaV0mOWHux3mUEttQPEiTyI5TxqTz8VYWkoakR7iT
pdXTQSghvdLpcILSvx3TkaKlVBde+pNr14gqxdQgR/ypUuTsDv5uQqlMtBE2
jDpf9D+PJCrHzqitFSepWxCZggDZhtNwXiPOlFRWEjpTP2X1QP9DINQK7e02
B8jZAOGdOe/7RZy6zgoJsfAaCKtorQoeaCrXi+M5S6frNngpSim/mGDq6oUw
/cULsEOVBx47AjsaZbIa38YzrtBEHuQdejRXkKZlwvJmVcpsLAmQNqi57Fnl
FY5h5mOg6863PuYs1NxILeHk5Pw/wnY1YwvvDCuWHouZvT6Z0QqsinU9Vnks
j6rJd0hG6QbYFq/6De1Rkpzr0maRDCthyHOuFKBj4AnybPuv03mAzeXMYRy4
ifY5YPqXJUixLHu7Rf5DI22ImkuAN+6nly6kp2TwHIl9OXA6IZc8y2OSBCy0
wjoZghSU9b/KT5+JGyU+pLWPdWRrEY7PjT5957gHYInsJZtw4IHV2bk841j5
3GTcA9zOzzCllIzyDH9HOrlL1G/3ApZlC6JW3zQXVb3jlw9xNbYgZG36IRey
kzm84O62QOqgP5H+DQltVGbx4L+zzIBUETQ/92tIYEibOlhapQHoaTr1SLdX
DHi+c4DZGzcM1uHR+wQmW1BEjC5al5shEDYT0qIVbsgqEX6w9aShGJw+XfMs
PrBoEIknSctKP3cuRkKjH1cL4pUtUd24MdWRn9ZPRKtET6n2zNkJuRK7NpVP
ezvw4e6I74zRmXr6Zk9ylo0ok2MF9pjwoxykP6+xUIIwvvr2stZpzXJKlal9
pOg8FRPFhXvMMi3ETgUJjAhynsEe1aMnde7CiV81p0ZflzJvwKmQ4Xfj43fu
8pDE+BkQuH15bj3zQBqA6FaQ1BaMa+apbzZ1YHTT5RXWMlPdzBCTD9vak+lp
TT0ub7aeXT/shsmr9gLO0SQKNBlqCrbDAGggaUNz1a5BJbzswtqSiEgeIcKG
4kkaLQxLcqoxXhoDceAZWjRfYw9V97myckqrrcY0iFCDnQVfBFQxSFDI/jvY
mwwiRMPKA2ZSV4M9wsbl+GMxRWCy03I0ItW8D2Qr90ADDfRoW0y09caU1ERB
Wz/5I+EB7rEZd3Wd8ClRCcKly5SqokAugtG9tGS6v3xhEsnikBri44Y6nZV/
LrB1ccTnZYTvNEBMqKpRyWv9mzyG6rdIV1HOpcG6KnTlfSQlpe35YHUBC+9+
bSgxRZLC4A56g6Uu9xKdCOZjjzKxua4/Ys/GsOXzWW23rdBVAfocG0wgAwPv
YUqwxOtEjLGjFMxMPysqAklDKaeYsTBiuzkl00CnC70u7QVqDVNdtRj2AEhA
PpynthUYM9OESNc+ezKEv7MvbuAym4Q9iblcg+doTMJUEf00YxdMSdtuR2v+
xRpz0kRdKSCRbUqMjlJ1ztOiyznmC0IRXJxAlCIMEz6h3Kgd1K3QxriW9qrv
MWr/XjejQjL9vAvbKbI0/f5ISlv/u4gJb+McVyZxMF8zs9Ry3+Z0DMMS85td
aBOXoxhpOe6hVU50wFqR+sO/XqA1ha6Q8kfIkTHSCASnfVDij8FNzcGJMBoD
Uf8zxQeoA7/jnVb4b/4bbioaoIFoJzn/7UsA5SsZjcl28Ekr71BZb1IOGMYP
Q9SeDQ/NmryEDmyvh2xsscP2dK1XsFyEOmCLSmAhdh70NEmasO219EOgQLr1
Sjkqko+btRLjq6TYQl7XvvEc/WyTmO9sRbuXXtx2DCHo4Hb/gEuI3ZcwlEsT
Fo2b/WsvbcrmufWd5g5C8SAvGbEkxilOvoEMBiXL9SDxRAZ/EJji44Zjzf/k
SIinajCwVOeAdMfgAyxh4RxISAf3fYTfRr3XV10JMhQ+QzINnUkFnJC5+p5c
t3nk9aza1GG5arFpCgnmYyYJXmY9TV0JEi2mWX/Udt6swaSyPvWYqhJSILMB
zoRh0o+XjNiIGcl3utkof1ILlw7hqitLIU5GyR+xmjEHVYv8oYOZHHRHvaIv
uS0a3jIBMu3d5wazYRV6AklmUULOVpjWzZireI11YvRvQMwG5F9njBmg5hj/
7ELGtANYhh5/AGZs7KdqBn2OT5xsiC2DYYwN6qNTzCx6L4rLQfckdjIvLfDZ
KV4Isv7w4mtdoPXPyZwqE4KVVHoohTgu+6nTAGnPnXaLo71fFfkwhZ7yYoxM
BRRQ+mYsB81UNaw2E0Vay8X5BBlZR3betRrxYIJ8g8ZAWGvm3K3M50ar06r0
uHrMlQfXC1Ol5XyRYREsy/Y8yVhOqGv6FOYrEx1K+tFxSkSgu8sY4tnh2Y6C
JxpmjXQr2Kj/4Urz7v6ZFjSM0VjgLIc4p4QTi4BQCmlG/SyRGzXm95Uoi0+e
gI27xBsrzcDd6eWU9QvD5lrrjuAM5f38MQPMNY+H8Oo7sUbWoMkFPzVPFaCP
W4cjsqjnymKCQHGs2GPbqH1gjiXDqKhXpf0c7uYGeQ/bGlWWZT8V7kuaVD+d
DWVMeqayHzX7OoSAAPMqrmEOX/uZFsUhoHe+YQjsgyHLaeWtq0wRIuzHmjL1
kprlrc+ZZx17s/elVd7TuSphqaYKtfbBODQF1Cg3KnVp770J9Rud580VoM2x
kid3jiTI5wyhXOqDjHzTjoVpBPf8Pewbs885tjnDopsBQlQgiiQKn/ywhOTo
Lug1E2gJFkfRxCZ7XHyLtSw35EZ/lBE5pnNWrnN9nAqWxopp+rhIACDgO6B1
q4fr2HBm8bodGuN0ZuOAGu4nyPsG8Cgl1xdSdjZHiWYz40RpwdaVCuZNG1T6
HUgzGTy85RaAIcI32c7WPGzE//Z+qjMT5AUNEEFMN39awcSo4FwhbSN/x4p8
8C8RDfmJX9x4oYk00yEm4kMBxxVNwQFASpIcXmEcVbm51QvvakLbqFi99ii+
8AIVRtVRCMnwbkjGRZ60GbQt+dRYtRsZfrX0k8dPVJFjfW8HsDX6SFVjjfsy
nGDTS8mzvv2h7jt7ZJhJN4dQl0f6XGxXSFilJ7+wGJ8nwvSTjg+brb+IfcmR
LQePIRpc4FkB39UAjPcn0bK60fTMmWRvWTXVwiclxykCJvsuADZOikqeTdf9
W9ghBTQ/PNaAfOvHv3hSathDapVObTPpH89qqZGLb6gg4/4USMy318THIlp2
o3pyh3UgXmVXK8fyxAq91SY0gW5t7LQ2eSh+pJLr7fy+pw6q2sIR3pRrB75O
0mwwsKYhyf4VFHhSF4wgovvRVtFZ1NWhLcJDj4REoxyBH094WTtUJTj0ULLd
T9KjKfZNPaSa2M/X7/QZ70uzLVv4pcweXe6zaSetQvKLOhExmbq4qRl5+Mp+
IoqFe8DWZXGXtWd7ZNVDbIMH3lalyuDDuFY45UkDCmUekpbOcorS06FqbALq
U7hnCN8N+9K34cOXktOHupn4SThQtZ9RJ2BbTx2XvP8w1Rbuxfw4vC4PFBGF
EH7B3CRPcf9p5w9SjUQn167xzWUu3QktwwIZV4/fLaqQv4lwfDu6dKXIYS8G
6+LmkQCTlCECx1oaE4riVgwfw1ifY8WDwDVr2lWZHjHG6n1/TOXWAJJUCuoh
fqPbKzbGO00dFYybH1X9jNpCF7HjEw2oIT3RY8X5mMC1vXO2xFLm/wslc6D/
XAS2iv8bZ4sVFLB7dPy7uFi2gg05uPMcZlR4Dy+lEqop+Ixn9oVg29YTYywc
y/WjMhpYmydw/62jof4SOkfWi/QyYgw1z58Y9EjMd9bxBU0tl+9cWUJdmhyT
NMuMF1HlJ/MHLsCGCIqeZJwl8EvIzlzLCPLjZ5SQ16BDlZX5/gIJgJy1fkwP
mkns3iMyaYzKETDFO81FbUgHLHDv6mYML/sFuSrfvtCP45N/t9mz7XgzSgJa
JIjXxDXnbkyZAe+ig0D0mjT4xuDSjRA1uDh9z9XXG5jb2RbDv+/LH5rX1XSD
ZTPG84rYDBIyBude1mcrVPRB0bcu9/vlKMIqb7f3dcc4tkV7F7Aw+FVTN0hp
iSLK30MGEIXnQjXEwlHtNijbyq4Gv6ISqJcsZGMtmQDxv+5a8/G8ix6rgXwo
w7dBVZKjdV02EttF49qVm9AtdWuCWRYm/+RlrHVFvIQaaSOmhDeyNejrzrJt
qWX//A0LwsNEhqv0+gnMzGC1VKPJpRYk5RzMzU4D+A6u+O6Zgc41Tg/U7cL/
orHGx1QLGgXNWLIHMBPo936ckRgApW9PMMThBoumhvagvPjTaRHSxhA1dcYC
izIc2tocR34HBtxRnJCPJ2dO5NVn75U1X2lcFsvbzCfvREmFlMt25nxtcxQ7
V4lNhSvAv8SjGZ78+ybf1SKh1mWPO3hGqWzI0PlmZzuY12FS2tEusTZp8Kf8
WOH6U4ErTH/y09kU4O3i6Iwtm7J/837ZjUyJgmD5Nsl5we3D5R90/iYNjQmd
SuL4yMGMUw24hyLCfBSPVbo3o5fCZEV0jsS+MksY8250u7+iLQrkapzUsuM2
XPHgMLe7abx9174XVwrsh4IKZvEMuHieksE6H0v1Md2DCQmpYP+qpK697cVL
8Lb1j4UzvBopAibrUnFqQuKQzAPABG9eLI5rlftyQoleEpp1py5NkoYufu27
94lRqAq2j1UtiF28gOwE362LvhrV5Y2ZewnnVeFJWSq+xWNaJKsIwEjnDBiK
sDD1vTCnNWvS356Cgde6fxpKfVulaXNQOTjNXLkFKuwfw6MnG+E5qfk+Yp/b
2/eKZOSENKd4XC3Vb2e/7J5eJ9+AKwskhnmE1zeUO417nNcvayv4dwAdBJ/H
DJoS2OldvY+RXdnE2wbJxhy9bhNFkV92ZojS6MbG96sLI5qKkzbS8S9/cU0k
85ls1s3l7TIikmogzRx1fyzzetbqW5quWIHtc/9BwczloEX3cdXRAaP2FYAV
vGFgR3cEQnNUVizewo//QTNjXicZl4eTfzQp/przTOAV9rtItKlYCiPESure
2bhZbpp3KZoHw9uIUCw2kcc6/BPec2ePyoTuOT2rh0PqZmQfFJa6ytadd/94
sgVKn52q7yHDbh69jHQn7bdXRkUAcMEQ1kHe1K/MoURUHyjUjc15cPohAUWq
b6/yomBfjFFSzy4uQ9I/BCilghE03IKQ+eIDtBS9PCSaapoExitghxlcZ494
X54l6wbrp8Hdq09kHEneH1uRVPCs6SAi1w3bRdiqO/cIwQQV0askaGwVOcgH
AzLU4HQ5V5cXqrY3v9uojP8IW8BskmvzQ/Cbip6J9LBdT5Vo3ECce0Jz2tdh
XD+FaHoxGK/IEdrKmJ/Qa6yxT0VFGdRFax9zawWWH5H1M5eu5y06SDcP+Ekt
bE5aFZJ/uK2y5TxaVyB1HdRLCArIqkqacGcEMQlney4d/CZAxQwQy0EHF9TX
0kW572fsSuEelK4BA+y/972Amhun1ebXQDHOFnA8clvyeFm04liI0VNwTRe1
MTs4LGkwNSfahO6Oo1jr508ZvR7z8ktHjHuhEuoN6F8KYF02lSXXpEJJkDDm
gm7qGUGhYYGuKSIYuoH3cKIgxz+DuHW1wAvwhUdN4Ip7ufTwcD3O6KAg+4HA
FWfuIrlN+80hKZplULrOwig2vXYTXwnvj/Mz5w/NbVpfI4H6atUfWcxUJ2sl
a+OGDpv7WHp5k3qbuTuUIXVfhTwB0/IZkhDhRpfmuXCBDsk69uV8p4Imd8PN
aP2hJg5g6QYJkCMUULconj11fp2rVRpyMNVf69B6yzA9INGnZEPo4xQ50DjF
NT6UocmPEBegVoytQpnkdZItjBsy8k5G1YVb+zbyYBNEHPABUCEyX4UhNG6+
Jupz1/6JirV1Z7OrKGGX/rVl8qEIiolhVfAzYz60uEhkdQmfFL/eWxntz19u
Iq46x9qUy4ZausIYNaQz6qE+8/6hW6+Cao1dwbS9FEWqPlBsrJQ49Am/wwmx
Zy25uc96/tRLSEXAwm2EUo8gSpkEqaXy4kvQWLvH5V/zc9X6uKPy0ri2vfyx
Tj7NC+uj0ivuVn8ImCHIZjZCV0/IiA5BZSUB4CEqXIJSgyGlaZ1zCxT+/weL
T8ErgqFTxKlG5Ua1iCWQ6FeLK26WsnG3+oiHTgp8ih7JapS5O+Go3yAd46EZ
/meDh++ogZ71jtygbfn8MY2vpxc2aA/HaY3he9gCs92ZGF7C50hqpjjV1L2s
tbGCOXN6tmtsNChCfmp7SZpmZMLL8OEFZgefS44YVeaTtEqUQtfQxjpiOgfY
T6uun1BO/yfX462oj9nO79DwAqyfuul3H2+v7cwJfJubhDK4lwqJF0z+koLn
YULspeEDwWQZv6YTOcce818+oZ0r/IgkVuRCNYcNcVt4nvG/7CLTCwU6vtWT
yzSEexgSzqzbQ03pmM4RWewRHxaasyTrFYJRJ+Gk1kT5N8QOorQfHCcIAwO5
GflV20pgv6NP2UNxS9Zo2N+eeD+IbFKIDPr0WKmeS6vTnEkyboTrjE99tQA7
rpFMOoYH7sMha7/rOBwUkCoqXk3VVKjbGR4F5umXLBsrmc1AzskzBTmtq2P3
UT1lXv+S7Pnl+g1TZB0Y3h5KiCoupAenxB6pa8ZvHyRmRbGa8iTXIS2KTNX6
UZAfYKHfuFRjIZvnCmmFSlLC9ywMCO2fDgj0Ztghz5ongouwuRC3SGqLljhb
GjYcwcy9cLiQF/J9e5OOzmtXiBRHsmtnqdX+G5O4rLGK3dWrbW/tN9uO5xia
UhpPAQ1rjQN/Lm8BPZ9cyaElRFHs2DwCtKwxiJMBsBKSIk0hBR4EAbQcnJ6M
4+AXbjXXwidkcOzWkuvMl87apw7Dvk8vjT6//KzhS1NBdRnx/QTV82G/g4o+
h2Y5DfQFqGVBtEcqtduZu1bhthBYk8PK/oksufFWVMCG4U1ple+W7EPLqJKb
wd0JSCQnPDzPU6W3Agc4dXfi/D4MaJnd+ByigZg6L9YAsBiiRlh5K1aYC7Bm
/a+j0xN/lKAHcf7yBd2Yg0NnQNhdI+6ipLJMZ+xmCO132eH+Bkn6GBjfcPkF
7yBMG3smdtsNFzl0/AqxxDJtsLrWTqilAInrKcW3GTmqA28mthTQPl2eDjLv
aqGUVw/4p+XAxI8/mdlsr1WrC+AazUR/ChUfee/US70359jP5sjatCyJI6Ee
+OzNRHvdneQZoiqTUBZLP3n4guNbmqxS68TvVHhuPqxaXlgh/iaiwz8j/CTB
h1Wk7kioWNPw6rFEdITFMz7ySNIGU6UjdHxRq11ocNGJ0FBnEhay+Iz4mXMw
Q5YVMA98qDTUrAwCh3Nx99bP3/rAlGT0QtjRGwhdZ0rcvZpZYBLbYCOys+0T
hSqE5YejGPdHUBFOWr7nfAlZn/VitdDJoT4xA0IhVnnYdzPZ/oczXHsq6N/x
8so1Gx7iConV4qY3FBZBGb7Zl0apTl1oW+BnDLiRlDE/TY/XGg7J+NNDXiHB
TFIfoU2nYId+MsVfaUaFXTaHP69CGPXXgMLyfcxV4pdoh/6C5S+M3W+XlrX0
uS+eHeKlTPdAR5pfByMPZq4CJ+P/1lVNRmO4jN+s/HfRjdwJkynyoQAzyldA
+j/+Zn6p/xGiLhdIEmfD9PARsZ6tqtrzprktSZs7YVoeHG/8mS9UzgeAS0OS
rr/KPF5f5e0vzmQs9eJrW+jUK1c/4gn9gzIZqjttlnShm/QHa18dLOZCgUev
X9p74J7bVgw1J2jYkIuxIiFSa/X2AtO+AvpGGEyrfmSGvctCUvAvanKISw/p
kqArKRvI+kMEzzdBv8hYnrs3H2DEgizN4Y5E84Kik/u09v5g90ZbARSuxyGD
9KOoccEkkZbLQlvQlPRNOr+94cf0eQTlypf6Ms4DGoqJi6jOl3iQiCQk3YfX
TZEIGJoNg5ArKRSnS0bntqOKWobNPB0eW5mZxRZIHsS7uF/5NLSA44LB4Nn5
SkcwnXKZSQ/h8Q5jqDdIWKqMk52vZPzUoCu8vDosf5Fx5SzMceGUj8cbWNdJ
ctFyBxmVTYQ2mESS0k5ZRt0eo8pFs6P3T1FqOKPpFABTmlHLEkD/u4fIDAe0
YLKS9ZQgOJRVIgZ9dD9EYuTA3AXD5S0K9xQ1EVrC/7pkHfmD4szz2PdpThxP
K+tAa3OaVl34M4oj7pxRUAsIsqXyVueVqzWqcHiBxfOdX6MItUJViMGf21RR
j5Yyd5kIQcA1o1zsbojvalH+0jxpVwzZ2l+hrcwd1VC9WxpwCoQX+0kMeFbp
NAniJmQabpxvln3Gb0dzs0JaaHFhpYlrCc97cbc49EDJHSd9/v+gT5cayFMy
jzrOjZH9snfDk79yFjvbIuypViuHxNVgoNGwXpq1uzMf7eER0zZlJtzgaA2Z
5fwYqqqSUDB3Y4fyQNa0bdlsUdS/8Y9pXCIezGL1vghYt+jUe1ixdQbCZSDc
zGNLPxdeacmmSyeiWs2DbbHE/ck3tQ30fX+6RzF0cCEhlYoHPJ6Sb4XjCJDR
4xnQ6CrP5kvi9ARiL3tmKSqfmnnsn9zAw5N0VnSnDM8IqegLznUd9F5bY7Yp
jp3x7vv/Z1C+3Hs6CVhZ/j1t6E8ELlT71ID1Skm96nvwidB5byK+wheYqX1Y
S88CK2j3PO3qrldYhipOfgNChaGwvWZS8C+pEs2WEbsbSO/9HscnMH/cpy11
EB0rvJh+ajRH7EHPTSlsA1xuuadehKbASNOAZq8viJ7mVM8xkdKr6lrBsVfo
eWxZmOaT2vr6wmD5EVE7PycnEHpQURHJ+TM96eAqKrf3xxTprpnqg/SD/2dv
G4j09pTiC/1Xw9SQOO3uymlzgBf14moATpzM77ClCx1Hj0w7c16380OzTaX7
MRQc77OQbzY28ixXd1DxQV7Yv6zkzMOpB1hIEow8zsnildG1hUQgNWgxDEIj
v1QAEHddrXpUXSkaV/XUD9/7/J2Yct3Rbs9tR5bmvTUHQ7AvuVOfI1ULI2gl
kCKISaaD/0l9EZu6NoRwC9Vr1Bmcetaktgy5yq1Bndsz/rqkZe84KdS+d5fh
Q0ttfPTcF5AHPZmGBsS8+B+TEIwT84VpD9EHA9Y0i2Vn7Oe8zA+Vk/GXT8OC
Y1OJiiV4Srvelq40cyaIDGFkdOQO/FuZn8LausAJo4hjxABjWI21ef1SQLmu
5arEyS8yQp2YnwhzfGdiZL+tNSZoH5vV9gXnTvtYN+g2R1wobrBzQ6bpgzwM
yh0i9FkBT3SGYTf6pYepP68cuaC7Gm7BAcu6z6PGjV/NQMwGiU69X1wE2y6B
I6+aFOD6k5bAUUyKHVoqcm491+hUD+NHTVTBPEk4IdRszHsyRtkmUswKjybi
7gHmdYV5HPTEsHqNScrntOwLio+vzN+eQUQTKQw4x2ak77WisfrNJIfriCOo
dATY6zJp6H8OSat2M2qfAa/jrnJLTMWZKGaEBo2oLxz+qpzjXIUwa1ezLqAN
ESBUBzlhO0Pm2rAOOVf/6j8LQPmXCyNev8/najdIdtb9iaTeCIAsV3oYQa7g
vf0ncxdLYu4U5Ho2hlrZ4vKUxXHOz6aXR8jZkTqY78MpzkzGejqOFngb21xo
IBmZm4qdwD75krvBz6uUHZHie0aIklWCqK5bOHRzLOmsmrQI9fkHLsmBzX4Y
+XgX8atdzB/W6RSVgoujsu8Alcxn3tSk+PSRaIkHRXGnhGHdfpJDJCL2u+QH
Bb/pz2zxYFZ0Vg+rymKISbRxIw6Z0jZGpqVGjLuvoLHS9t1zWvxRLDix25Mw
arb6MZ7heaKCeJKKVuvL/LqVYud9EQhqzsO2nNN6z1whE7W21Ep3pTYWKT3f
mbrvPbCW9YoQZzfII+lA5cTh+DwfEA4B6cIoLz+buGQbfeNXm/KKFdGwPk9a
Q9RRxLpfFVZah3tW5immZPaTNX+ssxQfUDqfybPXtkAETubllEUCueHoOS4o
oxvy1cZdDq0MZM0tPFsT8bROTD5uUmAljJBEAUPhNOaKIt2VS3yHvBN/VUca
0OK/ajExOwvfKzvav430lTbizdFIpA0/DMcv3vR3HtfjU7tjYsRRXGGfh2D+
9nlb+ApSrpSrgQJyu9ubzYdFVrHFaIZ3HKV0SBbodjnyjZD5gmlFP0JSSkRi
2oBlwOpotPpmf0LRP/fDTen2dQGBlkc2wv7mw/MKzPHq0VoNAue6fxcRlaNQ
inU3gJZhhHNNWkTl1SRPTaKB0Wn2CN+8yWn0TbX6Kz7QwYI4S81qGouFHMiH
lG32iDsMz5f6AVmyiq2wRm0pYakYFv6p03MehGB7TnS9Es9jk1Xewt/tZjrZ
wKRgQDp7sfWfkrifX09Mzzy0HmAofHrTkXDOxFw2vDO0zFJcwiC47IF59B4t
eoU2uyolK11HZdDLO9ZhoR2yADqNzkn4nK8I2urrtCNR8QldyaOldZjc35K7
JnS88+QYjKZvCNWd/btGg9B2jmFeiazl62GqYKTiufwiF3Am8+n974ZZehy0
stuFH5bVzA+cvA0jjiEofQUbwNsmJVOwBgtiX2shBXTUeYNtULjIWxaK9K2k
iUZbpR4FlXkKrm+cdsopjSbo6YH3VcYB6yR1PazjOeXhxpbiOUcjWzsz81kk
LaoHYSpiNxjk3ATd4fCTVNVRoPdby/MBUmffxfXb7mOc9BARsF9AH9tMKRfC
TUorCTC4ZD1HJBInBiZZ0bwaPVyGMJvGTA2fUUwyLEJzkUcTCzpHLPsWPAvC
y1kWWwHaoet0smw9RZc8MFIa/8/NgDbWL/wQtClpwJ4F/8ouR2lwOEkjJ3u1
XgUiwRlPm4LFO3tvIcr2mYB5QR06JKTfjJRdWLJ2b9B/jqR+cHyXwIkVGAw7
cL6hBY27Q77Bgna/0usXERWsEwGOmd0U52g/CCsJBj5m6VCBlSsTLR173eV5
x8tRbEc5l9WPVtcTr54CQYOqjzjbRTqP2kh4Rirvy7T6+ikjU44ClqSCGCI7
sddk4vYRC49R8X/ijmMEIksZDJrQDv4YBXCxY4xKFO0PKZEG6xu9eZ5MNeds
GAxUV181gM+89feAfAcvhJjdoMGclcFGcOLsMGVvgFfKePv80mtIv8JSvRhp
2S0iEhQdL5EdOIEYcj2jz8gvmr4sPraZfhzlol9zNKkkRP/2QThxkVKcqmrH
HE6oEDOd5r7Kx8xm2eawNnyqWdlS4+hWHm9Dfm5LaOg2icnau76uSjLKK4O/
sQ0TXLTzalo1YOJvktfamrMlMkUpras66b+1A7kZR4M9Ns6ohORC/3pD6rJA
k6HosHfxNMEArdK6J1OjlleFz2iEjwkCWH8evDuN4/AEP/W6vRcJoViqResv
7NbCYnuZdM4ahqaHSYajmTg8byMyMcTqmgreI8rmUEZvZv2xa8ORGkqGBTjc
DFwaqkmp/sgB3/vGVZvQuMJj34QwozvH3Yb3ec031U+rcE37lIrr0zGC+qtc
mwOmNVVad32Hd6hq16rsOkYOvBFegHn4qbCJIlMrn2slNezwZwnjLQDO5HoO
S5jnuY0d8hW883PnjHhRvqHtsn5MCb3fu0WQy16mmOGHCwwWITZiXlzE5EbS
LwQ+a7TJFxvtj21y6u2FsI05U5kNO4AU+li0hsQ93w/rpYRZwI5NEf1CtXbY
0T8kj3IbqOEKqTRoC2k0qjH+Puri10OOZ7Xka7nH9VQbucYkWw+B05Iztvid
6cq6LEVfu16/b0NUcAuNRYg/74ecPoEYXFkS4RHtne6utbiDcA8t3gaBiLQt
MsOp3FfeXEa1ye6lieRMZTNHY+LSFOVF5KcVGBtSYRni44QJi9Vb0SHdx2qf
aX/K0AR/s/H5B3a6bUfCm6EbAIFoMWn5Kul7S+F+2Z486/z4Gi5I1jpynSx3
TfdteH1Yg67ZpadCxlzLDj8NWQwQeb+6rZO4wXDmQVV8s44mcsHzhQEkGppA
xWKv9GAx96hz2OJZzgTU+RxfiEC1hySSESfstbdlEpu9oe16FmLSnrzok10i
Gn6NYfJ102N6yV8bsIYmKcKxO9VDFNB6DWcSpS0K6NPPr44wOiLo8G0dfeMO
9GK9H9wPq9L9DTsW1gJnMEy19tecdwGD5QuL+PrRQImXLh+zsDnHWCijTYmT
NywCfO8OJKN9+jOzEfqkuUXfLrI+lQIogFMDikwv5fepHqN08FL6/UnVqu8p
Wwc3aSVn+/vHfgm3LhCvm15S363jLrb6L2fpRsPOU6+q77PrB0vjwHx9zwZJ
mhQCPr4AMmsSraP6klqkfIx5uEelkNjPr59lqXvvOYzPcg7lfTviIqzncReh
xhxmjNVZzkPH2A4VHO53BDzhoXzyTTcFUDSYL3ycHqjanOQ/f7XOH9FVqXY+
NnO01X9h76AjB6YzNFhqEJxI6dOlbs+7fOux+kCNsTqtkcbBnlq5KK+imZzS
NveI+UozzZYA99Ke+AOj1B44uRu+zMIw0QoA7umVQoxHyrTKeL41J2JR9F1o
sTOrowKHQ3RdT9Lab9xySiQa0GucY5b6LAB0C/T/wnD/wmK+JveIGxHxYmRl
LaYwaucSVnFb5ICIBe3facojdgLJY/pBRwCm+ecrUxFa6LqusHPod3/3tZDk
T27DRrbaYcw9mLk6pZECmhzbZfhsIWb9FI530J1XH5WzF5pA5Pv7C09LmPsb
UoaFpdAfait2Srwy+A00lfcPz0zXbGXOxh8kqs66u3u7v32uQf9zvR3GDgEE
oTGeNvc093mE8YwvDx8GGdlC4VJlg4zlBJC1KWh/4vuuHpVmER8ELVvWEKzB
nVRENKobcWJvFpHGu10vIahxjki0OARqbfI2tGe0vF1DmYfWgZtTKuEFpRBq
JsLliuJ2tKkr65T23566+/UorUeY/N13A4uTuU3kDViCsBtbpzciJUy9iqpB
GKqXH5b9hT2dlN9xIhz56hWNVSM14dqpnGYAUBG0Cbq6nJILTVso1nkJoZo7
LGxeWtWKsv4kyEMwYCYZ2O5bvp8w/gpZ174szfmGpbdDlH+A2YLXpRi+rys/
NatMOrPfu/Uwuk5ZWi8LUHJB56tuo+kWC3Y7JkLDfhODHEfWKHpY2JzPjmxB
/ucfgyDXYH2AuU6gvu3DgF9gh85eYhQz7mEgoPXF5GeYzskVBViI92lZxLCC
20+reNFQojsu1xrJQPe4PHKwmt+vpzlwPe3EMpQJusnBPPKejg4ir/ZbJfnu
QpZVtuta46yqnyJKTGKUxcoNmjxDePWGG6wQBvyh9tzCJfVwEII4EA+F42kC
Uvf7rCqp4dKca0mnsuTRc9uzv0uhR840B/0wQid4jpgKqpmJMZkYufwm/FYE
w70k5an7l9p99HAORL8dZrAUQL1NVhMCqjdEtbP+/8GJY9wpYY6yvwcBcDpS
EI1BTt3pVMqULtZz63mOfzZCs662MaoGM343TFZRy8yFMVZtJA0sQnBw6Xvn
Z5qz3IrzWAN8kq0U0oF/qd6a5ijCSnWfC6KYYtolFe5gLhWwbGN3OQpKjXIP
XgwkL/b/khvwS2w5OzVzMaLFBwstLq/tB/pbu76PfVyIMkAlpRY4RBwIfbtv
rXUYN4HobDNOS03tMNtO8mpQ1iGLRXH35naOLEhh6CSdNfnYttgdOIWF+DZ5
Iz1OXGFgNEZn5B8OqO1TXqW6x1l+44Op8JZ48q42M1vJMckt3lqPIyv4g7dI
JAya1ElZ+G2oDYXVEL2N0yh31NbV88nMpBYYLky68Cu9q43CJu4PATqcvCDh
aR8dLtUdNY8j30RiCODgMHZICthgBMiG0/M7pnTF4xMBzhZdQPb6trguonw1
jv1oPfUoxkvLMOjLKtp9RHo+UePGy7u3alhW/Lq55Qjou8VzCqoXalrmas/d
Objozce2YlRrvupcZ9Z56FDpeKN+Z7kPoz3p/XCPcw8cExzXDXHALzc8ch01
yO5OZNa8x0XtWUX55xQzinB45Tqk5q9AaQID9tsfMbYHlVgSzLROqqlRSoSz
mAr7f7XRtLOaTRqK2GToIYQY0R1wp0o4blue+QG9TmgUfutWNKCc+0fDmwZF
K43RjEvOm7RQFvklctP9v9+oqf8S0XDbDpn4yUwTzKnLGPJkuHLHI4GxtlWN
UE5K3CdI1zt6GOxY5TEV2CjuMqSjHbhMGwVF+esnIuVwqhLb6y4xxZtQ4GGB
glp2TApaA95SBZktypzkF578NtIzK0Wi//cFIolgaNS9f3KoDoAijAVEs4GJ
2H0ElzgWbyPs2ORKx6TPJPQS6UI6budfLQV2YKRQ9aJVqLYD71wbPt+g843x
47AhMeqkwHe3loVflXDnZH2pgaFMg0cbwgr8sE02GEX3znJPzaP98la4bo/t
5oCDIEwPtAYDWTXdkBFOEEjlIepCCSLSMYyfLshxdWGGtSLPDACOAFWXsnPy
WMYBXJGC14h0JjAz4Jefgi0k7iOd0p0FBcrjaGhhJ817sXFlJaOcCJ/dY1PD
G6wu0P1FsiWEDZujnDQkSo5cF3mBii7AFyhk8u3b8g1RffcMIm9OXJBzKtNb
kvh9axi8+PkxNZnoruhL3KRdrs5j/VPSeo8tdZAkHeoZsmaywqRjwvH348K1
s3i30PA3V6Mw1Q01X8WCLWrNwK6r/hjelnOBMKWRURem8bqaZctofYJQCGJZ
o9/5qQ9U0G60zBP99tRuE6J833SVNNsy+p/OTlW12RuoD5GlrnQzv+hJXUf1
726FqSjjrRXE523DN8x1ct+WwH7SOvfTZDiMw5ZU9ACkJLE4Ijsermk914ON
7DzgK8yqWHOJyZG/lCkwFvzXv5RIbe3mJ+Waq7kvAWOYXaXsz+8dItjoclZc
MCr6lHtskmImTKDE1HWdDKq1Et+P8jBNZpbfyHSjA1lYcE+37ivl3r3NgrTO
IRzwUweNkfSkEGkwa5vH8km+/uCUq4pYxAQR2RGT7uKSNxQsipaxpnloxYQK
4rPDI7JRb9x8onTqqtvg91nEboFhrd+g3ZU4xNnj+7xKGn1c3r/tCRhyXhnY
SfJOlJg2RQbI4jp/Q/cWmCJX1vqz5Uq3rWq4C1P/xPNB6hh/P9KMJJASD5cS
Wzag3WY1g/YiUqZ3QHbolhj1ia0YqulEm7hUSZq99kvBiIEggtHvMW7idjTM
ez1qlZH5ILyAk/ELKIZHdVrGI+iNowjAsMj+YeXY0YH7nmcSWjU1gIMnr8F/
d1W0h7nLynGoCCWx0bf9rT2jS5KllUSA7PsCj/opLLxB8USEOAYsFMyo60ip
l+VGetVmim2X8nP71953UhkmeZHQVC8cOp9dzxj6EUDi3Xo1b03bskLctG4U
GNKoJLXPsedwIQWJS/IJQjgBS/cl8k2A0zG1GVrif0O92I2tFF4zRezJTDEL
RVO7E0C8srXupxS9e/eFho0bl1GsucKeF+/m2Wnk/oCutjbC/m2L2a2cXYqh
nWZoxOwg3uATHaoojo3vs6t8cIspMBhL9zreCORqcbltBxTBwCzDhZmd08kv
fp3k7yl63E1VrnMcYGn3hLPX5h7lFATRiXG4Slhxb88mJLS/GNd+vItmVE1h
aU/aUPlo9BWF+TD6PY7TS7nbMLW+XAcbYBFbPfSRjg8a8u5u+xc7838J6Eb7
B57xXBajErcnEmA/5+ktl7juenZg21wpCg909LCSSZqrOuIVuwp5UcpyFE9g
I2Lp0HUfq7HHJkLGBLMLwla+EfXtcn0dHfkfkMe3hsoar4IuMqEcQLk3NzVA
MIzeirYj4ZB8tCaC71QwI+fnqkQDUcalsNnw+qTZ2Oe31/mD4ANvVUfSDkjL
q1GMnJLk9zaGr4gNc+H2yf4mLpUi4fyLiUxvI93cTbw1XXfgvDq25SuU8x8X
AAxSOmISqk1y8umeii9O3dUA2rt9W9uJCqWPQJqNQerulN7so97yCIFctI6E
nVoNuBpUKhBYTSBXzNU+LaiRgmvu1K2hGZpNviiwwvqxmOMlROMwv+1C9cCl
QkLrHJ6gdKn6q5tQyppwl4hEWRMswGK+GiHj5gPxJ5JduQChDlUAVgTPQYM4
kEqR3Bh2NPptHnnSQ3Hj01eEjvdVOYNnbq+ea6zqD2QLeQb6mtSL9PwsBq6c
8KCf0jfqHEWsuVzEV6Okc0TKDZ/5yBOt7p0GRh/M1SBsjJHK2OWex6zrLva5
qi2mxracvT+WqDeODOGXlzefW+ThomTfhkXlIEX24gZOD+TvX2bjc7gX7408
tVwHgICCVwdVqGRT8QA9cCyi356Kc8hP4+FaKflXGoT2OI5sw0W7UvAR0J1I
vXuORiqcEibLb9NlEDzECWEdUx2psg4m4e98dRmNXiUVeoyQZ28jB8PHvNgG
I8BOJI/g5EEnaZiITttZlmTbo9yqgxAxiHaqygnFVbMQtDCy33QOlGXeHdHq
eqakXOg6g4s4iS4+SmqVLYz5GqOzh/GZL0o0tc37lpMpgn7M6F4ALrUFpyTp
Q2HdKltKS5aN30McPoCYqAJhqeLR3t+yFJ+ZCDKmDvSHQtoPprAC4UGzoIiG
1QuQh2YQWHkeoP1C/9UiJFhW7RdUVCS2RWmKLydB0MWbUZfYFcBYJi6feX36
j666aGaWmSpkLu0fzPcaiaII6ZzsKIKFNCiGs5ggcTGgDQ2vv5trhXZwcW1q
raVwVaCocjz9pqwT8mRAW/cmCMOtPUfXvOh4KSFdbaQLsNi7aKCy4g9uF6i+
fuWJO0pVugLTZsyAq0I0RWg9t5kahgDsOsCPNlRBDG7i29v19AzGibdhxEE4
vrJOb8TDAesIoFtthwMvr2htLixgtINvbiMhS967kz8IXy80gkYwHhSyopP2
VH48TIPLEXtv0TXo2+Eh3cxtNDAp6DSTn3kAxhCp2hJ6w61mBhpmoal0oNN2
0uuAY7lxKmXZlXxqsCtJ0ZqH1Uz2/hkbvB+yF2SzyQkQXGu+xBilZnSTYF6K
HP5z0BX5Tsdj57u8UphZM3P5NEYGWIoQqZmrfphaWS7/cUn6qIehF6wQzvxC
+6o6AQJ+HvUP10HgFQxP3dVUGGgM1OiK+r56bmXESWdk2K4g+j1PivMRL3El
7zJVHu8t5tRoM+3/1ityHs5QPkM73q47mUw9gbE1z1KnbDUrx+pGfnVxatWV
PI7BG+qPSewUqAYFsL2j6mpko4sDMmZCwYK8nhTcxeHWY3ws5RUYx9QaxWX3
VyZ+qXi8lsIKSDoauy4bSc7ZXpskSgJS+vsWkPLx2LvaEKy18Gd5ZQpqGTmb
gaiQuOOKjFzLlfgzMY/ag8ZKjjrKf9JfLE0Bw+xbRW7LNuQ0HatlGFswlsrp
8l0M5yIowtbXGTI1eGjm9NqaFrHTwQvDev7Bv6UATwr8QnDaIwPNfc7rsssf
D8kc3UATlP2gefQtA39paR9a5uHR6PIPy/+V5Kql4nZtjgWSTUmVY/NxtTlL
p0eBQXd0C6DS672ilxnwazeM1HgB63QBjxeKUkGqh37FGBGHogJ4c48iOCIQ
gnN2Z+c9ohoIAYQlCQyPoGf3DKmUTdHYOmXK/hNoRWjdLGRoI1mh9iPKygTg
PZ/hnuNGB2OmI3aa9SrvKI9AxLfwoy/21iM4wUsUmNkalSupbzZVzo6SRNiQ
sa77bBBI6+WqorFKFRP2HqQtheGmp6o7jRMOhhBoXe40WbrPQbOrK5puhEga
sK8gZRsi0oOQfbS8UibZc/OzrG82F6IqBCb+7lpgh/V0FD8WDWcpSUKu8VOA
1iS8pYJg3ncw13KHJMZ35CqX6ILn8+5ExK+rXSm03oelvU7SZyse8roUEfUD
UJSis9pVQEFhxR6XDptop0hYkuZkHdGqoxUOgIYgG2psQJgXrxUxsRygmld8
j9gPeZhFuRBT7tVVxK9QNGYR5ZXiBVrkL1IRDkdGBc/tdcEqL/sZvoUBVai7
OxFSHkYzLKq2VNjCMAIK6F/dmmLvzkyGAP9jfpTyZBByYZX57dgOlgMEIvyU
SXi7aARLpH9out35ksAjbEAGkBktF5dhneQJ/au62RXGp15ey8Ap2ogSKYIl
AlM9BCYulLG/S+KQ8l8HBSTvJ4Pwn++ZjWAweV54GV1TNfPQpaiIT9HP9BTf
dJ9RCW0x3nUFgIVlvnV/qfGcZGO3xrZ4HcFCNWSbWyyStLAHQjNiJL5dy0ti
YGOK6wmAa623bwbHXC1YGGGlQuHxSVTuOlti9E4nUeqzA8kEkRCJTZYwLwES
y4N/gkCS5S0A172dG81mvZR3ghgfMTVwERucTCKqWkpzAlBlZIlh6DJVPguX
a2POHsvrp0SKG6BVS0ucKfWVOd/TeQLbIht98vZGodZuswAMMfU4sTf/pVEs
l/iSd5VrhOhoOo3CdMAZ0GA53Pbte6jAmRSfAvGO4BUyMezxi+/2YNMmALBz
PkbVzZD2yyPxqdZW48BsboZoz6fulWfxzWKiBAw67u6WnpVSSXHmsP9Tlgvd
JdEObFnFNBTQvSpCOAW6BuN7eh0Tihve288KfhQD2uh6L4AzUGDfViZlmC4X
TY1AhgtL9ZB0W37jbABtrXxcYcsetnb7T354095iS2brVyufXhda3F7aCmTe
sKcmbCbzdhohEQtmoCxt+rdROMlV4xqcSPf21txA7Zmpyy9PcVF3rNotFjpg
oqh+liBIBluHNx0KEWXgBemF3fFjpuXzTiBRS4tBZOK+YWKSjEjTrohsPnU2
+oaFHejVZmtMnPHpr8qB7PysorynN8cvyPEsaNy2Fd/cOv6U2XtIWmZGb6SE
4fwPX1rdc9mdzQ4Vcm87LF8xYvhnrWqpPDPw+xTKfw7bGPfswdXy95mtGTCt
XCrATt2GEsqxZOscfKDcDh9TuzsSh1wZD53xHMQJoeylGqC2278J8DYBn6QQ
2BIeJRo28kdDD+ZIDL6ROkwjrzS7D1kMFdTNVSiSluFrNqYDqt7rdOrOHVVC
GWBJPMVErsTaT+wa30V/pmBjNRiPmsGgNUuGRBswjToVSm+ara3FcYTRQuX/
i/IO30xIekm/ofz69oD58StAaBMdL3E8FRqcHDS6xt5i06GEpMCCApxilLll
TKk4brQLagjr7ftPEoD00kkzFSNIith6ql9PyVk8jaDTkUVbeww8zkozcZ70
aYGJ1W1mB7R47YVG8X1ys9oaAa4cRr+8ODcaTkN3YcrS7w0p5rSI/1cldUev
52d3Xm6aNR9EHhxwMmJSE1mdcWpEfabRg9zqJY6Ej8E8Qb0xxz7ps1uJqjhW
YYEY1WnUieLcta9pyHdhBq3OGWf0gX0SX0HTcj7tWNg5CHe8+QKitp2tNO17
WQfqmZxFIb8ICrcmd6UOlGqSdu+YBIWMF0D8gSxg2fz9+fGgORORUBCVTuiN
9RiNWwcT3ySpLIJxIXf5mgcEbOI227cvyRI0AB2bTVUCcEd7T67HBjM8OPDf
EpdlP9ukAZCiBKqGsT9yGr0QP3H90qLkB/fvg92NTMJTau4S0dphIUIj+uz8
9cl4zPDJfZi0lqYVmq8ISqIghTSeTDWOdKpRE0VP7lpvd5P/xACG5hSV/tc+
s6ERqkkEAgCnLlbKsPpx7BZUpcbp3GNxEFcmvcfMS4zcvUXCP4V9uHFVOQqX
Tl0nCN8zerPXfzS4C+uOW2w7lvij6y9UVm4DNs7U+ZEJpyPSi8Fh4YVEmyjQ
pbwklAgN0pBgt1wOnIGAx3vQF0zQCmZTbMo+cEXLtiFaGd64R9cWxE3HMk69
LZI1bDUZt+NxZe2oBOL5cjqsNldRK0FGmXZT3Pk3VrJTzgq776YLCbdsUgod
3JIKHXQkaWjqRo9os6IVWGzfFx3tJ0GFKK2espfNIicY6b9XVMN7LCJySa4z
qFs8fhQo7Bz9XM+O167CqhU29t2NzPQQ63Y5ZR9vqCI+WOZSJIHjul+mQrbk
Yz1nXHYKIOAilRb7Zdx3eVsIX5FX4pg5cCTeixyILcJgc8qhtoo992KsL4qX
uJBFLsUUbElpEdQKzlhNl5NRog7Xo1RRy+Pw2m81TvJmF0YwsHqo9cE8+vnm
hgq0wloScCDXU0RLG6GXhScr0ImLck0DCHU5Ndg11gngJ7dZ71d3daxJCKnH
ttwHEHUfkeXA/PZobzi1+a2t57GQXE63ffe1T2CiRkVB27FJ23ogJcLgqcxl
aEuxBrmJwfT5GYUi54ipI4XreZMu5fe1BiAPEyEUBH9XKBl3tR9Ivci+CMBl
yThPbdBXUFHQ8pDWXTYVr6cv9+MNWGqVWLZEZqBx8wslZchZqB3dMKjUhp1m
5bzR2n1aZb7f1zD9OBClaUo6UENDBnAzIahKBGYdAnUJZfdVNS5uI92rAnEd
oQClARj7CNKdhhdXWoY9E4mhEXra065m5LYQZd6MfvdKxZdHqHrUJhOlRe/d
Vn9io9JxTz/i64YRRERe+yeuNRixFCKvBm/eMx/5xzOoHIaT+JIX/KPSh9jn
l9wwzpTAwuCuJPlifj7Whk7Z/UlQT4FjmdbCX9T6hb5oScVB8olWWyUdQ2cM
mpZT6Mj6G8R8mIV+WhW8kHHLlnPMJ9j7Ytk03nLHYOvPc/bzhxMnEJ4BnaUB
2y32ivYJHl1eTM7moVlbKbGZtULrgxYMry7734UThI9x/Q7zzPvS2yVox4uX
ABrnlOk3dRRRHfGKWTlfqt/5PnKanVZSinuPGC6JJJUvlTrkKU5/3ibWroVj
+qU0pNZZ85j3Ppycy50mXwupMth5knwNsbAnOBbpX1T2jILJXQ0nSCagEYMN
pZNP7kd3zEP+fCFUmG5fc5QlsoLXwPpO01IlRcNax3wqtG42oo/w58XLAMfz
A+/FLnqfCNnPF43ADI3Bw3LJ3hjCEryWSx3zA3uM+ohRYX7zre+EeK3fRbJx
0wo3Ga7SsBn2SqSNtOhOR1V6p71zD9eGTp1vmPDRf9aB5wbREybmHZ6TWKaB
DlA8fjH85XSJ1NkucErAvIk0IxMshuoueLD0NCPfdY4AWJX04/C5cYYOi5W0
9TOSvZyM6l0/g+VGC8H1ohYUzJUshL4AzoUpU4+ghq78z1/Z6uCmhFboUr71
FV2IcAdmYzqU88PiGLbDDZWjX982+QIC+h/olE/Sl7geLyu3VW6tLlyyaoUG
n9U7x77ehAJwf3BKUgcRQd9CqMImW3ZW5o8gnULwxCnSxzRdD84oH98scIGc
rvsMlLUeJnqZzr1W2yw6Kue0V01iNFAI5fkCRnVE68VcvXFafR7yG565Q/S0
v/1sJoQ1NExHSa3MPpdpcsiyLooFyJrmxSdSfI4dj5IyHVcIy1NpdF3FBrbj
XjwX51e4q+liKgSblI7ISbfOEbYnP75col64bYz65Ll4ryje6c6y9+aOtpLL
6oloPkYmVmYHkpxmwZZUqFzaVe94gO2MohASc6Wz95kHmF8LbRdnfH+bvDVP
J/yczR1om84nzxHuyip7gYyceUBuCrZKBNLAv0G6V2vEAuVKJIv6aCOQuGE5
0O0uzQPLVotevc3cUICqeesd3JQiX/b+wZwUZnK6F2BwouRDRfkKkjs/elWk
x7Naox4TofDtB/ZLQpar59wjyBg62zVPzwcMt+R3W+zYECHBLnO2kgdljGUN
z3iMP/ENCfl1VFSA5dNVb+P5naOPzpytDz1w7wQ8mdrlpc6cWXPXo/GhDDMy
N1xylUWspfflmAk+5xfPmsnbo+JfgKJisNi4nVyWxrHPKSIu7iEQ3sVdNZTn
dT2wySbiHFB6icXalCD4al1e9zncF+VMW7mqkWpJK0KYlbNoNwDSownQnuUF
DzjGKgT647qmNAkWeswduhZrND3B2Dp4cukRtxFl91hf5P/AiaJuVOO3F7X8
1TONptr5bZ4fvaMWlSsXKh+60z4SLnZda+44lpJ2mJjyQhq3eGwmUo6kNeXp
HW87ewT3F3lKw1Czrrhg6VDgUwE4QQzhQuiE1ujwbVaAHC3IL2fLlzOe58q3
o3rIH8IQ6juoNqGohCbsyV6A0fOqPZVEDlPHxNqxagxx1u4H1MkDURWFnOvf
AP5pEn5o+VjuKfzJwcqQw8Zh9GAiCIS47c1fr9OcikndMGPbsrxSPsXKXcjF
hpkqQ6sMbFe/shLSgVJD1qt0rYiri1QF+0h9+uAAwJ8qKmcEkdhN4eKB/+Xv
41SBMSp3N2Jj+hKOPf6qEKBnYqXBDiiHXheQnOx9YdhkI0EcCDzIGFmWaeeZ
iJ4U67WY8Argutj3See00QRL1aGOl1nPbp2nxBFv1k614oTs4HlqoRKadC2n
lBa6KZDP8WmuXninrbufeVwN6TgK9j1LgAwyosTCaS44JXuzVwzj9mm9LbMP
mdBHhRm8Dn8lH5JFMMDjPkSFpmuaXvjC5RiWFx7nnkoLc1I5Kg0jDwWMphLR
dNPDludIjsiFil/YJrHV2jcucDj5nWoCOk2JwVsWriJ1euDnnqTNwPJfOk68
CgSxLBVxIPjAk3CbDjF823h2arT/cEVJS3VohcHDcg1o963IrQCFh061WAJC
vb2IuzET9UFEFyiughsTDZEuB4TapH+rLTkf/RHZ4Dbn6UF1m7PhhbofQRtJ
IadOsQFNHqy3J8TGiZZyGmEUCJzmhuNGG7396r+FCA+fpJ86j2gLYjccGDAE
Dkwsxn/VMJXOi+TesGkqOGjq7YImw9KrWa3jZ4NAjiY86+JxVS1ILtnYdi6R
VR0mLv1ao+p1GL6Mi47ZsJECD6gv1uc7fLjyFxjywVbptaJiW+KGszKKHOp7
ReXaqUmxkzIuc12y0xtopVw9P/NI01+tsTCkX3AIo02D/6YZlpLfBfSRDzdq
WU+wUTQrROgboI5ZKYCEUeyVMoChduA07ADwmiFpUZ+W26J89jn8/lOCYRWm
QTtgt0+arzy05dq3hPxHQSr84852FszDE/weqeFTDrmhN36KWJj4jFCX3ZX5
sz6B1R0Ir9oMOnhiAolTESXcBEOL/50UmY189Qvd05i9TTPnYilzksUwOT0d
WbaOwBHHH1g74hVncnXjMfvqg8h6CV9u5yX2kaPTA2QY1jq0Tp0m4k5gW3JE
oCDKMK3MY2M5CBcVAH84xBl/O4+XPLD1UUWc1l6oyEbSi6WANr9g59tIzMQj
Kbpd9uJKLuD/fpUBGTcQkR6NDvS3MWTpSSWSzfcwEtx50tZSm+kVJqFKf1Xs
8erX/yCB4+ZVFzguJ+ll2o9F5SEv/CjUSCYKhzlxR0MFLb2UmLLLLmave0Hj
oUeT2hb6juF5732+XQGy7mAlrJeUGIyULqL1AyMxNIjnveCnog2EDwlEF5Ql
uHjhpRchJzgBBFsxHg777svhxQMStXj+CL5ku61+fT/lf1sNg4OHxujty9Cv
sMsldL3H9aQThHIItEj0dwZxXvHx5bKmdG9vQcrZZdUM2bShPwgfI995fCMF
ZGKoCPi1rtzsZzau7FvNLQyiM5CaRYBVYbQ7bWVO3ov7zHYiNNqDQ2fYQmjI
lGxfxKsUDzTZfwJS5jOtmpS62s9bQ4i3mGnU9K9xTDLdBWk51u3VQ6nztTAt
v6D64t7bz/IfOj5mcCze1klhb2/WCqvHG9Hcxr9tjCDRXtIvZrF6jQ9joUcc
INAZmWDn/b4x7FJ7dvUcM9vj9fONYDBkvRwohd+JvxI8snaorICXdsxcfdn5
MImgujs3GQmX/dCFSHwI09ACVhwtExInOeidErfOKuuVDqhNYiVLNp6pYNoa
xLC2N6UA8i1cIkcsYtfCwmOO1LlPF8OpyoY+1oJI618As3gWtvG98Vt3+fyN
/uG2+FoxjP6KvBrIxO54f70sXRAyg+Ul60wNnulb9SGTJzUZCdM+9gQv6RHW
eE8rz8KNANVJQ0VIAvbDUGd7Szh32ATJ14tMY8xIvR6LturuY44C6ql2NB3e
dYIuiyDr5vN9QNAT/GwG07dAxTEHjSFIzxoucNFdctJSpJcx/b3C94BJgutk
j3V5DO8QK9Jj1ZhS8LVT9SUcnlmpbfXqpd4uWvT+ff4mP3uCaA0jX0ugtmi4
mmEHg1s2LBA3IL6H897Fi3l7NGr3afkcPvuKG57dNhrnrWyyy47pSl+vb9Rb
ACPTCU1xhxtRz4dFlYvF9sIVYy+m+rn8UfGrOzpBGGJhpyorfgrbwL046P6D
5Zk5UsaoY/vAlPN3MPOXFbyNmZvKr/I4n9hv/6WyOrPEl+is+ayOfOZpKIHb
EoEvp3D5sMQsi9iTs5sWHW1DE3USjzL+YBdGZLx06FzDTT1pyQ8oZ9xfDH1q
DGCGCCD/96zDUQ75z7NqJD3D0h9TAygV7+W1uFR/54HZcAaj5HW4lkzEPDUj
UeYzzeVFD+kcRcW297EGNzhXIn27C6YoqPWJxCCGTAldl1u+kMSNnx6BOHFW
U/qQCbakZU1vKcasNhYwbiulpLLf4mAhP3qNtWXD0MMV7BvFr6dAcfrhvIjc
GZsxSiEPx+5hUcAezxpPLifgVy4I50iUKMgJaTmJUpvWKMLddB349kJjs+jX
gq1haegwFehtO5JFRv0pkh0WzXRY4NbmBVFO2l0Rvqhtdm4aMaopT5SzYBSp
sj7uex5AsburaZ5LpfK8obutaNHpZ+zdJe9FELleVkvTzwpZropYWKde0Gwe
ecc6tUnFZFw8IHiIwZuRseEB0w8tbCPrJ+VvJ+2HpkeSki7K0Aj66sBD3R+G
KldUHLJnzqSgQLC8PkHKrQZ6UkswgVKHXev+S69gIkrnjAMicdY/zyksfou9
ImJgqOJylC5DeeimKBI25wifGBVUFRx5gsTEYY8Y/Q8/J35rU9gOJ6IByEGp
f3ZLjCkkj2cwtZ1VkKgwEQFjxpv5Sg5l//JsMoEAkkQ+ZncU6RwwcCWlvLlf
EWI9SEg7an3M2SS+f5yqlzqQI/K/jAbq9jVtWi4C9G8kUdpM7Zs8lWaRP5RO
DbhLeixisncb5B8893zcbbYajb50zas127q1BG9WbqCxgCvZX/tH79Qhh5SH
mJIsdgTOePljQ2/AK0FUs7j/uxbGaweq1p7cbnYZTAVvmevJ+Keu1bzQrslw
KzVwqdF1kVVuEmtoyfkeRdKlgtIFCTuB/BjTAEzr419tpSdvB047uy7SwezH
FZgNAEzK3yYEX80uIKgvf9BEdrQ/30pt2e1vthtBdwzV0EZ2fnAC77i1MB0r
DMAScFGyWpon+P1oCONAPa1YtYf0LFV6NyCu11IXB6jepTxnxSygVqFTpEZu
1Dxwxeu1x4AATH9uZ3PpQNqJPj3pJsKh0zPT7gE8Q++XMRU5v7ElIiTn3+Lo
QMpr8YKx6xZ0QghxhaCmmpNp34QGZuH1FrjcJgJ+QZ45ZFV7JLh1bX9ltIkE
qwnF0NmD1yhkRdjFsm5ih1weNjwWdG6oTDQSgQWv98Z2Kj9hvQ6J2uCiQl6+
iEBI6zbxbdGaEoVGO6KvgWRRuhX6Fa+2PJ7zLZx7Pa1gD6Qo4D0mhCUpzJ5Z
wxGcnHp+aQT6V1Cilgu6L/ZqqNSJU8PVIT3HLfd4vqYJg0URHEw24BzF+mwB
6Urrg42bq/V0hH7xqCvAMXeJLt4t0u0hNXDpiSTqjQoLCzFOMKqhdgvpcb0U
lHLdnHP0/WTGscc28yyNuNCBweDNJyuOVt8Ssok7yt3CMsyugOeBCI0fvV5T
Gec3MGhNVKsxQFEZvKDW+FfqIIrlT1NPVHghwAAhKCX7b8JEhgrXikV4FKqW
J4HK2ca/EQyn5h6XYD6iPOleANYmA7b8zgT/o5gmqSlJpk3wPlVLCoTdgroR
cJtcvYcnvXuiea/93d095DZV9uFCBOc89+2zuJfjeK8/1eVd5NYCtN8DgpdL
J9QO4ca1EIV394YvfGY6skqiBTVNK3rbmzLs7hpsoI4GDJ/De3Qu438Bv5/Z
4tfSdzV0QrmVGlh7NziWDZ85Uv+3L2rRvJC8ZXFE0Sn6yEaUHjMRTpt2dPYj
u6Up0zetMLQ/qbt6mNKyho1Yr2WL4uX3GDS3G3xeHMvtoSfTsohzIk7zVcqo
YSqluWVoOz6KORp/ferVXZSi23ZqyoQ9UScUS1uIkICyHpMDuJ1IxEP8NYM7
vzVUTc1l+54A27lbY2jj8QPqtKkSu5kaybmoycvtD37M81palGNU8N7XX35D
IdrDKEEEPTSUvUuOfxQdgBd5auj3CgvMEqTITCPTzYQmse23+FaRqtYpH0nm
AXXNk3m4xFYiBcXBHLaWvih2HLT9sBz7zt9rWI21ARvJusM7GMKhsNBYn8Ck
rCGwHeRGjuPzlN/Vq0jlj/fo4w96jRTmRRck9ZkNhMQ1Q77jwbkX9FdeCET4
wY9Ee3T4iSTHl/F1yJ24WUrHY5PxAcT1XK17iBcfXZFmQh1FDV3JxpwGXhQ2
itcpSGxKnWos4Zn0p3K7gMDNcKaaO+sydmhw5pAlOOw63ODzOOFnkVqONuOf
Kzbqj/b0eUzQtq0/xPTzpSR0s8QQGXlBz1yxo38K4TSPROLQCzhUvAoEL6xC
xCJzCAYO0XmlH4GUwwJsse6yfm90vweuRo5wEbEhHSp8IGtWG33S2BlGqj+T
TwsKg+J7AWJjf8Y5vly93b0H6nWDfWxy2F6EIzdbdw2jdmEHE1UUenA1d4dU
SB5BhT7sP0fWndCGBNPkr4Ud8yp4A4bQf1K1rYdEuAFMInO6/l7HTAqfX93T
VNri1032ceEeJtVnx045GkOdeC62kAQxP4ubDQgJ/GEhdz1L+oKf+unNDuLa
tw3GGkho8M6t75rZ+Fo4mU51OKyr2Uj/7Xp1caRlDdZOyww7MC1NVVwvFxf+
v7oqrXe9vILFIKfnMitSvCJJbQ4CZT907LuQaz/pgpi//t6r8/HWbZh43lg1
YvfTGE1oLC9g9Cg0YQmIFrxIwG5jfObWvnIp04DUcIdx/txNqWl0LN0lTd6P
DKFOdKsBkzJY5vN/zXpQBl0fhQaW8pj6dYsKGo+ubexCwDrYmJAHUkDLQpzS
svxgTwQSHa93zmvg4kuKcdhTYQ/z6ndSWtOr+Yi7LOkmFD02ZYjMx/swmA23
nE5ntNjQSMQCeuneJidmHk5nKG3RTKGDywWJmU+W7oC2vWh9Mvuhqm5trepS
RkzrWb/wRCmITAg0jhvJRK0Rox7lgr+XyAqyi6WMNyZyHqSbuJDqIum9B05H
1IXvXRATAcwcrKd5v+vs4X7cIWR2bm6nrjvj5YXXN1RMIygmGQankHA6Bec2
ovgIxsQ14CUGhZlM+fqYthu9GscX/mcYgOKPxW8w7QtenCisX91DQAwKAzns
FC9qpEU5rOcUPkTzME4UkkoR94E9D3xgmvSTyDKvFH47CW3XYTaX02BkZcK3
Fleh0GJsx7JTHY2wcL4TMc5sQ7KLAbeoOIVsLmhMwhbeGC+U2LSn0JHCARbo
c00nlWxTsVjync/UTPpl488B01KpJZaCxR/MyKgxTDqrgT+Lk8XZfoOIZ62q
k8D/ZUlR/Jhmyd/0NGCt6F9+JcpKw0gGzvPCgfBlZW+DHHQL2DKeKoP3T7M8
29eq6xlb7rG9oFW6dIcHFUFPHQFWIbwlRGkzwYXW9Qq4TLX67d9lMdTdgEXg
1qa9A8r7NX1A2IR9xy37j/WB7zlu/szg1KwLEYGvY6SFJOX9LWef/9KJyjJM
bjROmFfd2aXhraz20JYmPL/Nh+8VcR0DQkg/HRB4KlL8to611o/fkaMCBrm2
qcO/TnhebMfMmtRxrGax6369N+6qmJBQowM4L/lVPL4K4veKKnZIDGyngLnf
LY3LiT/Llp029dc+tqUlMR9kZE42OUyzuoJ5aUGzjvW8DzX4RPiXNl0aVGQZ
OrFWtI45vmetvWJWFeNr2XHcg48tWJdBzGnJaMy5DCZK6WaCxr+RN/xkrXWt
mRmTiRhO+7ZGoqhJJ53mUXSbQTUBlmbCMyOO9csd09yLMUjGDGxbc9aopcHp
lPhEyvtZhcJ72G/7DGAart8ybvfr9d/nhgMgWNAyXJIFPEXfj3uYUN25Mw6o
G2Ck1IdCMRmEujcT4bwe5oXfGi1WXREXH2nAYtE0Opf4VGokmkfV9J72jbdj
3mPETOu72kQIoJ+pLPauSqWvoBIxjpXwUX/mYCzN1/Sx2MOdEwbcrMcb6M0X
tSgo4KflDxF6DQhVSzy4vjPSRoRpxHI2pX3aK8aTBpQpz4qJ+58O0P8Ff5hu
oVYF3AT+5PHYcC/Z7OL/76tExj+RX+drOff6kq3KiiFhaFJuYdIrcz3oFU+9
fKTEx2vp2NvHdFblS3lPAh7+FhPvJ76Lr3NKsQBmU5OAn5x6K3EhVvNmMTV2
H7IvrULHm8vA5KqLh1f6ZjCpxsY98JaW4NsGLrBIGDaxAwhxvwTa7vkeOZnE
uw77dpPCjfxt8+lXk1I6lxRp00l8/VptaIhk73q6PYx0XhMbkOUkqZ5/nWPG
FXjsEQyDEYre4lSNYMBaJOgbtA/O3b2GoGdcr1Sf89gKEYZxPMn+No2da6L/
yrQKz14NrNUPjcGhjewCEf+TDFFyf/zY8aqr1422wlYKX/yRcPl9RVgTGnDp
UeisvICHivxPI/wwGMeZHURWoPGj95d8s8exTSwSKAwcKp45LbYbYntssAw2
aLlLVsdf4eripdLNKhREW8VF9I51nD9flKTDzEPrrwg5hHwE4J5CtlkF2ylD
9WSWiru4klKg0IXZ3vNdIFe9X7b4Esl4hpvIuBkv9cjDb/EDm/WxVUlc4aEw
ifqU1Gdn8aCNXVg/jfCOCT3NC1Adm+BEFovZvt2a6GAmkUG/MF5w6eO3LFH7
7c2afthorV3BjpyWHkvy56OXnj2V9EXLnOFxb9CxZtQhzZ73FQ2YvGYQaB55
/0XGSaelUD/2jMNxcXV6Xmuba2ROFBKwxkmlEoQVncRByo4gpJ2lpwXkMSxO
rxXXsNUbYqgs4aWcQSddqmYYO0cqkOdPSrC1Jx0gXL9YrCM4+GxVwhPT+fyR
c9z6liEyqwF1aJ2fmDl5N0InPuq0+UEpi/ht36XHJYY9TK+Hqm8u8PmIG58N
kMDObzmeWRwqO82Xc5vZeUtvncZ1EMLwYfWIY8sjsE4+poYDKW7jwdnTM6lM
vCGkUtYfpsU/dZw/P/krY7sdLM5TplcK9vWXJjB2SiGMa2XUr4XdVsQUbslS
hZOwPKm5nDRsHVc0y5LC7GuLUGIwM68hsHjSFDV5pBnb5FmHjFrbuIqKMBrs
SVTt1QKeO3G6ExCLLFmdncp0tLdi+YQCWjSNfUKfSC0L4GPqfPOeC4t/2zxE
6ZP0kpPVQElPOCtULYNefoxAIaCsYqT8HWmCvYIzIjbXww6XEoOjmVc41pjk
G3JkVldEo6EKU5FLhqgymi7LJ8q1LQVh2piq2jHPYSijwH2vZkyYde15YCXL
+bVa+MSH2DNalaFDlFvc3tQoZj81Id+w28gl+Q7aj8V5VvuUs2WG4zY3F4Y2
eSPn58nZWeFMxvyOuEjR9Bp9T3DSS6f9KddmudzaosYZLuGPqm6vZmfXmWBL
EHtRZ9HOPILwhylzC+zUA84ybGVESwafP+y7uwk1T2NnWbWxUyDw1GmG8iBV
FZT/2DoFSm4JqBXHA4ZWfN7v5r4TCZVgxxrHoyN8mGjxq6fhleu/Whr+WKc8
cd1NfijYNFG4KTFYJBKvH10bnig0fuSDuJbpIQ8fR6xb8mf+/0qhVZhbAw8A
0VXWUbFq1VFwRlBetJrR1pPoPGkAv35AnHlWaKzZg8CPBLoypnPcW7eWR0j6
4m2+vhBGpQAwIKkfRhd7NawnrhdqiNzOi6V/txwniEO2f1OZQRdMNm1Gf908
mpOJtbxMsUGP1+TX8QoBREA+LAkHdndaAetN8UYMoXVobkG1BKHgHtfOYdbP
fcnbBsPWqhROkD/RVdgNuFkDZYsCtSpCSy9Ab07KH4Td0vpC7JlGRuMV50ll
16zSLOCZ0q+dWZWhSjlcLaNQ6YciiwY75x60WAsMeJmZ4ppBgsLzlKid9Gye
WAP9OxQXZFcTvXwtoSV6GSJQ5YjvyD1hX0S3nE+tXLHz2eQyZwEosGYrfUZt
VYajnNi2hpCvdfL4vVAmz7IlpkTj3e2IF9GGAUkAZkmpkAOPm4TCGo4G40iX
mcXlK+KxmCqAcrhk5yRuE/9mLXahv0S8/sBEJDtLJuHPqXD4tjUYgpR6XnKU
pLzC0Ar5Ht0Jvg2C34k/qHEamLHiYzGpFVQC42EwUSwId10BMzjFgXnXdLYS
uqXXzuE5NBxTkba9UIpW+FXfxdi6VHm14nhnhiLnxzCmEAawgjxv0Qkx3qql
TgKNyu8qeqFowNosdQa8xuRvFBu8dI8dmKJ/S2C8uuzrvrS3zPWcbyJr0vFB
9LJaBwWCgg9k0mB0q9Cv9G5WqGEGJ22Xgw5PE7lo/pFJpMDavePGMYeRmUNU
+7CzSI3U+y64jXc6fM0xG+22LsVLpxSIt/NaP50BLSbLlelvgC7pJXylw/+X
EgSxGwq0InhLo+eSmuiZMdA8Mq8/rL3rmheVpRu74UTjoD3lo/CUuJqjKcAR
X6nuLuOyjFRYJRzRjv29WEt2YOyP8XcsRI4eSzqp1U4PfVztSpunzjCNGpss
rg5880HgxokVb7W+c6XgrrcN4vGC2JiYsAIrJLhagL5CTeOJfRWDZpdo+rK+
GCvU8U+C0DW16gZU9pi+ziCoiq7Od+6Quaa5PS1JQ+RVOzQZR5nXnDJVKvzD
bnuLDdLrjV/ys4OV4YRmhbi9uV0RNk3jaP58FXsr4s9P1E/77ZsUl7CvKKG0
01SfZdJMk0ck4IGjcwAiL2J58mj1TQDVwCRqOtDqw+UJatXZlh4W/5Y85DMc
l0bsAx0xwz5i8YzGimK6T5BIz0JRmLCxAnHrSunQDL/P7QkjGmABAvHUzvZH
dfjI1WaivFi3S2Ce3DSZwK/0BN5fccS8AnJhkbLQLXtnDd0nKCg/ong//WUH
6zj40EsYDU4jUw8ZZm1czP2GmoDoeV0IM5ax4iCV0GYH6uAOuYlpqU7vZbVK
NSwcb6kMC37HRE+YUwvmgsOKhfDVSfz5fBOaaZOXcG8KSGpPqbTdDMPgZWC3
6Cit3y7J+PGxwazQNPxClQcGmx3MN8Kgdp23MaBS6wBgpOcfZCB4UMgL31I5
zP49lu59cjlrphHw2IOly9W+7Qspt06mfdN3HjmY76+oBtLkPssDxqbSQIZ5
Spc/m8ossqzF2soBT3f1ItJJfeV2GYzT1uWeApKY82oIVXAYuJiJC37wT/Js
G66BjSq1+3NSwvKQxU7Zu/Wj4ya2w76FaGlo5dKWyHDCtc0HDgoByhEzpqUU
+chFcLekvS5QZJBevm1wVGfgIOJ9so1Zwt+ML6sPqoe2CTmPkkgdl1CRAEMi
rfJr8Gnc9G8ChTfVGExI4cd+rPoISpOokirxQtGBnBHyJ789vRIs16Mcxo3a
gIhze3RgBTSGeIMvlXaXnMWGIb2tb0R95ArWyfjSfRidN89RuqETxR4m8rSh
Mp5MYeJsKKTm21IYlikY3AEjnRyPOMgqYBc1r1bOH52HxXsMdbrHv9worelh
tursLbtT5FI4JbxqSg/leCGUywbjyUN2Y5unxa4dodGOzvn0mgQ7BCxLFoq3
DVieuVXkvmYjgcJt2ug29XPQJrRy66z/mC9FDYaV/waB89li+axX1vdKkp5M
iSnowJaalc5yX9SJXQHir7uofZiRdHrxoUyjVb8Ph8OEpeC9OqcZwiDkBHBB
BQ2W9wbu5fpgtpoY1OMLD8zIWuwEF9HthszbtnXW6Ie5pdsBQrddw2OG71RW
st0VJaRajGUG2+LZkC5D7sAhQ0ZdTrsUknyZHpflA2Sd0FnfTly5A4ryvplH
fBaPuesQh+b4CYFiqFPmWxvOkDPPIYaYwxa7HXc82PDIw7w/hCPoyP1Yjelp
5x3y6oZvdjJDmVqxB0V6iWrukmpWsTTt9v0t7YJAcSzUInQeRlzm1Bpqd4WX
vf+deNf+tRyuraiTwY9hg9QJ7mtCiEaC/mypz+8Tv7fOuURmF/o3alM2Uvss
nBB4eUejj+sOD/wB3sz5s2DdM4ZMGsIOjQFn2se23WfzVtXuI4YD2NKGor43
iI/MTFzGT6k49NsB9vE0N8hVMlvXYrQSSgBXYNi+jAqajI7RaQvwtOsDZRQ1
DUHYKqTKTRbq62I2Ov3J+knGrQ5pSZxwrtKgEqqvHL20tZLYYjkn4Awznn0R
XQ6cygm+81ylleyqT8uSmXAkjXIM05QAKeJv51+22W+7u7ls4Pr31I904xn/
0e/WkpphK3YjAsJKPyRquxx6XESGlVnMyeS3S9Y1Kuy3Ziw4eyoVG6NofsmB
ReQVgbPUKS/1fUj3MaNQVlJHIBkGU4Fo8mWOlJks/RoTWe3aHyYJt+hp70Ws
DVIUxHazcMukKG3wMmJ9n4joZ25vKf36uNzn/Jps851Xja1LYqmqPkR22+Pp
3muSlTK1iKxGVZiRmAO05MJsk+mRBHr40tnCKWA4fts3rla9Bu2Un5YSmypM
YR8N6FR6kT/ikKvrdeFSAPW5/VTCKQR/XV1fx+mPu5p9xIamnZnDSXVFx+f2
jS4lZ8HXHAiQQCmgZ+0UwH2GSTiu62uWVAdI4lrmdppJYoumAjUAWol+vZMi
vzsdj76BsD5r4CXRVTmaqG9Av5UUG+MtNVgcJZgh1r5XR3Y1PacuA3cHgkSD
v9u5ja8lKpidyUbuWjCvmc+nE/poSPntb6p2yFVtvaeoF33n9ZXsXTy9d5/W
DBAQ+0PxVujXDACs8UXUinJAqBNo+E9zUUzWjzRobXkd5TSlyD2DOuQLhwpA
SEEEy5WXH8rx1TV/PtCzppqBDNMuSbssWDLbcSqylxs7tVEjjJTMa5yLNmBv
lml1RQaEw+Yla0bqfNnnAA51ArwlQGtcwSPVlhuJwO58MIf53w/w8k5u2oBK
p5gsDMoHeMGVgjkFLpe+lI75sY9oHdKo9PuKzivZoKi3koXCFwqR8BeZNNSL
YE94jPtHsVaQQ0/jWOaU7GpEJZYETpGf40oMwe4QiQFcLgHLpryk1uweREdQ
r5G43zOQPqtieilk5e7ujiGAXwDfJGI5rPCeWotxBF4Dc7BKcN4rd2bRRCA5
Ozdg75f1VEO8JW20AByygKbwzAt+6m2mIM+x5NQ0Z3wdHzTGZnMfQe96VBQS
TN4qzqwddutImThctghDQTFcoKpUnaBDcSQuX6qQiSdmUFp5TBF0NXuJXU7J
WB7Otm7MMD5mH8Q+9/M1r2fT9CxG/vJ1tyW7xOJg2JUiQh4a5pjfsPir1RY7
CQW0wdU4PLwj0aev1VYI7nN6Vkd5XOivcldx5Qdr3xDXtSsO1iGpDVdGr/We
40gCpX3mBdSvZ9ycA1D180L0el/JvHbY1sMuMA1fDmzbmU1YsKxKEL+x+u/H
0FV+LAOOvN5jRW1nPpuMAEZq4MFy0hkPhOrfE4cjhUARzY4UnAWoXxSWm/bh
mZYmPOR3ORfKIV4bFW3cMsyPkSLbmnPGXiDB/HrmLnIEdDoiki9pBuA4A/Uo
GA5cBuEDdxdZHh6Hf+CYzMzxj+/SjwDLQLD+PhGsl3xBx9F/T4QxoG5/c1gS
zeZ9/CZEvsiu311xS6SHgt/R1WuKB1xjtKc8fPYihfHtDBbd0TtBs1O+anhi
dtJ56XsBLs7GuxYaA7zV98isUHy52hs7klH6FQo9ATHAc10Y3ceYopkKQaZK
3TUMklRoD7THRKGa/ImChdCMWBVO5xYviXMZkoV6R9rre6hDpLFYc52ffHTX
mAzr9apag8rZFP+EOOItWgxFn8PgU7htIjC/4jCcCEFnV6IEnX+AR+rcIm9z
Vi69O8gPTDYVzpkET58IsEoZlGHHmwoQA7CmDPFIVanv63JWGB9pqlsTDsW9
315UgouNAZVZwCZf/Uad3ZxphQccfOxRh1rUBhxEpqmBYrcJObjZRXWHT/HN
9NJn7EbnamBxSqOmKiarzLWH/eb5Lkb/SIumNXTTBK7ygwDcW6YAzeFOsigi
qgF8V4GDLqeSqr6vtTlqUSkP4g8TkHj98FNgISMHjNdk+ACS0OzZH41s6wTA
OugeinmZ+xranxYVbGBmNvAr8OqgYNF5K4pX0jgVT306ijljV9K6Bg+58CuI
tpZAFUMKZ9ey/AbRGO8JaQRatJ6Sk6RriDLUyY7AL+pUasDsD1ojj1wWEjd8
OlbMNicHqgbqyzfkWMlkrtljtoqs0p0pqiDGYK5oSdnybwkVqLp2MVxehClE
b8qcYum90OSC/O9EI3T90Y/aUl1KTmcVyRoS2T5DsdNgPGq8WICRM+tlXUnQ
N3beS+dNfozX6sK2Uv6T4OynTKy3LndQAQKbWEoLe6jM17B5cR/f6chj3oW3
55vphLD4eT7bt6TCT9KbRrTlqVOnnM3U0BOblWCz8N+3pTBgbqoFzS9Ul215
2pDdIAy+BJ3u70APKFgOmSYeY61gyY5CoPCHVVO4JdpJv+NULapBYOeohV1v
lBo9wRYmTbZeG1cNHKkEaTM5nrIXp5IB3wVh4XF3skLsadkoCSnyBVOSP30F
bMGqJTi9pd3RCgiAQjhqkGAnBgyfaMTmCSjSPW1DHrVOaouhb4I95QW1/n6R
+sDByaybzd+AdKVqRrPGKHsubO1hgtXXJuRbu3mUE7JAFhDKuwPDlT7Vxlhi
46XjGM/E1iCXnFlDY2UZwQWwrs+TzybA1m6ZaFF1UmafBshARQnKxyhpXCBv
07ar6mdAM94v6MLN7RQcIMM+7abREbDuxnY0DR7M3j+3bEOBiJBG6iYVLNcJ
ECYzxJwO3o6YlE72pIBrTMC1Y+/TbOU6e5LjLokUSDomXUsDvwoVProvJFAW
ohBUspmKG1dLCa8GwiAUXsHj2niuZaPLlcJWrGznCfLw42S7bfPsDCAn4zQo
nG8LCAGx4xUe3MLeOwShgNCJRgg0rDG+EuRv3nw1eplhzg2pSRSM+YxmDrUm
3Xe/uk++F9+BLP0pvifnLZXbPS5tDxvh47fwGANfpiFWH58YXHvKfA5zjdKi
+S2z5Mu3viBj3+ttfVvMp8IT43lss44M9fJsviIt+CWK8SmgTofODK3iaG8v
YcOtfIcJPG3xwQkMgNv7+cMVOftBlsYPnBhZpPZS5WY/Ri2R3DrxWmhaOIEX
dJs9VbLM17qOns31i82IfYeZNqOf5i43MmgtA6d35M0BcclAPgp7PUIs5Bgy
7H/wDRz9jorNaQ6op8pKTkKa22hmqauGIqVuv6qfsB1aWQrIkJM5+TjQmxbB
+1TmEOX0VyKNSgcLbZnD72xyn0CFrMmfMoTkduIxBKykSsar25oZeT1ek25M
l2JfJD7XNrD1r9mMFWj6RE5iNn1659v3tIYEDbuW6w7mCHO3PBdMcUK8gE8J
DkHVcV8t7WeNwcsmy9BxUCGYbmTOLNavmI4fYiaNy1m7IO99JYLHTmwDxQ4g
OqKlq5UvkuVjDXo3w5lQ3KMxixTnpJO1LbHhlWVlggPBJ5Hcoi/F3mTBlvZu
AgfYpjPmygvVPB7RYeIDGi1uQurXpfJZIPmz20tpcIL8W4qszwEffhUDvdvo
t4K57Q2dnR5HaZdY5Uuwkky4xfgspAmVIfoDHOKJVeVLLo2NrN695LP2QpbJ
ayQbX/HHr2xI6rQFloeG2asc0ooZ7A30ivjJtXy5u+ErA/O15C/8WJwqwhGP
ybudpDYxhVthpHuRO7v6iyVDP2FqyYFdmslJxOVcRfgQOj9snBjU88jCDgYO
Xxin2IltJJRUpb84HdQy9L+xqIrc4kUBx+kMkco/IL1esfA4Yf2kI7ETv+K5
qoLxkm6zNZtms8lxPsQIAnbpXbO0FepXYw2sjN8mcroKCOg82cKLggJs7kwO
kCbTd2Hp6MNyyHdGgG8f8aY/b/DQ9o74sqWNbjmG18Wt5V1x46HcylIgAKTJ
7Hcm3A7RlIYTm6OFXJAclFtMM5ryUMszFgzdwLhWt+hO3zLHaSlIounLwQ1j
3Xsx4fKXmj5dsbr9dTvJ7dlOUjQsgj/PyEffKD9WMN55EDhSS2M3+yf/1Lqv
Y6pTAQwIuZvVvKZP5N9PXy2Ny+XDlgMc6AXJ/uQMtR9A/gqcPdzLg03ypDfG
Hy50xEQ6o8TKD9plHet/yEwOZXXN9pu+Ff4DHkndyGXRBoGlBMZtjMnd1RYB
UPiYNEUn5JSwhpq+CglAF87O1Sv4m9rX/pauMuj0eBA5AJ1xEP+Fda0Df+YR
3jA64FuKcD2fl0cA/k7G7KT1Ft2rCCKnG/LhBYkEg2f+NSyADmLbpts0ULfU
uz0G+k2Uvx1efIbFH4iaW21SuGQ9/XUuwWc8gWkX7Dv3WFscXD6GsxBDYOaC
eiqgjfdlNm22tiC28xjNDm9YCisvFEfuwhgTDB+zyMPcXjhbNMuUxwDLcXsM
WDPAuZO8p8mnOG4mVcZB4BM2CXjSjmdUBgJnUtzAiHzeg3qJyM1Sq7IIHEa0
2mPj7bafyx2Xssda+0kVh5DFROGME/klLfYgTNp8rivx1kc/DoYh4GRYfH4U
+nEjDKEmDj30yffkV+hGx5Tl8FO0k+D6Gyx1qKPovVxRLqaRcyy88JGwgPTV
q3qQmMOUxf/GMLaRTqfs59diJUWSrGLq3oH9AeYQ3517c7TQOPqn1B4cY5e7
gwXYscuUNCP0kZqGCZ+LufjKmx2eLj6/WTHY7eCFIS97NrtGOpze5NBkdrAG
FF44N/5jQsTrMT/Em8+UvpHu5d7XsjTLrCQTVXBVs3yFb1q8mE4LQ5fekZsF
BsrSL/Qjz2e5+qmjlUtnQ3emQyZoa5CkkFHeQyoKZOqSGCNUGpCgb1fNluEN
veJZH4yvTrk/JAdjoM2xuSW0DRSZsZ0iZ0nb6BlOkLaqBJ5JIvSQbLDQ33Sq
/k67Gc9MO0zuZxwV0VcGD6o7f2U4VHVlVtxVbALTSpkODaRUUUdWfoZXkLW4
NPzc3p3UfKwzRWo+/JF2ow6Nt0v83q0xLIs4mOxFcGLavrEN/36ECBwhPGV4
3mSUoyTmXcFAdbDOMjdg/weMvvoKJlKFIJmZ8kI9rXndMYFK3uLnyOdm/UnA
JLyfii3QRavyUX90m8DI8D3DKLh/peP3Dhss/V/fDSAEkj1JEgXKDYMfKcvn
jyLKSfKdV4g2h55RIA7AFRf8ItbzAx7o5CAZ3gHBcdBsd4hLa/3m1AoUmeRy
qtKYXQjVQFnR8J8hnb4P3N8MEcQjvTcP5DxcHH4Ba+XikOHxEkmFbJDp2pOC
uBYbjff1JKURB8bocXWdPN9CyqW3HjBWuYStIjDN+BrP4nnaFWS1875pRm4b
xugiHxyjJTcbtxbjyEoGDIQtMqgPIlPB37q7tiz/yRuWVPb8rXOEpY4tkXdd
U/fY6Uz2uB0Gyocbi+85S7PZNuz3asjSwB9s3zqJCsVaeabIJx3xbJAHWq96
zFggSGdI2h9rVqjFd3A0GpmU9OoDotcJdw17xnx7wr2zUAVhptXshpPnz2Iz
PZxn8maOoDGBcjO6e6rLeH9ADrFxDf/zTrUwGFKUSh486wN2g0LMtut6dGgB
b4jdRDLD4/i4ys4k19WBylyHsqBMUeEwZpdB0tVKiE1KjZ3cYMPVn811vjMB
S8Je2mk7KMO9/QRWTofVOc5AI5y0WOwu9SfO43FobQUTIsNp43m8+8bC46q3
bLepGfw5ttuk8rQcNdlz27Jg/R0VVbk/18etgzR7SyQIPaV6djSqR1H6yHAe
0kBGVZTSMW54PRdOkBnN9GxwaW2/BV1FappsdlQkKeBq56wSklsk6Tzxo++9
BzDv7rJwaJ1YZsK4Frd2jl6yaW2BXynhUn0PRd4fBBipFtyIBcG1/34cT3BX
LyF9T1wsRIWcgnANdQGDcrFEzWNusDjlo+hBJM5bGWdLjQeYgOWMSYYYR4Mz
2kLkx7ONg2x96G1f4lrJ+dNGtbmNcqyLWNyi6KHfqZ1dOJau+RM+PkfnMUC1
2LnTreSb+57kjo+B9oNw23FKMKKL1RjVcflye57tICyxNb7pFrf3h7dvEooa
UAB8CIjoTgDZ1XzGbtDMEucsUf7k3cs57i9BWptrMedCMcPL3mLXNqk4/qM1
t7qIrcafcU1fqTGtLMxmLL8O594zW6/1XXKk7l+/GNyv6tU8Qn5xC+pcBC/4
avqhEgPUbRFpu+a/KSpqLNyoGpsYo5AJORXJjpjr53utb2gZaIU6gX+WhduS
zFOWBiqs5cMj8VRgKZv0mYJ3gqr6rv7vL9MLF9Ur1v8RfBXGg1R1C0aW4evF
7Eia9HAaUTREdrG2QuDvED2NzXbIeP6SGXMb9lRwr1BmOLNU7tBvBAVdovsK
GNrOiknZ4A90ZZQ96TVbZD17rHIDnt/KFizILOGKNy3pzUR3fds3r4Q9UAGa
VJtzUEVdpPDem5Evyx2R6meRy4wtjZsrdoLA52APCFha8wvarvuaF6aqNKkW
j967TtuUwy6rI+7TwOCnYCX5CXyGzwZXXusHgRpI2vIPTDrz38dkEHxy6Nui
4fFXvDy/2HQ9oI3OEIgjD6z7X0nULprk/ITH5Jd29Fosr+tjjsRxS2Nia+NG
CopSUqx/BY+WX+BClTIzB0h1Q0Zo9EB0LwTZjPEshUaFRhRPg+NhkGx0m1Zu
LbfBWfBd4ZQjACge03WDv0HmZRX8mQ2fxxYWAVoW7xqLcjaShRBx4joSLeFd
QCEilnsha++2TuxF7lYnM6ED2X5lFPBK5wDqG5a86jexR3AzY1E/fCK9F/Wr
T15XgfKcqcpbrHIaO9+7hN6aZdTtlf6qGUQj3GiTtM4iIv+idhcSX6xFj1Kk
rmSQb0Jh1TrcRpw+xGJzfW1zAwnzCB/0w95NPFft3fs2UoN/3UZ1K05ubb5T
7Uk9ruABCinVCN4bxxq5ilyPMOeqd8lMekKVN6AHFAryfczdk8yMfghaYe6K
nfFdEdZz0ecaLFzq68QuibBQqZudfG7AXEYShGNAHtBswVyir7bgJhkWeatz
uYe+DXp63JxGfCB+5JOOMhJO/yhBAkGdQHxz1FtX8g4snKSzwq6yV7Rk2Iw2
RPyh7A3SI5OrlkkNImy+mYX3aWCyem6w6u3VmwqCRFvI/HAgQmjWQLhZdA1B
ttXLaLQ8k+eTbwiafC9q41CezQ4toOJZa7OnSylC5GZWdU4t/KJU+JWn4LOa
t8qK51ygFv+ZwbOeMgHQTKrQc2HmCaLvygW11uuUH/8qMTs/tJuh1jjCV9S2
WmKFc3pFcKRi8czEBlsq1XOCyj/KWASG1X8AUJuIIw3yYKbjarhnd0goF3Nz
n0uPHqF1m3S3exz0ws9siCCimIzWfifZBsFGHtijFPP2zn2fd1KJPOLfyydh
L2XXKvgHIExDXDT8HEFvmoaAaSWff/RBLlKmYguh/jqFymqRJRzIUpGilHFS
2ttpW9smPcUuDxgX8c11zORpUXYeG0w1zJurQZLRkT+3RosbX29vz5ep67es
rYUq2cWQjHQoq2ODCtHw7qwCKTOJVYWpnrKLdGr3G7/YKAo2AKpJbZRVCYj9
+rd4hbvZ2ik1yxVC5ic/i6/bh0H/+VO+n1Taw9ryh/1XJAPvVzeG2f1T79z7
xQcvtxKsJ2v7el3vvVBSZzjQL5E4sHnqhXsNcmX0aZV0GOb8kLeUdqgcUG30
+mraeb8YYGZudrBluuqPRhnlVgaHwr5mhxHgmAeVxn6VNrG5hROfmuFsErr+
lRVXUqPWM7gvYGVnawaM3HlsoAWoZHbfUW1cnpn2itdbaUzbuh/qeCI9hQ04
rV3ssGKdVgeO7Lhw8kyXAvKiVyqgrN+rOoLwlxVlrJdk1dTmoaM+EZlLG0MY
+D7zeceDNRBQ/zImcNQ5vqzpJWEminFEJxMcXhoVgf3eFVJQFHx+9XzMgBHN
7YlKuRljOmeSISQnzXRu3G95Ok2xaUWnMqaCa2MAUlL+ZdywYVh8POX89gb1
OIvNiNIuwAMRsvB36sew2KQ9i1pz/Xedc6ftaTpKRhA6dOqyXtkx1RF31lH0
OOCw8E7eb2U43aptxRtIuYxQMDYly5ehWb1uc0n1YKH5+GUAlr2Y07svw5/x
jJ0rcQ8ceVjLECjm3xlETkj2nI+7PeGJRG/dmY2Ac0DzuJjHYk7mjuID7ygq
Lb5/ItqTdDKQr30vT+IgAl81Pg2HgGQpOmuJ1j9m8BbMcefLLXV6lcDL0h2B
JtDAX3fS7FvG5I84iBotZwKM6eLm1/P06IgKloQ/rRy/tJJaPbMAMOAQYdpc
pE7f/IsLXrTVtMyKxfPMBxfNdBPqoVWP1XVzhBBsHBvwKhpkT+9p9UJKFlUo
dpYoYfvSD7vj76VW54gL5UoJwQUznxqOX8EhpJ9BMgGWWod2WXi6RR+FYFgs
3mM18MB8RL0QMYgzrqNk/xxA5n6uA2hw3DmAWW7fBI6hfbvMpO4S+mu4cnlc
3BqopjtN003rwH+Nc1zeIP1ZCSXPp2o1sMW7Hfshr9QPIarwVMCJeDkeXcuL
bjn5K979FNbyrRhvAt4eoBu69cOBvnI8DBwOebzy9nR/fkEB6lh6HjKmf0Jh
aFc6DVmYeLtfAwKy3pdTKf+h9eQnFO6VFEXjoEh2uQ9398SNlDBBZ/45mZAB
U2GiWJ058qOjN6UthHjOYxc+dFlgLafSMJR8lEbsKPEHm3Px90bKJphHXIvN
JUQI/p32bqoaWmBTCiB1D0TXfG0LPJdunoDEBQCV03h0cQyHn9au8SGEN6qE
mS+W1TygyX/thQfZEvSBk3cfOgIeYEqgwWfe/2ZZoLJXbrG1reRFeBr4aGU4
9BplSRZDG2OJUffq690b6Is5UOg/R2fUIUtdH3Q/jzfJ0p5J08o524RvY1Ii
oNg9lTTUfd7bksz7Ldf/DHQ+ktzt488UOmtSNWOr8JF30zlB7SM55/CY/kGF
L+Po9eJlycF2vlUbDjfqGTm87xCgSzQlSdD0ig7Ii4vy8YiC8t79bVLWdHZ8
+TUVg6fSVVkEIAMQlfu7zMqF6JeJEu4eAaaAQN5eRbcXDJD8nalxdssqfgLi
JEoWMUvY2oOi0b2bzK72qJ3uIkPliSutKDTSMCqbJn00TBPYDWGRrAA+cQCZ
RG6jLIATOx4/NbfZPjw5Ck0CWS/AEJ4VnpkAPLIivwQa9CnTltp2d71ycV67
hAfiknMhJt56qQZUd7QTgqxjEHDE9wTS8L2Uxw5bcAQsrRunbRqdr1XmSBtY
ERvBjBqgrPzRrT9hUBXQYZgKG72JpFUXh+2FD8zyt0g9obNVBc+8txkPyi5J
Q4Vn6JmoItu3Sbn+kL9v4BW5XwWdwcFu+xh9jKWattx0bvoy2gRQWHEP3t/9
85msXGoWEBdZ/oqinAp4NZOKLveewH7HAfR9V+UmoUGurvBpDvGmVWNswT1c
DDufRLcP4UtG+B2PF01EsaXA593HhPi8b4S7kv0tltlX2VThu2ggsvx4YTRg
o3r4MeHVaMlrcSw5Sq3nQ/HmDlulnkmBHo/93cf6irJKiyQ4INipX0siUySt
37EbqTbFZHmr0b9OGzIJGDrq7BFCn6UmIS8rQjwZxhDLAh5/W4cf5I5BlYA/
kITa5aXPa7MDmKUD5PV/NnN5JLBMgQqffoC+9kxk9YIYIOeBYHc9uHgs+yTl
3Y5MqVPyUd7bUCi6KGHOWGbO1agsyje77AK7V36PbWLlspXfCV86F+Zcc5Bq
wZG9A2G71QeuqomIizw3B+40SszGF54F9cpsUeQ4m8f1xcZmGCV2I9QUHizG
qxpTWIuPKEG3qb+YWettLT4nSRfUy2b5LZOHCv0ofnHiY9UOJtYufpDccIwy
t/1jGLkQR4Md6hPZHsyCWwhPlLIBxdWip7TyzvmEQE61DCyGnIRFrJezxdOG
suQ7wBLcsWh3Qy2nOV6O8a9xwvODpkWLjzEWzjFFaHTDAZbDPQ9vbnRKcwcR
psiYggnoN1g/YWwPwt84Kd2gHgslMOWdY1/EgN+2VSA40ttApsd1IBlehvd7
ZvxOtAIxrpt0IUzuyT27U9wO2bZfKOeG4g7MhOolEf7pL4K7K/k08j9BMN7S
n8Vd76KkEJ6Z2wcUVZYzKdZxTqYjulmSxdu5y8SGCO9+dABTDkAYuBSzJPaV
zD54I00gT0H+Pu4iAPKmDZ1zsii9suH7mhxFiIaI8dKlAuxG/fKhXSbNcQxB
4slsEfnKskjEqJdUZgtey1mUZlDVdZU3XwBQG4Z3fuQLLCcEIg1faHvEN4HS
GQqZqpP54WApErV9mIh/0G9la8KyQL9QLAnRm4HF7RuDVV/Se8kN3BboHVpi
UsuZbcnYi0ZW5FO0pBBiY/7686PfTibhgx8R7pD5xXRyOZDM1tm6+MtJnAav
9QkHaxXGX7850YNE/trz7ZYWfaICSt1niL1Gt0GwA6/06R9yzdkp2fXNlP81
n5p+oh1WPyVie/CX+9HA0R64eFX94NiKVUrZn2P7DQUIIKC1ezNhA/YRixlB
htam+kHgd2wzQvY6F1mGklIlpLYz3xhsNvmzEgzuIseOfJ21Zab4H5eZzqqD
EzCaE3KDGadzecsH5LKxKIeq+XIKEYvTDTE4+4CTX6TVcDZT0VpIwrDwvq4o
wBog7CNbji3ISaSmipiInER4zs9Q5NAeOHwraYXxzG2sybOgUFTH01Jp7vxR
HEtuNJFo6bbjoDLp8csiPR9nh3se/ZQTZd3oHcxecBOFzE/tBGjiVwRLRWOr
M/xTXCYKGrKyBXf8iOFoxrJ5HwkThCXiKZc3i5jsv77GmqWK4lZIzkMk4nL+
m0i4oWYENd6/AmyVLijIqn4450F+XMa/zRByzrSZtD/RNsdsiHLZoEHkc/lg
Fs2TqAMejmhJalw2TWoLzqgXjXZtiQzN90p7kcvU1ZDbbQaZee+Ap9F7GJ5x
RCvOyad6TG9e/zWi1byrAjGEsi6BCAYR1/HzVipkpRUXHqHltG0yVKV/hfXt
lJdv2kBAdcCqBsSn8U83jBLYv1R0K67YeLDm3sx72ZYiwNJEnfZkAB5XWdFn
vRYO7ABzHRDHMQeKtT3NBWVQAFN1juGeZXiyN7oSzEcel2/ESFfwEMKFR6Hi
tOXhzTSSMps6vM7eGkB+GWR30CSSHifk7PtJN6/1Aohbhky5IC/v5epFHLcg
Ev1xt3n625JgZ9WQXz3NAGWKrvLY74POxMYOLRRhY6ZvqH/pVy2qcW4YGQL0
J/BW1QaE4R9nQvkQ59vEQ/CTvP5MrwSA9NUA0CZb5hnTXOxX9B1j+88k+7h5
IrccOjLpmAOqTqYR2L0JwlNa7h10mxhcueyiCZD0cpy55Tuk03q3Etbc26Mj
fkzmS28NSMNBmYg62DpsEoTUkiWyGVly5tnApXccYQPy1YQl1QiMeJ3A6mVG
ZsvOHZkrXvUnYFQovTOmQ3bz62GiMW8z0YyQ+G4a/YavKDNKnG+3ho8gEVzD
wVF4cBP/L7bcvWVSOVge0/beMGZzoQPorIoTMKZyjvrvopgbFiPXK7MCGt7o
ImVGf9ONzbE9xllfre3IWlgiFR8c0x4kv5Ht+esmv2/3Jgp0SnVBIuARcTUR
DcBb2nlnLlIVXQPHr7Xo+iRI2pWLUM+eePG6kdfE/3NvOrpLMUyzFBf5FJiu
RSqe7a/J1v2FNrH3pw2BE/40PTz5BdPUOT3Y0061EQ2io/1CUhfpjVnuniW9
wyyoQL3sdsD3GSHhaUZ6C7vgmLykXo88mWNNuTsgehgbx8Z9Upw/NhR/dy7K
F2A/viQsEyfVgTuAwVtq1umERPdwdIEipBiDBV9wpuBKKGDHqVwG33Xw8PU8
CNKZLn27kZbft/xE6i2ga8t0vT6ra+xbSwiPDmiB5pqZ4drrthaKJo42bq4x
ZcrnjhDWb8KmpjxwZNDLEkgk62/F6d6X8IGoC5mpKTE4ZfCf62ydeTjdF5f7
aRoSulR0ZrLqWN4J9SlKQP6XaLTbdH8CP13P5s15NxlGZWiuaZPkRpp7bWjU
GvtO8MRSD3vzcfB3oJZjqQ+ohqj3hzv++R2USRHqsX+wKO6BljNdEfagAN5f
OgyxJA/NNhrKucg1cRO5GxUNRGJRv9smhTKebw9Wz4S/s0F/jto/sML+It0l
aexU/0rp/r7IflBb/yQt7n9xbRIH8l5ksHgSU5EoKrBAtdxPrTBOZIIJ9q6J
5FZ2PWIe/sJ5Q2QXYr+wu6RgXJmiLaJ9/nzOo4N1p77csSs5fHYOcxZ7R3CF
bK2si/1O5NVzO+LqnPHAdxBoRc7zusuLbNeyW8rV6cTq097r43VPxXXvKfG0
EBeTjXWN5i3JsY0yXTaaNXr+HdYRYW+XRgWByaxFeY/lHrcuLkgyfOQYhEBB
k/42hL+PNcwrj6kyfrsAnPdkYN/zdoE1Mn5ecCxL6fflhTHCR+BRh8PfDex6
zwbzXcHbnhJh8FlIj/QivSQHzcdvCrYcDRaLhU6PWXblNap/YXqxHaa+6IXB
tsQH8EeIXtLr1jgV9tLtKCIe+AzsVqVhtAAHP3WYTdWisfp5jPteBsl80CJQ
mlXcecB1TyfwmqySEXxP7tmGgRHoHmv36CzADBK+CFoHDJMNOEU7+Yxyl4Nc
FZSBN8ZwWz1lnhw2DOP8arHfFXMFwkxOaaJFq9a0Dhf3WwjeXo0ghq8rWrhY
RdBEEal5ztojYdjBtuwCFwDFy8wX47MonciLoYOwQiL4hC5yLNr92+YDnG29
9MeHu/YBlpXRPwXKhp/lO7V24mEEGQzvjFLCYAObxIUm6QkL2waOMKsQkUSk
3vC2GzUDOB+I688A638dX4I47TIhjpYXkscdvlMCFz7Q/CMbBNqVlQETDFo/
jZVbmrS0duV30v/C+zpo1aG1/nuDVYY7xvXtChhSqGJi7rqtZ3Ak7y4VYV55
k2pOXJnExQzDQAjajAEa7aDZigfEPdDO+zskPnm4Jm+xHe1/tsE6SZqIbC48
o8AD9JPmeazSLr//LBPcAAoxWKkqArsw5GqiMgljMXzLOTEbRVrvExO/xsHp
hLSS62u2EqB3DTqFxBSI1xp2Qc0I/XHHjzU+niOG5e4n7Hc2OwtiMoTMW/JC
L4CZ/zI+DvTUV2jrgmjCQEziBNVKtc07+vcifribTBQuY/pxd0Q6EuLUubrc
fNJqbiMsq+ebHUO/HPYqzNSW7Q3UeKwiSJUNjCx1+I7VytJEO6FoYEP3Kk7H
MM+MxilxighNMabcoHiWVcFzQPYsrxZW1a9rFSOs9OAmL5WqW+szPCFpHklW
qvTR2TsBhUBm9Xw2FiJUOwe8y1IF/2oFyDnJPlRC5mVibC3Eiwc+QgfzYmbA
r6ULokT8vs44Qpye/kg0tkFks83BxpNprgyVHz2idjJ3lUuO7bJA/1+cLtEe
8P+uW/43ZE1wrHpLmMkW6fdxtB2jnZ5lXHNMkMtAu5mZBQY4BrI8iOGvLYtV
gd45BkS7Gejw+Nch8x9ikmeT6f72lzHVMoObaiGAGvdTF4UxFlQ+1JHPnLab
X0+dRiCvfEsQIuHZ1N75lFEo72yWJCjMilp2r8tpasx90lJ0LWlszR7nikDz
hZaDQuMovlrKUShX4UDdHmuAoaxMiyr/0EtMXC07Rlravmlgkk8Z7uFC0PRu
u83cno/45krAnkLAMiIMEpSQ0PlJ6SCmOacIt2jWev1cOKNxOimv0XQ3UhdD
VR8n3U/PN8EudM3mNJe9DXjQ32T52Ekyo7T7i3laMddulV92s5utuAeJos4C
rCLT6zdEyh9Z6WVRZt2AaibTDF6VclCC9uDkosAIkbfuV2AHucynYKvxpZ5i
bkfz8EM3KbNGqbHf689TfUyNm+n8MwHtxEeKu6nrw9DUFFHv9Re4mgbFKTGF
aBqZD8YZAxunMNJzahjtL1X1XVymjDAMBxe3KjKbjSWc9kmj4UHJL6LmTlR3
jQLBPCB/3uZDc3ZFMs+l3F/rXmjrkmdQ+Cm1hLhy/4L73GfjH/hvOGRCxN4t
kCRWr8SiOuLYOmsb91tuEq6TkwLdUMT/HfXziXdqXORAoGastDiv0IMIPXo9
NRzwyD7VSnLw3SJ+6v0mehk6nO2T4Tqhe0TTpkR///l2FydUlocLOEQhLYTY
/WvItwaN6sdEQWjpQKBk375yOZW8V0vXlDpdSTg/gW/Ec9uBwt33Cz57aLRB
wgdJBvQXyDCn8/lc3e47QAHDNgEmhkv4InftyLs6cQtM7sN7qefAhZgLyJH5
TkcPrTBkYNOxu1fwH9u+t6UletCZYj4vtVW80oVQG252DK65hDML5TGD3UV4
p7mktYErPYXcZ2H7aXxBppI28G32fV/zG+6vP2APvxSp3dr0995zX6hrv8u9
Iov3p872qdG73OFrjzWA1BkwY8Nrm+BlXFE1lrXoNG/oIzmp9p4sMBtNG4gO
RFHahMFKikQi8aZR8W/wLa9cWpnRxSicbDkJOqFBV/OdsGYy85KbE8J8hHJH
ZK9vtOk7j/bmwm4b1V+YSdgrWCfUsszkqZ7qxuHsW5kQBdGOposAxnMM/9hM
6et/jJ5SokyjL+dxqozw4JyfkuWnHuY+O/kYFpmwAErrRYZki3569qCe38K5
AiM9CP5/b51Ek8bqKjJC2Ql9lahOp9mYBjMUJ6Ra8l1PBt3ER/yMtDLEdpg+
qj0NQhltWaREtOyaf/WUgkJ1uvpZ/ObA+1jQoQ6XHgXfL82YQFVdGgs6oXm6
vse6i5f13OXWB1RqlrrsCa8tbW/YZZFHEmAPDtnl8J0U+ftxobXyMJGN6/bd
X/MAbHbIYMSXhgTonwWFPHD9kMECyMLMT79AR9RCrazHIVWk57GyLHg+EAzp
tU13b8QRmpxhQmsa4bku96WL97Nx9ehF6LgWfbYPrbkwmqU3YfZPzXUfmEyU
v3+CzifvgMLph5PfzsDvXDMTqPb7YgxOumkGiIuGmxVvsoK7SY77o+n5c4cW
X42oKhkXZAT31IKvVD7prh5QKvZdZZ6bSdPss57nhfPt7IWO/JpvEzOPH28S
kuh/l7+57GSCYG+khMCCvMstu7XX2ELwLeKWAmBe484J5YonlR7CSju5bLk4
IHOOVniLY777QjkoX47PZfh+nwytN7jL1rWrBkzeQUdznjFSJX2+JuzKF431
XTTppe3nGoVsVV74Y4TgfkgYeZZHS2+QZHO92sBoe9Q+pXg1As6CHf62H5N/
rMM4A2WpVtHTRWFzwKUPk4MiWv2WQO3Jzs8iCoIq/bMr8l695/8BDyGrZ2rB
fI0iaKXVA4bPrpSxasP5XyMJqm47qAyhtvKC8+H2DjZgVJ/xToREY8zP88Eh
WsOKtPwZ3Pt99sI0RZLqd80UeegT804X61YuFtImQXtdhT8RHMrRLP88VKc2
Gz157lfSkZS6PDb9KHSydi95QljJKoPr3yL9kVhYb6rEMoC0lzUELmo14JNe
u/QfXTqo5U+c6wFTdG4wUUeqw7NMXczqsnyWctqgdHeDvZ7LijcQcOW+XEMX
nxouavZ0TIchmM/IvjGHXDo4tRpIZ8SttuZMpdXe2qhV5IkqR9b+dAxNlw+b
DV3DaMXXhTOp8RgLH6DVpVBt44GYhlqgVUoripuIQ3hDv2BBYcNUtbP4ns4+
UhoeQKup28liAw4IQZgmTNKc/BD2kuSN50OK/7yZuT8DBjunHjPf0FyJnqUE
cxpDNiI9WJRTAt3fhM72Ct15/e31ZfCiFdIiz7KR0LYbI1sbYWFvYzzcLNWG
Qt+FjyrMSiwgHd3D4IXObpv/ZzZ/jHNT4+ZshvE2TX28oOhn9Gu2wBv0S0rg
mOeYvHyC8G81Lb5Hn/T/LOAxP0zjTT5oCoXNRhH753ugNi0EHq7HGSI4530l
1XjDaNll5ZYTw5YciqVj/sP99sBiPmQYyVRk2lE522WslSmfpA2zZV/NUSJe
0tEgJBibBqfKOGds5iRcUGqWugvpCnoO/zprJtGqyIB+exStnSn/5wSez+JE
SJLKy4eTgXEBQRwxdH6iHRv/V4LbQJJLw501BqhA61hH97ThdKXDpZltTN6S
tKK3pHuasXq5kDiq6sZ4eEmIkVRbTkEuf9NIABdv7nuZ8R2UZ0nS1FlTOsHZ
bZrSJhiCeu5bPV85S6dTYh2NmOWkbn3vSv3EXqlBsoCxsqxvpmFnt6/ymKmc
U3QPHD3SUZt4y+7ZurjcGgzYHPUnoGjyVMPA18gsJL4am2RJqMeiuhg8cyz6
cs7o1yshX52JEZpDNdu/AIgZbIEG5FEHcrDGvY8/rRBjeHcl62OIWFX6UG/Q
dNbUXed9riLjzFVLy2jABac4p0Dq32MqvsRmLM35iEfEGOTWbXWlZDdJSoGc
OoJjzM2zxZXYXBcYdNdwFmuxIhwTlZZyeN9jDfefIcxdoK6Z1mQIVvsAx5V3
APQSM3WH/DbV6m1BCU07tu5R8v0TrRmb1ykwaUIleeqnuKwYOAC/NXnJI+/0
K95mzsLjCAiDLN2TuVE9Ny4Re91cPMdqeSw4EpLCPA//VZM4ne9WWPPYBuiQ
rqvGd8WNsbnrBayPqZN/cZ06AghlPGquPXcbH/CY09S9Q33Acx7ZbSEA0wdK
CrjXPU7y24mluzbMfTOUzpfeXbBsbXeoeyMdIltVeeLuIcVYP5CYNTgkahqz
TVVlBeKq8XYn/gGVqAwS5Gcg8r7MsHWxr56aBmpeMJj33bvJ1dalzql/1rbI
I8BvehJdVoVdt4wWkn3eLQW0RCczKABayq4fllpgyvgk/aDsmhl7Cf/TslyP
RDLS8bX48gx+J1Hn38BUcYFjP+hjtx4q/LZSyoubJluH51G24bwG233cQsTs
VAG4pwOuV3NCQwtMFPZEp3spHcUV7fglH4aiuhqpPtDAS+bcJ+SySx+lJFOj
0rXrxh4PJuZ+m7ZTUs2WkFXArUhtrd3Pt3GJYwoVcoBbIQEXepRKIE6NvUpu
VExkJy2oElBp/ah3Iq7FyBMlRB0UKD12h2G2wQxy3p50v8WtYEWD20FICk5M
Z+GAfvXOCPyP+NCfQMh9UhrcylMkrHduTS6S6fJ8KjcBCi7vDJh9tG//wYyp
tVLzK3z20TLiVjqjWnkm09NlLWrPkG0QQr+yRxDekoy16YQfu0LkhU+7oFdJ
A0xCswVFDTOKZC9CgHZf5jJIkH7GhWpvDnJx/Ce+v2rhfpM7oNB3BVp3Sern
1be32DJqZnVndXjbG+vpfPh91Mm3WrhRyov2x29bvu5ivGRvAxrElfPBiq/u
qkiw+vm7po4aWEWD9T1Atti+7g/3sAc7SLF1W73MzPzwQ5Eivv9S6OqR3axt
BKkc0n7zX9eoaXaRCWO0VPx3dBnJCecuMx8Mv6+4ieVHu+SY3zo+O+7echCw
B9hBiSMmOL4mi3HZDYnIOVc9xAucItc0p3HpY5ze5Qwj3Y8SmuQOIjb9TyRi
FVvML8OsGfD+JoYcwgaxHHO0QISMOzYkS9AV/j8Qye4xvXsrCKfDLlI36O5Q
8+r/huIRR36yaaD7KpETCrJh9ZA2wytQsOVOX3BpeyR5sCJT+8t8MpHXQ2J/
4bGTK2uQ84XQupzwo9vkEsXohVBWcTBfkLFg2jbl94jOQdIrraWgvlsroic9
hPgSNurujQEWyv1jTLF35uEGqt8VPVylvEdTqB8RTXRE2QZuY9iX5gQKsvVt
SuE4z2/AbhT784lPh+ntu/AWznIzW++2CM0PiQI0u0CIEllKRu21mfiJcAM/
7WX+VmVqa11GRdK0GaQhZVsIoTr2I+amAUtRSA1ioFi9pbdmJ1kbPJy6p+gn
qS1yC1K1BGTUqdFxUP7xCMStBj4K7vOlh/eldCMDDbjo3chD5ZNhdvvbIzm3
uikEyLgyD56Hn4l2GmeYhWfGKqIyK/rknBKrhRhGGUhzO9LTJSAvvfD6Td9i
KfEFY/llxmagtlIW88MfBefqEWGQ07Mhr8KjzDWM4Iw/eKnX0+qW52HVQUF/
UYPLYnauuSIfMPNYiEX4zE18wqAA0TX7OY2wpZ04x7QwapbeTECTd1H3Xpp8
K8Ehk7MelqfaJyYZ+JxMaRUpn0KLXyZXp017e94SzemJhmYQCS3Q/20iDC3E
2Q3KnfOOQbTM6LB4XK+GB3WR9HxMx7c0oH0q9V4fRAFwLHOXwqac/fyJpCQh
iLYD7EQo30iQxhxoCYElvrBcicQ+M6yH4WTynSbisFsm3udZTXV4WhfFJEk6
FEDe62DoB0Hv7p1rka9UUM7KdX85n695WukGvF6zVZH7j9Oro6u78g+omGVD
vYradxuzaNu1YpPPs1739KFnxB3zW2P64A5RMcVp3HjSjcqTzuCUtbkMpQNt
9lpZfEi0AEodtYV42omHjl4vDFP4Ka0IYYBOLfEjmoUiq7MnKMscJ2hk0Hh8
7+Yg223IzwX+/1RKOxYqr65Ntf0v8y7nxoONsuzBL475dE+afkBCM7ZuVW4U
0tG+dsWmRnzOnvENDpIA9c6pUhe8kRYA4K2heu9I3xH3RPYE6lZi9jyo8N/s
fEG/vx2iLpPjPO89/IBk08mwl0+JgprgskbZgMLL1Hq02M9pYWgxyVkQ0LkZ
a/jx/coXosN3YyUQkFL4nPRw1CxLw8TxS54t2acTyTkFFeSMvWsmAcqNmn0g
dpOyP2GLbehjVdlr1SjKmUkReOneVETx5LpN0+2b7B8mcdcqAGSVBVnWMV8x
0RjK6xmAauY/B9sBf/wrcQOFnoqQILtEsvqBJUnadECU+Q4TU97CFl3i5lJy
vHSs32K0m1+fPyIKdOSmhtRFarJsp/zUZ+gkfHjz48HeY0NEwhb4f/HH3cFe
mdhxD7corAoAACsZbII65LWna7kP76rh3/aa87HwWW2Tjrw4eGZgLOygJgwW
vcxtqbhyv9lt1nSo7rUFZt33D9tjMRR2xMJVEkSArhexfVNoS5+aY0s446pw
E2TMCzfwjLk5rqpt7JWIxw4HWgWoEvVQPRUATvn8jX10MG7eUf4B6V7BoiFX
plmDWNmGw0aY6mALR4q/GCcg7Bu5EEztfQUkjoq9OoA16fZf4DY3O4EBK/nT
YMYWokjUw+oTD97nRiW6pefGnhnlalFUCJ9Wcs2ETeBhT6i9fEbZcXGL5cFk
2EXksghyPySI5BYNUkB8rDIQZjE2weJAmY1/Hols4dDHM9yRQqomS6h5PzTW
P5FgJX8K5rJrGIpB/KTvTc8B+RhDqi+ltaWPX5XaMoSmgk5Tf60HTnSoSnoB
W9KS8GQ1Iz57ewZQpwSmt5jGhAMTxHfOoJ62YeOuExOH63Mse3WbOkuxJhv+
WyK+1U+fZEitOmY49vZn272xzWgiPD8enFn/mZcV3OuAlS4DolJaGfguAr0I
OWgc2yMB9TLCb3S1XOr8uvcLOt66xrPjEaQN+jLxwvlvUB/6ilCtIb+WGImV
J/lP1RCwxcFNV/WsRdeMI+59dTsZtbwvE1Iy6XXwdFmcpia2j+cV9IwCqdoK
vyYUEyQmNLwVum3ouep3AkDYwX/FT6iIRwYwt8VrkNQlSCHzuHsUkpDQCXOy
VaXBmW6kmM8mHxmfiCP3Tt56cyiz/xHvt0pjGkZwcwQuFEXMG+WjYypnEC6k
5+pEsIdLfoKcTkMHSgH+eGJkd5qHGVr7bkZqtOcgS1G4vIPVb8KvdnLRQbE8
XEHznVBJijqtVFq/YKkMTZnHFkYl00ExEJgEQyeU4Q6dbaW20nlpXbVsa2q2
eq7h6KsV4i/WZNiN9BdBEICHRMmcXesFkos0hE0KV1oDzu5Wv348e/DhDBWI
Mgkd1LSu23YPEwArHx+uF/bFXlnmppkMeBZic8FCp4LLNCiSSQ7amlkbf/Gl
xFysE5zWiyTNO6NgBGnzSYXG5MkmzFQIVHnepl69QnoeCqigDNzpOoaTTz3g
B2QtbJl1N5/8IX2JEykmBB5vXxzEaYGWPBKAMtwmFq3CKTZOK7nhqof4TDLE
hQruqWwsqviN6//e9b93XoBq+cftrKE3w46/3tBxKYrp56cdQQabGzllmYpv
shTekF1IGcnNt4t/zbxCBrNecJ5oYrWUntWagm8wh4n3GjKlwI6t8lsaz0la
Bi7qdx/P5c9djIu9Nh97n6snKri3LZ+yH7vogdnbWQuZSctWtHLT5lm6GY3U
h/hhauJ/PEPaAtNBoCkWZHk4riJ0CtAocupyRpIzhh1FhOrkxHbJOW8sGtAB
vibSPiNGxu6Jnd47utppFMJbe4x/Y7u5BrY5hF0yzTQhpr6Yc/YfA97IIvzm
8T6kDXOK7Tt7O1PZYRFXVSEOkpiXTd1Odwm8mVHfU8spahrifW9KKJ37b79J
q3jy0Ep48lHMteh7emJ1sMcpwbG5LIeeslSruxHYFKeUAMP2mezoQVUXOFiS
E7W/aUqi2MFOI+XiHstRE07TTZJghQg7K8WZrBeOgvnxDvWFHmfbFiypmYSZ
Z5P58QFyojDhkURnrfrxTsXuoqCWMoKnxxFUfJt3YWBIw9l5pZ+13Pd1Da2j
ajbl6JEa4/qikuz5IoU7PUm+2tWQw0iDHet+QDctXQZev4Ah2YivzD3VwPYf
E3Kk97fzumsJtpl4eOWos4/9I12TW4H/OAeyRQK0cTyQGY4eDS2ZLIlt6ojQ
aLAnRN4OGjmsO2W10a6XkZ5yd/chC6GMwjLl8Tz1pNbIYhDCOclwYj99Nvrt
9KYcCkFNCS6GBdgqZgypGYK51SzNpigFtjsAyTwjasy7zFw8C90jPSz4hvHB
b9pf4f9LvDhFxAIOdfhUJiEYSsMmq0u+YIdZzbsflYO8cRKCi6oFpKyYce9e
ora6YIWA4OnMRvrqn6OO2SExCnWDr15pHT2z0imaXXXS0AvU23GnW21HoqAr
lrIC+x196xUr9d79wcL/oqZkDJMxL30hqemCXlOWODCNP0KFDYHm0dXNjxa3
t2FwaCgyqL8zcOTs1ZUJVVI12VJpnd/ePqmpmeXDPbezTQl9h/M02OvYcbyl
nxNyjIHPf/wzSyTSF4xz5g7c1+ubP/PdpzlISlKsrpPN16icZG6rdJ0a2PlZ
l8RWWqv2pizEVAFygv2MR1ADRYQV8bTPFvxEgtO807dFbqK04GFOTsiTp6NA
5R2dSQHMc1kNZgt4iG8MROhR3SBvH0XEsvFA6BEOx54CuhtHjZiw1kWc4UA7
2/0S1hv+8OK+ad4bxeBAsqNPMzJ2RqTleRIKySWx8K9pSVLSWc5r2/7lgppE
NFlPbVqh3qlT9JfTQh1uXdDvBufmnQjhrZzUkfg2y7ZOkd71t/VkAhW/xdSJ
qBAcuXNED5mZBVg5zM70opcdQN7Ze9L/ukwyrrGibjWlji2AnwcoPBFWK9gf
SbWryBphTUQB/CLQitmpL9VAPgxjEW0PmNlkpDx8M1s4kHhb4Rnwm9UBfbre
JQVLxsNzC6w9LLXE9xhyAJmpR9nDP9oBNSEQNrZDhRWtT4WQDwx8IdeSYhuS
fP0pmjmzfIbcdVDvlVRPnzHcjzuM5tR2n9Y8+dnyCfDB66RA+HdCpQ+bqhSL
DyJ+2tFmIjz+LRt3CPykt5hbYQci+kAPeC7m5eXGOoSQ9V50KwCECo4IocKb
gnglngdiMECFbhcHIYC18yG2MahjUQup43VnFJ3CFlyqgsmx5NV5uwxV+P9P
r7iRzGBn6wjt+tppneMQgxLusiAacVAWdpP8FE9ywe/VKroB7StwmEh9LLgs
JgcGN7WsGOmFK2OKYojkDpq3J1bGhXNRVr3x7+3kaj3PJ+gk+fVPxlN25tEH
f33/xYF0ISshdBsyauT6AJdKt5IYH6KT12gWDR9vNYLBwguVcfheCquJdQhC
Eojdontuhq1GYVfGsuqEDb5IfWdAgMjei5spfSfZTW7dNimjOSUSiB74o3yA
7GEll/DjF4PLo5ihK4dtd/A40rU3uuNBGqorjYZxrYjBg4OPe9Lj2mF10eck
BTLXsNHFCn1XAjEH9TwHza2WPk2LVfhRFmin0pMUHbxLq7BqsrTChHJTr8z9
RNe/OeeapFdG6NxzQS7McLaE1nxJFzwSL4edMmT9lowC95BdF/6LXeChnHd+
g1UEYBFd+DtWhAEwfhzNa7lnKSoE/RrUdQZ6bHpCMunpkEOAOHOH7k4bhvvH
lEpBqRdOTN4upWxJAzRwdhXaPgapi66PVOQbpMzEd30ufMUI1Q4FkzRcYRea
L4vhk5ZBfM+8gEHmyXNVMo46tXVuToToMHN80Zq0cjUgQ3z9xUDY8ScyZ7vg
XCGGsqeRT11tMhUlJRjRxL63OKEnUh6qRdZtkCr6sm5FRIGXrNdUU1c0YI2X
ZiqSiWMO9yogMCEPQUB9AGCGTrZhn43T3Gd7G2FPovrMAmcVs81BgS4z8Gsj
xoxkld4UswiLMlsJRvvg80Hmqw+ARx9U4JWMeKwPIdMxtqLKvLCPTw+qgE/S
0A5vaFfREEchDG5KWkPeDt2VYguQuIGOJl17rkyM+CL1MiAx1UgQlY/iHASR
rKPRM54blqfiuQU7ImGq8cdvlSHLfAskdh5Kjcqw1Iz4yyCWHXs1quOSrQlG
cOFbIA4hStbZ0EBtq1i49NRJcBfftTq9nwF089gKlED6DLHQiRJZVMaNzUcu
o1ePmFPYTqV7UPRNqO2Zrsvb+QsNdftQq4royHXnsA7d3qcPlmqLekHvjHVQ
fXDGjzgHfNac03Z23PvCULloFf+YLYBIMrpRim/8JjihLaSG4J3h4/STJKOD
iV5tBdtxr01lsLhPiX8wihlZP8QWVuyBWvgWVZIHVVGwpMnxq4izdMJsFKM/
+gxbx04bAI4+nylEcJ9px1p8wGHJw29JLjtqrO0r0GFZg4bPHc6vtwuXihzA
nJZfy8Uewb8+/pB6HXMps4LKgJ/ygbA+F/FXL66qVI+j9wmIk3EI9j1IiZTa
g3wV038r4qIOMR4aDb9TJ3T65bCnKGg1CcIK0Nce1KLCGnbJmmtEpQErN3oa
696gCSh7Evwt4QThouypPsSEcziNVPNat+VZa3I1cYNp8/qZdAFzK0kSeoOI
RdJPd9VZCFlRrlMZukJgc+aBXJpXXiMPZch33fYkoHa03hrnG/nQH0ovTrHz
GPm8QArnrShqX6f1Xie7phNoNJJLe+JIqVqQPMSoU2RWGXRdaPdhNIJX0us2
n8+6U5lxYH0Lfdfxyex/YetWu9ARjzlhYSfrvmY1Ew9hL3vVJJmCB2yHLdBD
AUwl6JEoTqHyauaqBFtuIZjSLp8tUfCMq7XPfcRk7ZvIgAA2wF58SDIPOl2I
eGjuUFD98aqIxuSD61r8gIu86EFfmDgPPuFWca2D6qQ7leT6HuXZKuvdTZXx
KYhHm14DLWW6iQuJGKtJWBYEG5MCeG6U1wqEvseF8iDvewKct/JlvBb8F7UQ
2C4z5/L+CEhQpyaCMHMUzk3LeHdPOJG/RbDYf0kK/gmmonYAb5HWcXHPT5HR
3Kwk/NECifDs9fCT+L6VhM+ul9gAVYtNby0COXi15q63DTJA0WJC99fK8Mlg
S+eZ8qHSmJIMtVVTEZr05jtZZK9Fegt8SnK0UezUJTo28RznPgfYzXPTG8rn
VB5HqMiCuMIZp+p/DX3r03mk8q6qbcDtiFVTFG/US04+ADyFHrGeCpwwBtB0
pnxEKb8w+gcS21k9Q+WS+nq82xUkItcImk2M+l5FM/VNrqskVnsDx6xW054Q
6YTVk9zWvQbjmpD6gGWcLLfrt/Ucibf8vGe7v47KLaTp/fRLs0vftuer/tV/
5viZUkUH8cD8f4LwOpJZ4z4FH/DyewVwdKBLSU/U4o8X/EGJEiFTIXHZrDSt
pLJEZWQ5SS27JebguDEk18efb/sv6Y0xMY6zbhH86dy8/xU7G8j6rmdDlAfe
3p6ggWJlLH3gaYU1MgrPusNCL8cbFkGys3agoXw0XDzTqav5Bnuj/U65aviR
/32t0ro8kpetDFSTal/AtRZ9juknI6mZUGxhflHMqBWmaX8wu80ShOgSz3wY
ug8E/shJMrRTmmYSFICBIuUDl8NwVTPQT8AnGFtjjjZKKSI89mF65RdHrSmI
25qk25TWe11ud0c/fDgb48KkdENI27ZNW+iVXmB6WLuK3paYMCx6lD3gCdjU
5dgmBA5OSNYQ9Z/WSetcxcM6J5vodCt/boXsaB+KrWHDwhDbfKWyC7gLcUYl
L/HUrQAPEn8TpICcdOUjBLRUrKtxANIbBkEsM2Oej3AMJov/XWFGUZOmFo3l
xKPuD8WACIsOANPfrefCCxP25AtcoY2/AhRQqF/TnjKXIaTLdOkNR1+OBZuV
u+58KvpChOtSyOPyPpNH4L6z5ssTfhvhvlsd7D7bSTTwBNHBsQmxIer0hpan
r9hmY+z22gl1Hw2BT8oemP7eNFvb2llOk0J9b44h3Jy0WMOR2HuYDgY7LEwd
jw0flY2IQk2o6fS5X3N1yZHC4bR4b8KfUl5qm4yO6lBs3wzSh+wp6j400+6P
GD+0IU3H+M5IOMqvnu1MXJcH2/kV4hpdkh71HUjRoMhnJf8uHWdkEdAUV19e
Zupim1g9H7AJDlwf5f59eOFiJTJnVsZYB/VW25GoRoZ7aP+VwNmv2Ml8gUpG
ad6eFVwx3t5PqCA8bpIomzSfFWxkvooGjK3dwBzb9jxo0Q2xUb5sDPw80epb
RKUDMXLWmbnBJ+wjpH3MPa6IKsv2Uuwnn912jYvfV5orjbbPW+P44oTHLUwC
YbvKfZKcokx9ps6DgamBqa3B/bD2IRwjRLvNEWPIMTiClL+0WjjV043lfFLx
OFuo56wx/p2NTiD8B9UdoT/g3uMo+tvRjMmGhGTHcS6ZsClF4CmukD4hgalA
iR3CREDn1a9ViMqyGr4npcDUB7/UElMnCcU/MdL99RYpC8uhsQ9s+QjxTwej
XVn1zxNyEdm0JWwOxnPbWRoIF2Bq/+9nOPGQZJ8fhR+2iMNAf5ujuFLSK4IW
lbL9RMCEGkZ7x9ue62IMPrRK+KTcprF8Pp7aVPlcMmF5dvHA30mKpT8TGjn6
HvFzE0txgoMdBONPSN6b3rHQXZX3zqL3lRub/KrUd6ekdyCji/YJOvmnWtnn
uO1N1ZrRf/cvScqMk/AexJ4dCq4C1rTHRvqeAxaQKwKjOF0NbmRs9ZSci7g/
W6PsCDk8adEDcCH5wZUzq0lL/aJYCyQEsfQ8HY11NTy5NNgvuip9Ig0L4Jj8
Ot+Ka89uZ/nUyRN/CLboJZn7VutvtfXRPVznt+ZM5FQb0NxOpJOU6fCB5MmZ
pac6Ycimcw1Z/nPLQFAjZJc2bgaAFTDiR4dOlDjZhC/WPI2e3S0sIES1if8G
dOZ9Estx7X+W/hnzxnQh6CsRahRd08PScX5II+xtyZQiwTnAkvVrXjcpdtd1
+CvGv0Z/yIPfRxO2L++5qeJwEYvMRBaAHQY7Chgqh8tA6IuLWuUZacUp+IwI
xIoAyDCcr6PUk9Ts4v2ru4nGvtSQkBedrSjzZp+qlfC0SXo9Syp9gHyn0WOD
BdW+XvvyfWqd/GzZJBBacAFZmZ/A2RLQo4UFC8anZHdG/otBd3vonbshonAq
ol6P7FPste5BXiHYlMZ9PsuaMbnVGwIOYbEeJvJW84+35W0UBuFMf+9wq6K6
UOtTMJC/nJ1LEXdnbCgwA6zUZnyeC9o5+lfXzk/fFTbFcItZP7Nc0zY3Zmcw
af1IG56SZpGziIy8zKKGiRUFT0mIKTPbZUsovn4/89ze+8K2qk7r/RMfFVHq
ah4kDLKGxSfhzVNLBHa8/0FPUDxTPDfyyWWEaHZjCds/xsiu3aKhLQPTsiAo
scnIAQi63kps2xyUgQowuvmuVNZMe1eVxR6EbEFUAxJ6SBGkh/TOVhl6whno
uuVJFoLQHpsx+fBTfbaQTq3BlB3qohZURjkEOIOUx9Bi6zVNUCYz17ngCsHb
/09sSQRlU/Uykx2zWLMx7Bn5TyjLXjYhKV2r47IJXZPexhUDOqPTPSelFQCG
jltXphKlYVIQ2+kt7/eoN9WUfkatLlilY8JdTk6fxX067FAHQXkNkfFB5lyy
oVIdgjyjSgNZZBEV11m+lqveHBa7+Ax+4Hltk+CUU6ap2t9dDzgS7TUOraxD
3kaDWE3YurHajJDHUQEg1Xa3d366TWzQbDjpnndUN9XwDaZs75xpt9xr0Qm2
286Civ+8A4tu1IiZI20X9Xa3VwWzxK9I07PE/TTgB/XUamhWl5Ms0xeVXAZY
7hRWpIw63KHN08L4TxoXJOB8kG+m/K5kUvZfUAsiWFOMEHb705Bo3gBQnaRj
Ot39x6iOjmfxIcl/YUUpANembVrjKYLp34+vYQRmp//O1Ny3Jh/6+MbdKd9m
mT8vU6LYC0vXsQRPhfPQ1gLSsagbrbLhP6IRI05wj2m2Len8OZVJma0wpf/6
H471WnAZMfRn15scVhRV7rbsKvTb0q5zrljMRRPfmwImCW1a6JVa49+PXG7Q
oJ44soJ5PxQnnRd58sNbqATId8XDOCxdPXP+LjbayVkd0VA/SzP1pjRxAm+o
1YVGj/uuiL4AIjJR+WcpELEBf3GgfzRanohNcc1zcMYOS/g2ID7jaGSXyQNK
tQSn3mBjo9d8ofe0SbgPcq5fMOhFOgKEZBQz1m+NEbPQ8exkdlhWqrfMilV4
5d+HODV9/07r9CWj3lYcoMt0vqHMZqFDS/MYSJDI8EDG6fl5/yoB1gDE7My/
rIZ7GaSjGCifyMj1ysR0GXNDK2j2jQmkey5aYWViUiE0XHNc51zPJJ6aUU4Q
ZFyqVkbOdv/zSLBeQwS50qjnJQY4yaVUsy+pO7KA5lL9h+ye+sW542mic4cw
rdpVfPmNr8MVQB2fwzXcRTa9KKGJm4elDvfGNycoAYElk91u0m6+HLIqzT9G
YQZ4QD+m3Vue6vWdjiObBfDbd5iEjKTgvbeV/4o/TyuG6mSSSpMTTyIkxHvw
5XED2/Y6H6OOvQMJ6PoF3x9iJUFhDde9QBEFJl7flZwqOvUr2JK1h2nPiLOn
qyP/Jn4HWrz6yvQ/GHg0DROk89uiIHOICqd7NdXVNEROkQGZqPpcUGc3+/Ly
noh7iZ7LfX8p07hnjUhVJVYbEHw3xSUttlO9SJlecho6bWPH+Yz6G3sq17L6
41jCA3fFdCX5nyUUTLCQN0VhEarsFYIE+bWpl0HL62flaya51OEcjnH9SwGC
PnO/Zxii+WN9vVh1ZQA7a0CFCuqVDWBlUkTgKgdSDt2ZACqSHC99VVJBhTvG
Tj55fMlBDQ4VWgj5C+5D5KsMvnifPukr28LCHRVisJzf3m1U4XluMihgE7cW
XL+KB8DLVZA2dshn8CWq5ohd76/Ly+K35z3GHsIdWCJZ4O587VAb56F+8TwI
T4RYfifzGWiJ5pwjE5EWk4UoLRcpZYABaGJRYIx6IiE962bPTOpl0EwsLRDl
nNOX89A1N1Q9TaNR4va+F8ZmBDrOZk0lEn9aG2LzbXZuX/03Fx1n54u6m0V9
oAiu/zZ6CyETLz/CjQgqcBMauTJ0ZYhEnDWRGgO0jSH1q94qtYCuIwN2fSIa
KDO7/ooGWcTbOYr7H1ob1s5TAVfIMbBdcTyveupOx1V56c0aER0sYFoIztr8
VKfQpeRv3nxiDXtRSvjNQiyO2XRs5+UChOVebJBAv9KS0cLJnFJJbt07qyZm
gw/LQFR97bkyqiOsKSpgRJHOi8OvUbMcVQNlGi40iVRxmSNH6fv9GSV3RsGR
7jWxUKV8wV8SyucjAwVjwKO4erxMiEMk5ehxK7AM1FCDQvBK5MX1DAdDUgur
5yBul/okns+8F/xWmEIFxREcm6q2BEGbprfkgFhz53I5aerSl1sN6zwsMhG9
xAV+xGcTFIroNvvqSMUKjJFPfIJSfVGC/9etzMG6Nev65gXPSc9ldVz+2VIy
h2jZbV4zMDitIuS4n8mNgakTc242gSAgYVRs+FtfTkMN3y1oZRkr5cBMNd2m
srVxfr7fU3J6hbm2nU6T0DaA3i1PxhB1yPKY4nncmfBYy0nKz7WSKRw03FjY
hytV+Lse/IH+rXy8WC2jdKgdESSqm3Q8hk3re65zMT1rcTxPvkiqpxpoR5Hq
huwX4DHdjP23ZahO1I2kLplaxXhis0OT1DhO3lLULXEhEqvuWlN1jX8b34Ws
CJmaaRZEFV55TNDYMZP2ACYnC0a8oerAY271eETsMvHn5cXbQvlfK0ivhkMS
F7iP+x0vg3eiUxSIiIbG8JaIcPK7LK5V8pBGHt5FM9H7jaSgJMKKEs9URGnl
nGVF75Y2OoW1fnhvy7kW612q10D/611qmaB0HUL8ZgkSebZh8W8kTh30aVTx
O9eAzo3zGpc4IubNnE9QpBRsSO3PAHapzwGJOhpbyhLDV6tmrQHLgFOHH3/m
pJa70y9yDLEEjxvUZop98X+rGK7TxxEZ5Dym9DbHOXNM7vOX/c7az93JDS3j
eZ0M3CF/quREnZAzoTr9qsNaOmy5hBr4jXFPXACpCesY0heCauiLjtMOBWhw
6IjPz+S8ssO221LxclazJrdl9vvlBjwfuvCnSIcrOBJolAyQ202x6PamByHp
IzWqr0X1kjp2Y5FD4IQXUEtu0om1SbrauPan7OgX4rJ6ko2Yr1LWpGsxQGg/
TeBYgVj2OpQt+SUTrnN68Id/8S+DBemwHmatb96c9yae3P/OmcNN8g6ONCGp
IywY79WM4wGOgAz2YCtRwX6Pbw6b1XiphXutJkGDwa1A3WMVY27gIWL7ClQG
XCZ54js9G2+2Z/pmIhL3fbHsXxOiaQQqTCf4aLMdQ/MpqobHSW5qfsWGgCaW
C62C6AsJ7IIWKhwJBS/42Hip9Pd/YoYyygIH8rT/u9uiwlTf4Lsr3Z3B8IxS
7bWKOBQSPkOQHHKwFgUkLTEyzw3wyNgTYYDHqNGLs84QE7Qod9XEu0Y8QGdN
TR+4EihQ4/nK+wwx8CbBsR+aWxWJ8/4q/AiIXOUqYxFIiWqWO9N5YdAuFrCH
M6X1uV/8/Y3jZw7PiCWHituo8C+DKaPh89/2GJEqqqCkws3IciwyQGP5fUK2
gLda1BHD+ieFqBjqXws1MI8u8NCajU5jc+n85Ne9YLPidsGTBhcxQohDrHSr
qZOAzkwvpQwR5Z4YhglraiowKWLyk5a8XTJwCZCduJt3IcYTtG9FhFxizdZB
LSDI9DYkwO7nUQcjmC5OIXQ+PrOwl/yERZ2mEX1Zf4eNsVujPOivg831DHnX
b7niFOxidIghrZKXxPp9Z50+UIQqkMM/tJG0TGNgB18QfEYLbjYdUCQ6BqN1
K4Yae4uFcmcBiobGTvsbhr/3KoTRPkBH4vIQp+HVh+43yaVr1wfGrY0alotI
FfMMlTO9EysKXby/T1Ja9Y5wiBlAB8EJIFltp5UxYOFeIydPBOuGjCF+zWOw
JXiFdoRJi6cvnjXQHEl8G8zMXfSMsg0wVpVIOCY4BP/dYBf0EcWDXTzgXZp1
Weh1V+vuEE+6f8KMpZXdiNRcJaWjqvbWTPz6nuljkzgxOzzwQbdWdseId8RI
o37Fs9oMlTbci4IZPj6HrL5vqFuJ+VYrmXcgDSlDyWjri5OI0nI5AT46nb3T
y7ot7fu/L2wc+1N+krNcz82V5yAGjaX0OeeU3SxRpFUZIKcupgdDutQPZRHs
4OtfS3c2ZnquWcVlxK7SamfsSVcz+93LqTKQE2u275YajvZpJ7eeM+7RGJUK
s+qcsPU4z8QOUg+hY54OulIqkWtbHF1eHq9wElh2AsLqDoyMERRpGZFOWRHs
0wTxnl5jkBbPpvqdpFiA96KX0C2nLDB1Jg85VMLrc4up+exwAzpZUEzwiCtf
+LMl4ajf+GgnLYh6H5HUBmFVPtQAyvB8OMvESgVXCQtFLNrlDGw4nDIL5VD6
ykzQN6yUKXuqCCwg5tcRwFIYvvZVirmz5Tkz6dXE16fJcbbs3yfugBMJm0X7
IXwq18Y79H/nlIudRziaIFzEwZQtgOsFjRrcfnFwwkd/jZNWimqarQG5U6lr
ld7DyOBcdXQIzki2u0Oj7tzkYyCDMCmCK70Tj02/izaKHf72L/qUr7Y84yXh
z/Mr0FoZKZ2EXwXyDDTD3+xC10ihoVnpIC7GY2mbJgN5n6Jnkk22a/LyJWJj
iWJW++aWvLHAk3AHBAwFwlJxDWl2SUnrFYRX0rIZAKPH+qrDn+nsPcrvXBUM
dEvJISBprqDsJbrfo0r52TFKPmJyvru8XSHjiXtAbPxY/hhlvBSKX6DpPRnZ
UwW7oCW3CXZIqx/nqJ6U+oKX8k9AEtQNhgIvfUwyuohjPByDvtrHEwAI6daB
0hTwwbUnPjhkzyLl5dtabHjhIKnGI53k13Mr3wVk4q92+N9hAcXwZNaa+9Os
/3r8IY1R/rZMQBLs19m37SWZ9INX/G9e57V7vttD7WlpIBqAyojB1EXS0puN
Y6R/WuRDZNiRDiOijx5ohbSGQBvFPCvvUti0xUWqa4HQDqj+gYFO0AWNrqR/
LQ1FnZNgSV6l13cZ9vbNC6qAYpG6YwLnvoShwN53rVZHQig3/ICJn+pfG7lT
lngQlpcGiR8wirR8LZYYWuLcRyTdaI0+L/mgfAtsr6GKS/182OnIJJkBLRxV
dTeaeeTD0lqIuLQ7UKmIJAKBw25TYreiVJpsLDKnB+oO3CnGbgS4tlv+OgZ5
bLx+MsJOQ0hiaIQsDbnzkMKRH876HrjZ7QFT/kLF1jItaFn4cnkVwNcdOAgv
seAetMPs53GrFc6V/oJAa8CQ7oggrxxyRVPmTNIE4lxpC/7TrndKAd9GVXVG
OOHlPfKJiegMiBNvuiqg2KaIq4reHAlthFWZamEoqkPNOyC8BVvkp090KIEx
ZgT4ysEyiuwhbEGuOMzh8tPZT8uXrHoL3KPjWK1xZpHPwwOdSVwt2OPvnFnM
MJk2Rkh5VfxN7T+0O/PVMQoq7Az9nKoMjXrIjdcmz075FQS6RdWT9LQ1OCLO
SNR4h8qnQKhUbVMVJKdKIBlY3HZDaOy1VaAf1ezSRoSObaoCT6XJY+2/Ia0U
/u5lEUDgL1h5VzHqsX+XzgNUXwqZMBgzD/QnBfA21mc9KjG+9kjZ0YXd4OHA
RoH9u/VgfbzpI+VaZhTzrtVySJwwH7QMjxF7dB64J3RuS9KP5Q4kf1XEC+ok
9RmBxq3yFh1tr13PJlqb7fBQtlbBrvdH6CLIyz/Eeihsk3sp2KDrOC2vlTuB
atU+yB/R7tRcOzSBuWmkNyDVyeqos1rmSTtQG5CQ8lhDLrhPWsaC9fjT7pwh
u5OONzisXi8cHqLfK6wF9jGsDXL+k4bolQ6pj3KETCu6f1CMt+HaaZINSgNg
d1TbbvfOyS8v3VOZCMyHVePCm1jIqPi1S55yJPqsMDF3Sx4H9vscvVO1wm60
P3KnIQeJjcWaK9ZczaKepBLRVQLI4rnwoALiyri1qD0+XXrJSyeGQh1U4cFC
8mB+7OP+6U9FKBcldTU38ZX99CioAqD6UMVJEDuyngPtzT8Ttp91o+0/JWSv
yQieXcpkgO2Y6rog2gyyRaLob3a0wE+3cUZ6yp1tcYrHeIVVXu/8Y+h+gmNH
paneDgwf2dg70xNeWGLz+i4dDAnBtsG9RFZ/3aF+3T1uKPqAX2cf532nZkKV
EVMiZkbrm4T9dbzF2LwLlcSiS526OENrsBYCXtZ+ZhbiAeJyv4bEH0lzIS0I
PH3ChDPwHMkY5qb5I+1dH7vYUq1YGzMWgctxkYxDEaW4TTH/Whbny5abbob/
4lbW6cWtCWQPeSMLtDWlU0i2BiayVNPTfpyHcFkdpG6xs3g7Jkho8lZlNNVB
+5tUbo+tVpOz0JKuomiqTS+nUNOKXkgTTqLh7YTtDsllkmIQ2jy5Hgx6mNxq
D9dklAg1ar5vFr3rSlIwyD99Kmr1uwLk3YYZMw92RGiHVIvWz6EpOe0Vu0hW
wN8htaoTzEwD4hAPFFk3XdgTvAoNp6ZuEatJ49RzP5npVMg3zkVgVjeWQ9Nc
sPsAg7QiuxUnT8k1mx4KC6G7wFqkVmUnCjiqjxRKqeGUgyZAPgWzlE8qVz1k
qKsM9xKsh5+5dhhTT0etStFjP6Jo4WPYZl0K5wXlpZZ8t/P34FZ8IY81m+ge
3HkH1L14FhddGkP9eP6g+ODorV3yxmDkNewc9m2jLHCEQAObUu/smIH/L6UC
fySNBVXw9oTG2cRGiosljecRrwOLIQqCrtIB5KpySBqiDrC/TalIcIhKslzd
oCbFG9jYJYxYHNgaTXXF6ZMbC0064vIfRakaWv75+qV7QZQ91mALc/e8Bl5Q
6Qeb4UiRiSOtfckO6iEcm2UhGIHfY3k6sn0pMv+0MxXBqhsd0bcFoj+wlOWv
OlvwBCYWgAKKLkxbgdwcbS1A8wH+UBYS6zt9H4ZfFRuGa1OgspGrQfcBoKCc
l6T27EK6BfFabHfpqSUm5IBtYh3Hxzs90U1cdE3UCY5gVH2H1+0Sp6aflHxA
hHIp91DleRPoUrf4OP94Z4wINU1SBiybjwaBzbuFHUAvvU7x9fY6Ra7DjVKW
oCZyksykch6EbbcDFc3Xpg3lf3fYET6tOmQFCjEOCRzvwxtlyOVkzpbgUj6S
aBuOEZBkgcOPz0HPR841F6H97jR6WUPBHwyEoYngT5s/fotqjBgEXBQE7My1
R90ccQZ47WDez7j+zhMoc6J9mI2dnM9CorMDdWcfM8FkVsjZgcAcPkUeajVh
g0GAbj/lmpS+CQiPOng8AIA3hTsqB9qrhU+qzKx16EFJ3fySw//Vrg3UbBN1
cXb2XprWo2LjEK6BikFYxby4U7sxmbOz8Yj/kt0jZKHnjuLOxK8gIgs9+0Ew
5EOt7Osy9kCrsJWEDtDA01nacw+dioh0/3r2m6vt5H1XDaRROCzBU4CuBPC9
9EXINZnMdwU3H9o+/iLS7JcfaIRHqx/BEdmpoUvR2iAbTO7VLgofO5SX4ES+
RCw9eTmO/UFesgsqKdke/J87Y2D96IBKlS4bMp/xQIOWVZiZpTsj0Af8merS
YLeJ4VPYzd9tssfFd2cU312SW+y5FRRDOE6tR//wTBqJ2GBd3ogshpN8CmKL
xyAEV+EvXxLI2y8VneyFRspJ0qCl8NSIIRVVTqjg0rSb3h8TVh3rjULgaFgl
ul/+0W0ETn/FokN86xwXos4v5gX1wVTp4TaVesaNKriaQclzAlnKGuSUH2+g
JCZ7iCsK7lEQI55rrfqUyzHU7+hY22oqJfePM2S8bl/QvNxxKyFj+yplIABW
orxxDc6xE6S4AI4PGj4Vg8Q3h9bG9kWkubz5btDnF/uExtiIoXeKVHHa3U2z
mi6snNuSJBeUvv0vRTW+phJ2uFQvsrRODi+vDt0xJVL0wjeyuz5YsVNd+yCN
Z5Ci6ZCHkzBs3CM56OI7MuuZT1Q+sCIzjZEf3/5gEQ+LeafH0O/XIufwaTa/
dGdm8zcfji9HjnkM0jBS1SV5pjwpGJjegbzb7UbagXImuA5qZDSSwa5/t6eg
+8BUbeaYxJmQtP2mMne7WWvdLQCXVL8K2h2IPHdjS7kexP6NjBenDTAmm06e
/FjuoBgkXKGqafm7ckB8yb0fMaN/0P8u8STmYyWEuAWZ3F5b9m+mGOsPZBlH
69nG2yiWO7Bb8AfkWNwItaQ1BZk+OFjPvsi9xVHHKpBdPJnTE+hSW0T4+HUD
/0UnueYXsMUBINNnSSMDOdHcw6cW52cbTtbkFVUzfGWLoayGrwGBB+6L5Org
x1oeDoaGbZmzYXSkDGT6KbtrQHX8vxD0HWMGkBfnXDjaofsJ6R3M9uZCn8hB
2Kq1nlUBEUGaF4snjjLK9EtBt/kniofPCTJFfCDJKroTsRsSzmq8R6mUNtW4
Gz7kd0rOV5Vto11HNw1YFKIjwUfady4/cKsemUWyhsREFm/S6b62dCHqW6c1
yvjBSd7zYzMLgrisvb8O0eqMvvExLqJYhPRlvVdliTd82o3ETt7FwJqc/ncu
GZ47Xc42M87XwPbCFU18jFBz79bBVbN1Gs1q62iuuYk9cIIgVmLpUidX36E0
POiaEfFBE5hQyXk59PNX7dlUszphmm74y+FEIL+f6wm43McemTKCiSo28/Y2
04vcPQ9PROCLdtFgVm2RvJbwmbNTUv2iHcpWpi+Yym18dsXznxPAP7PcrWSk
8ywhk+gQGgho35r4P3TyEKH8sE49loJqY5tv1uQh4wcmot76qZ7l/iHqmfMW
t9XilnU0GDLVEqdMUixfNyI9WBqOH3IFxiXGufZng4loxjDHq0bajiMw1g2S
zQrri1p/j3fhiHC2kzfH+LfsngX/+TouryHEFcu4YcwT1G70e21X5zez20uG
bfbFhLQUWCJQ/wI9bQn2k5Sq29pCopI/4GG6JSBnQl7qFvuSH+vck+9wzzR/
ZLx1lnHMqzaARNwoPCG0BRDO/goy1AqmVsAJA+DqfKp9SdnOgtoe36F3sPTv
1Pempsolw1oupZqlxgmh3B6Pv/v9k1P/mdJct1gGnfiXB2gTT61p0HdNuRP5
yFovw04ddHB0YVA0PD2EbF2XsB8QAkWKhzXG6OC1QFAnC8Sr9F6hbqBteMJY
N6oDEKPFRf/Ce5EDLRV7YmATHBvSOa73I+xRY6loQ9pC8cGWPMLO0ITpQWvd
bX95pYIN+5urRMgnwzqgUvLIQccXLtT8VS0+7cTcsmhSBurYbpztIo9s8X9r
2eWd9AAjPhqvnfUtd1dCTKRAdA05ri7fvOkqYNabM9OEnP0/gZ8y2SmyE7mf
gl1BSFlBEg78ytNIwvGxvd6s1gzg1A3H95KGGebURhUKbPhIK2KwFZgcALtC
vWn4civaojjGA4kkyE/kQZsePhERNX4Yv509OjWdcU8f+QeztZB5U6ysSn6F
apQxqJJGvchsln3P0uQfeX5lbTFzEZL0jmDAM2KpkiPgcCsqCmFO8cztqlMh
c/sS0TL3ZIixj0hsBgs/0eyEhS4FGo9PWqq780f3uQB7iwxqzYiB8gl7ps0g
NqvFnKS4DqfEqgF5VQXSRerlmahs0BxTQ5kezQc2YL2oTvHiCLfmDZW8UpBF
SJcAqz/siw7QS3J5KUs4MjKPX+UtRqeBNdJG6M/Dygeb56i+cd9L/pcRstJZ
Kt9AGAVXJw0jEgI/tVk4QBwaUrEl1gKSH9lv8duL5yhk92blBYvwcj9ilmos
I7Zz6si3N7b+hxWQXYrtWzY82TzvL3/hvGrcrrSdZBceDHDROqgzXiMY2Hbz
hJxJt1hIC33W/tIm7IOPEBU9oZZcYcnjszmpGbFjUjoSv73GwI0WQ5+tLgev
6mHPcwR/XZZPU0o525Of7gyyXcz2631hdTa6wKGF5RhDBOCS3HJIM1mfYWGk
7rpmQ18TjKymCYiwi0szoHiNFXqRrzIEc9/b4Gg8gCVZ5P9kFOQcT4oocl+S
9DptOjvUj3OawtyZQMoFGDIupwAAuZdiSCuyCStBgj174qZGijBIsK8Z5pva
qa315rgYSqKe4QR8LVqd4WToC/haZXzUADQIxft4ucRorLYKLuGKWpLRTkQP
AFZdWct8Enooit1951KiMnypXpMuhnuoNnl1MHb4ersIeIdjlfXp1yPyBesc
ix0Pl03f2fF6q7Ihp67DZCq1p4gpdPybPCL6cTyt6g8NVwLsdNT5Popr5vXV
dus15zBwXvZD/oc1/geWugyASL6mDAspDTtYD87pa/KyqPBT5iU3cXWWrn7Y
7RnUUKnpUB/fROmm/qtvL8jwilZk7XWdPxReHkDlAgaqwV1iTLr1W6isgVkW
WEhGHPB6thl3HI7/JGZl8tghHawtPGjFwwcBdctb5Alk6mruc4xg3oumToUO
EZAC72sKlaDtMhYkb/ToIypKWfoN2YE5bKpI74tsaqjFng9ZnsAHYr30q51A
auGzNFLkyUifRWkY4wCDpoXe/11vD/7tAamcVtCDubZpHKGezOveWW8D0Oc0
dCKFAG532Twf8ixlaQQYezbu92u/h7xXGCUkeuFGrYKKF9vkMom8m6tukKNR
BoXiPzoA+yDCoN9BQFNDSZ3t7DoWP5KL/9BXfXBLUjKSClGTPtdMOyv8N+iH
DEIg+uhlEtk+NvmODICGWv3untrLPPbk3q89fioBjBAgH9TdE5G1wSof7+Nc
dym7sOZ71pQli15htjrTggFle1sdtoAwymEqvczQzsjcXW0LHoVhp74v7VEe
r8BliphMPLggjaOCG/9700I2iFUaXo5lJt30G9BiKp6wzTFUxqMmyyDW4ZZU
4wkuXx3xskWcrrG0d730SHrpMvP/W3X9TD0UEoqTWJ+ufLZSdd/OQwJD9qgD
eFdepH7DCTLaQWMypBP0HCtqyyGH1hDsVZwmNgMjD0UgNIPseDg+HXpnLEww
q2yruuXmjAilNEoPj5z1QCiMBsjnopwOIehftVHrBSBD/cGUJlYsLzdP3rjm
QCU066D0RkWH40S8Afp+PHFwXWnixxfSEgSUQA2FiY+9GCwmcyVJ+hqiAPMV
RuCMDqoGI/hl24AiD+3DG0ZQXkswoEmCFidqXQTaZsvJhS1IZ1lMvu5X3gfA
ZhO9YrS5IEROb8WeGqwppYr/kSZxM7LUj8RnKd4QjRtQSF7xv93lrNLrXehe
7c3XGZuZOpMjYuojIA7DqFr1FQE8B3pcrLAX/Qf+LUnRDHjKkatQ4P4F/7qi
UL7mj0/rSBAriQZKSxCdZnY8F7puxJSO3yPNnEohvRuDwlJ2rpJTMBVrw/hr
Rqkpg79GbdVmsWFhRpozobJWNDteHwVg3We0rqhCp/0R7toG3MC3D9qw04rq
hMVzhDRdptfNjeLNtyLfmrqb/MkUpk98SPjzaC96o0hwEjrBHkbjPro8SONg
XMN9ONCEMrFtbVACqjX4NMd4xJv1Hxqapjx/cMS2jyF65NBclXncF1Le9NN+
CUwu6t1c0HfgoVdDTY4O1f/4RF56SNqBPb6+D/BpWOleDSYgpHrRleHq8arF
FaM93KJVBxeKxPqbEfwUdKCpAaOtEPRKzxcelK7TsCiCgGEAlFdN2Gxec1P5
j2mUpXBrXmvh3ewq91ySqn9kYg/9dlkuB1EyaED8I/ilUdV20BsRDs56Xhhi
ATaIGFpMjna1+C1jBQvzT7sSRHxWZtVjQC4xaG+syfeiSGPXF5Pfy3TE4o8m
znMvfiMN2xzDunXOrcry/ZdPiNerSS+/eQKhr3I7C4Gzlj4bc1GcxiEF5oqV
w/RJCp/YoGNEK1s8q5fxVKIsyGjM2pglbu907mV1AhG4EsXdf/GPoqIpTNVh
vvqmsKwgWsn08AaXLznltMxINtoPvBLMRquJkkQDVOEEhO1XOrXk9/2gRHIv
lIK60lqnEWMNjkIwLNUPDaInKbtBvxOaS+Zbpnj3V9d07CsHbRHjmrtMxixC
NJePy/O+UsivrU7k+/U7gsovF1AxcPdJgkBHdLVag3lB4DnUVa98IBaQ4wKu
PyHppfopEkUEtdDPkDbzLB11hEeEQhCEx0PkxXp11qnvzZI+T9M7Q0gz49gE
H0ao4oWpPVwFrgEJWGPQACKt+NnvbUZeF+xi/j+SN/Ho1/4R/ao3mEH+nC/O
AxWTkel5oov1FUOHPJL5pjdDQh/fgPX/edIecpxAGlGdYaEWVSZKmfxzeMqe
vlILNsgMwlo/iT/JykpIjdPQWzAMfFhKKfAeDZU24w+jK73kjQTVV20wmxe3
hOuKzAnviU3A3ipsbLkJUvECSbGLZZ8yhn8Ub9WBzjBiBsTGualMcEhqhsbQ
P9nfhxUAbaL/YvBHJc9IBkEi8t7bc5KYUOqJwS10Xvxgf4Zaxi5SloBXKf4E
XxV0OVF0efQS458sT9Gfz3f18E77JcqIKu3mWNYHsIiZH/oDaHXjJzNg+Uk3
09paiPkxXjrYG41f2LHvPEvTfkmXrTh2apPgzWjIxT/iNTwAY0HZKccAIi47
jll0g1xp99kG+49R6qpwUISnrXXlRnunohoildtpyknIfokRSsKFsMZBolPY
mtkNdz5sVFuNIj+MI98GKajD8zCXUOGH6dzem0j97/h/L4vNxwNlEK3emhiP
YLV4t3tlsNKoHjP6VI1DdEyGkwol4Y0bVvrNbzNTc2315KtwUcRle3XURt2/
VGvHPW1g1L6rfA6SR3GauIkwgOhHfN9y2MLNbOdwd3DG+UEKhvLR5KVn0zYD
NJkG5hq0Z8hpY7xRhGYU39zLJc/clt8yMrw4hmoZh/SZgDwPjVfgx6Lybllm
PR2fd3O7jcX7HuORFdxmsiRT6A7niPIgqIyxyBPAWuSW80OYI5PfLwQS+fZt
LsxUH9C+KJRQpR9NsxJqvFVeWfSpbsQXsVnx0mUT3E0iNdnMGJuKIYkWTXYt
roV4JPkgHnfZrfleCK6uBI9ASi1Vfgei8XWq29UR/D+KXro8E7Qx+UcmoO8t
WafXhaS6JJqASKTRBXE4hq0YW5/XRyOzxtujQsvxJOhhgcyjscN7xjJ+inS6
nzp5Rcyv5dc9/Wt1NwRn/x5KldQIV1pj68eZ9E4OyXJ+zqSAROfDV8KNp2e4
xcmkQJO2AKMGHzJ/uTXIJ4e7Y/b2dZDg51vljlTepikaafWpOrMNRIfxwTxq
k4dFydRpEtkp/rbQn/NRbdIJ/bS002n94SgorP5dKicDQcmXwXSTPrpZdCNn
f4ZNFuJTZTEVKUfCStTmRfoAg4QlomqtaLSAEbfsWb6L+dPq0gfInpdek/wK
2IVu9AelLULwARKK/BgSaxS8MPAyGM+vQ0JEt8ZjryY7T2uG5Fma0guMEODp
aHP99AJRQFKjbSUqiqQMa+xL2+nirSYj5VP1F6izYDA7dbRem4K8gWmBYv84
ScDXo9TyUqgMWtRO/+XO4TzqznVuG6Ztiz95ng0WatQucXEeNFHzkwWARnaK
/bCLgcoLILCCychBdpGMnMMUF/CjsYwQj+khjEVLsO7vJIClHnDoXENOguai
Tv81XVk59ZJXqLBmjsE5UNpMDuV8GxHJV545L7ibkbe3/ioZ7FN6Bt0PUvu6
7HF5ey8E9+ZLGlgfXiWsHtCGe+lvzpmBpAgbIsl8VLPrqr/ters1ZSgqIXQu
VR0MkpZCLJ+F4uhqX8AuUXrw6mV9KJfhJzxqvEBPXpCcF12OPpa472bbfRKH
IPAbswdYpIfJaX4Bf0bG97cE2wApcWrWrxxEUa7PYev5r3inXsJXSdD0ikcN
asP0lUjth/8hwepRBKXlXtGOMJcZSl0OdlO/BT2tnb2kJzXcRTBDw/WS0tIc
qglILKilGdUMhCocTUTHk6XOh/sKqJAk/B/UGtxYX2Y+MguFXh/S4TyalHHu
fr/UMOTFaCra2CZtMsRRYbfhndl4+pU/t3u/wYxM5OMkf+OaxfnCmR0ERH1r
kJEt04HVgMlW+gVuxdFWyNHUt27fkYIviF7z/ZVBD1xdIth+XgUBLTGxM/0O
FGTHof5g3nxVC2kFMmERWW7U/ZbuBQT9v1m1nHSMud09l9eajO5o5wcxQGEg
pkXxjNLMXdomyM3ro958QL5KiryOBpMsu2L1OiFzWATfJ93YUsRzcDTEAQnF
pCqCRaJgYJHq5vR1Jvybyae4YjWqKsnjdCiWV007oB4iEwa2B4PinmAWZqlC
8UMC/oLZe8WU4Pc3+fnHptgsu+vcQME7huSLS8Rp/uqdCakBPtGohsAiycSa
W920w03wUpzkJAy19WClDr3D7dwJp5ZcmuJpqW2jZrQhA4sMMuWyaZmgcQav
7oWUtJ6lw8gaNN1q1TL3I2qX4l5TdBc1Mu/yUElbO3czTH0oaWCTLZ1Xqvhn
1XO5YwVNvh4vDaSv2aVaf0p+RKWCmAgfOFSAoRN9ulPeyO3cM86Sq1AM2Ffv
J53QYGCbJt93mbXK3zSYKdtNKvp0O9b7+AHdVaD8UAGAn7cU7H/oJ2NiSIeE
fDNxvjG65wq3MeHp1opanT0R7gfb1D3vd89fySyyrJC2EJavQRGPOeyOjx7r
ettDp2adp8hFOunmfORxeFPHaDcW8moR7cwcfbZcmqurMQK3wmVtGGogP6hr
Di7RmNA8F+bZKsgS23PrD+mcS2dLickeugVhvLUx34o4SqJnmgdYhfEXvaCa
lrXVk1cxE4tdLgP2dgN52CHTExy9QL8KK+smIxrD7IccW6yo4m4itlnIf6Ef
5SA1hABd67jgKdJe2arS+nI+rF61+Y4cR0xQoy3Q2cwS8d+WfIJradI/GTGY
M3VQrNMQZ3PyyAanBNy4jkELMlg/8yxdIZWpn6wbZMCeqaOYKE7lc1bbp/bR
FCJqK2NP5m+8EVXSdNU/776M4Zhaml7arRKoNbriPoTcp18D4nZRtjbY7e79
sle3NQrEhXs+X7Y+Qxb63sucks00FhBuM7HBORKZA1eCyXylSQqtzlIBMZRa
fl01Q8nDLAVfmN/rCV8GoL/kq69lO7I2D28QhWqi130JE/Pvy3l1Z9Sbb1Uy
89+RDCqZynR66kehcM+RfSNQw7MoXNbRCeDJ+5Ufk0S2S38KTGqmBG889hAE
dduO8X2uSVMqfrmjx7C2PEbDxI3W32gH7k3kYJnMBQY5DzT6IC8Mwd77xwjt
JZIaZ5/Phk+tnfZRQUm8I6G1NoDxDoU8sHUzoNFQOIjTov7aypzX+xpJvnMI
Ag9MP3pavBZ+DgXXHPUDaImlvOVJK3kommj3Ha7dFcxuDECgUXGyKGKVDYOP
e/fglrmU4vCc/fZhR0soR7S2AifCY/Lz7/67tHBf1QKXhv5xge5/K1cwF3vy
wP664y0u9XOYJcCzpl1Jfu8Q2oZt8V0Q8ky5W6P9EviQGWMwX1mR1p/saaYt
lgu5x32ICKEv20rev7M8Vy1KEpyQgoLGmOJZLPyT4qNG8jqmE9hK+JY6NT3z
ooKULdpfX9kxevWhUjLLJH2SUYpZ22V2VRGGvvyRg+r0QO2j9f1q3uLCoqLu
GzO3Zrb/gZDszAtc8+PaAmrjl9vHVFboJ8rkkeZxVWMk3LKMxqvHni3PZdcJ
pmfQljAtldH2fA+Ivrb+BLk+R36rylOULjdVdN8erVgJnMOrM+iOsWy6zDTN
hEeQ9tLblWaSdn0ylUc0X4FIMr6IJzizsKedGg6k8qUaJDdZJhJiuvsi1yWQ
djuXFWkFuu9a5Kb4FwJvlq3WF1wAdwpIdlMgy1900eQoLVBMYWnixfEd6kyx
QB+BGgwaZ5yfDOYrA2R7kcfuzIlOrkAYhNapF9b/aat0LAyEMrVBm+ZhiyFQ
azVthDAiISPmcGynSUvlUsChEatd3Hsw711O0kfLKPvy4vact6/tdvxCkRg6
/RnQgGYQ+PnwO0CwRNMpNe1w59rHG35y0dryMsGz24tL2E5dTaCMbS8mhTfR
OTh2hjqtEweJ2lqaSkDw9qelVSJzRvCreXWhAQxJ0OWUxZjQJ1tDQgJHFgqZ
FD96WfSroco9ltlODMxuf5ayPn4yG+Xh8RaugdUfos+Y3dPT1Xr1luThvl61
AOnEaxnPvws/SOrca5v0Q56iRXEZ5nFi2CrjKPv+3J2vTu7nO70OgOenW2oq
BgbUQQZBEp99Z1lKJ9UD5GnyyOEDONXKIv50MLOcugS1yXzPtDhjQ/mrzKeU
oaXjPovTzlxGW7iBLm7ZVwh5X4RUU/Qu60ra6HbtrJhVAWXFoLKuLo13NzSj
6z5wgMa5/lBv34QXE/ifMIAt1pCSSqqWWniJgTDhroRhCAzDXFfxQoOLgqul
ay0LpW4zUGd9Eg22QLn6fy/xPqsI22ecqOKMQXa3eMzxQzqcAz5ykEqxZFlY
ifU2eY8RsORUDek1xM8I8JveNSawuPqIm7bZulkf99TXeYvrsPstCiIyeBNb
nPiiY7zuhz/Jg90Uk/qRv9ISRqmTRO2ItLvoQTo2bC7ubH86d3rX0UcPcVWZ
Y0Hi0HJKxsyESN3JL//4PFFfh4ndxzIBS+daUbIRDXWtnHPkL5XnCuGN/+SG
8VN0V/hiqeu9UgMGOQlW+3/XR1bOjyqKkijqrsU8j0o3AkeCmGs1bqhrSpPn
qFycPKNGTBI732NM97rZxi1opFourgRslawqKqQWTH7EdKb1z3Gx2mTp3/QG
Al2ebyqrieNfe1dsPyMAV1zy744hApBCsdKs0AjxZwDoz+sT1Q/tstcVb0pm
8bjG6of3KaKeTPUI79Zu8D/fznUjtqqgvGxNHjBqqgwZVghCk0qWjkJwq3hu
XFUFLNX2+Z3R4XVfrNbnh3wBWZzNRFAHIN5bz6isoTZswvouce/NkCIw4oo0
VUoqRy2ZeCsV1BF2ahYskUIqTQ+kddaUS9tMGVRtcpVt1JBc+EJrLpeSmR2M
DAx4ZOPvX6oTNPLRNeWs0UUO1S63qqgsVJkCUotxQwX4nZjoAx05JzrYSjEj
D78FrXwBrM5OWU1g6UdXJSj3OaMLbUmVEjyVcMgfYQXNTpDtvaPEUABrMGxO
IyRhcNGp8B4vRyJmvmbON4WELSDTeGJSJzKTP7r5pz9REE6hE54DLrLOh9aF
RMaQVSC4buGxNaVv1LVg19BdBV8yES9h7k0y5yTxkqFKDPWJfFG9A5yCY7Jy
Ff4q9cm0wwvBDYjHUrksVNvlWR6s2D+jGJsEU4V7gyO/ZEnQ0xgZCIqYtujz
dLpKpr6gBcUHOSL5HvccGDt0itMIrowpvTi7/tVzaMW2Acd387vdQIsRSmnv
vrvKGUnR2emptIOlfEWNWvfmb9Nw7hu1RWhIbGbu2Pl1UoNB8GmO7zyN0PyH
2grLJBVYQEQ1SBpE974/TE9JmLFR4pbmfqXqgBXL9rBIK9aOHmsxXUL6j6Jp
qpwYU2hjb9nnio6+HCi0v3gZlB2JPfQ3IyCmC9KXMi9+DYa/qm3av2gibPz7
XRR0v/tlSQLFmwjWFyOM8lKZIoJAdwYyJsS67NuQuAOSpoZS4mWyCSBMysj8
sdTIWp3/SR82UPJE+9S+H/BsOjC/2CW9ct2zLd5Rh0UTPxrYdKWCfvxasB7q
zTj6KevNfPvGOATWHaWmH1XmtlIM50pst/sERC8Z1TwCVMRTdPkCDnKmPh4q
RVHrNYLHE9BHlUjUQZRGrF01Cdkq3Czls/SyVOfMBaQdnKqVSh8S5IGNqQYY
3uZsQexBdLI0reHdEWkq8jGJURXkboNldjGz2PWiIYGC4NKSpiSc5c2SmCEH
YNuOgW4k017Dv/z38CtlnnjyYgyby6k9Dns1vDOmZfvYbuSjVreYhzxdJ1ft
WKkac5L3OPNB8jve17p9szujWQ5isqwnV3dgpS2YwRZ+aRY4vcY/YpbyEnoD
ubY9JIwSshGPArvACLalt3mp9CuakqQXbTr4jL70LYRndPxypyfVfrbQt13r
7XjWsOwg+BuLulsBiJEwVAc+wRMa09M/oZVAlKkSPebyWCLqTBEG6BRFv2A1
C2IpjJDlZtEd/hoZegtlSUCNvm3iBKdbwBBijhal3GFh/mWk8e2KnsG2+nys
UDo1+yFtMkV4vDayh2uShW1CIp2OP6SZDGLH8H0J/DC4E0w8KA/v9DLpKly9
JlNPdnpkuM1eTYAGgEYK7a5qwbO8+LBVNqOP+tNNh3Tl1N0bNyT2QzpBo0Cy
DXhVXFMYrpZ2l/ivpFbBzITZjWUgKwKb5muH6MbaQBibkWkFhx+V63SmVm5y
lzXC+aeICuSJEw0Xt/S67kPRwNJ2SH4DY0BSUrMR90vNhxNPiDkmIxmfUN/3
hcjgIHj7J4GCnNceVuVe+TKwyisOZfyJbAi89uzUNfHFC9nu1h2mAKJvyGV0
Y0AJSxN1Sn6EPHjwivtRKr+lUDDjEwcfso7bIlZBlZcHZR0KXUGygfWfGTc6
GwHmDmQYyU2LWNHh7zMVEVLNmALR0c9YKBkYf4ey8e0EyCO1wFgj9svxc60B
qH1NSqjzJwl0MbZDiJ8KXdCiwawoPh3zdG++clNGcvgADkmYybBRk4Ewt+bO
VorKXzy8DglyeuSz8ol8+68eLzsZh1OV3aZ1UqvRcVi0K1PB+PQMAbEAIBok
/LGWh+/tmBnxH5Pg1Vk8HTHohKJnrfm8vby/jNDf8wW7zcpI26RHEXCN4cJQ
CbDrJRfFtaxAQ6T/qGoGAUEAGmO5Y3qyvo9FaZgnOJrvVxFL32gE18KldaSP
ONT2VXBk+PSmO9dslySEGytVtDcfbn9rnGLmey+sRduusRyP9LrJY3Cxbmce
pVxLTYc0AqNU6UfOVi5ptPKoxVkRRcUwqzEd48ScOq56h3+fH70QCoHLeywJ
MLXikv2zQRaXyIF++eeS5F0dkwrQrqFUJPDh069MIyHTDcLqYQ3KYxBEMNIU
vdd8SXIDvlxMVDJEfFPx76E7WD1ZGcNGpIq6L8mgEoHSH5q7glrM2+4I5ApJ
5MAPsyoKHg+we4zEao7SY9ui2B2BkRGrMfG7W1V9FYs+7axA1zJZ+GaqaiWN
/LatZJ1M1CvsRluDRwQONalGYLZAFiDGKL+oFZFCHtQ7Dr68agJ4/6tkV+cD
SG4cFaLwjPKNFyIOjAeUsG/sZPSxiFiMPACbLaRMutz9nIoaw7T+IWgsDOmC
XFLZ7+bk4uNi2KnuwSflJ2GRK++m5JYAV83hDpk7utsOxPJ5FMhCI6zWhpSr
CbBHtD8EH2kveEdrZYVxEsRF2hiTLKpezaWmXnELNwefZ6P8Um6uVDHGu5ea
PRbGPECYq7yfnLrSZZGXB5rAOicgz11d+ETUL2+OVijBAUtFZAbOeMuJmS6h
YzgOh1/93y0HBilZC4tvyESga23FfdbaOAJgHuvp1aJd17xh7y2jD7HGXEeS
eeTN1Ly3VCM89znTxr5tAdaddK06Pj1l0LMsNTXklvnY+YPJVyjglifpnzsF
On/KkyzDwJzGeKdANF2Xz0tCLMg6sdjVNGcNvkbqfAr5JgAacAjIedNvRvGn
tC7h2Au4GPtfyDDI7g/dwXOLqOi6jpptgLNIUccUYBpSyy4nKBQRzTGWEvIP
12dw1X43wwNnHBmBWXpd4ioj4nrHqujHFC9ES5EqzO0Av4cQ/XmCdhksVlO7
Jnd43HTP+jUmjpIJGdrA80e9zyWYTXpuuV6YVjWWT50T88B/kEwWJ2bjqHsv
Nqyh8E13pJ35a+i30ISafY8moU2gzZJBnqhHQuEt1lO2AJcxkcWKmx3UadKj
r7osl84hkwyuR5+J0UeV3xrY9MkJdIauxc9dceootIK0JbsTUs/VFamctIjL
hwBXah89YtTIdCfV5YbnvIotjgx8s1jvfslQKTnb8TVZNVgWnk9b6odemoyP
Vhuytp4YveiMHLNy0tJuVGH+JWflaQXaOfPSidM0sEIZxU0cduSuU/bKdA/n
5Z1hLZe60Ve4yV6NA4Oddg3shu0qlHYLD2uan72E/PW2+xJwfJ91ujFn0AQk
XWIZvAQ/q5L8dArVyjP0FXJXo3aNN18crpvLco9e9I2fyiC5PMadnUeZfQ/C
BeEib6tCAwZoVEJRGKNx705lA+JovC6RZVChK+FLGAJufSmCLYyRA3b1Uqi3
m4eMiuUwRcVl/v55owcOX/eGNsW7Fanqk+njdmGxOX69RDu8pxnyYMT2PeLH
sC9V8rdA7tPoHshjOoHPnLNilKpTgp12FrIYoqZtFdJpvJK6KUZGhRNbsX+j
5trXYPvZncnsGal8ROk8aMd8eeffjedZ6oOhMDMhaJqg7KyLo3tWxr62YAlg
v/H26ZqSpLpwpViFWRBTGFsrDm0MyHaokcSBwt15dtAKQ05+mA6HWLY//Ux8
xaOq/dyH+AndOHy9JeEjDYRmgkYR/w8hskMWEWwYJiLznR/1vvfbUXWdF3v1
JKFNaoavR3FDa99UABBiJxbivsV8DKRQEprAZ5WWoPP2yrTR5MeuOrqBi/qV
WrK10buyRHrIBVBFFm8Yqub2EMjzRVA4JT3g8EqmjWaU177S41DXYHD2jw1l
opAkPcZnMbo5hZ6rFPtW+i+ayQF8I4pZqU1kRaxV3eYQiVP6fv1uGAbsQ7wp
ZmsOX6Ke8jF1957cTGQltmQxmcxQd9geENZSrrICxVykDGdjJ554a4W9/dot
GRUqdJKswgJ/OaKMSlHxRkJ9gUzpcb4cSa57kDcC0UfS5nkvT5bexLLOXq4y
5hvKo9+sgIck/yIpbdd7rMuQTxEyVYgZkNA64qf0vtMvTDHpWqGRn0FYbUED
+Qiotd3tDBQE8swrGwowhaU87ypBRtd4s9hnySW3HDIg+KFPisPBi37Yt7N9
m6rWHVxZOQbF1tIwXSC59JjqBpsczxlKcwcaks/JtWOZVQUGEcw0xuVl1hRD
Nw9YhJAMsaDf7B/+SFi1fjfbHjodsVUgpaM/e5r5eKmvJ1FNrGZEAOg4yvTc
fl5bWZXjt/Dz5nfkdxf310m74ZfExOjKWRa9argPKouT8GIhqVAQnmnFKpg1
jilOW3GZPjKHo0Rq9Ye0yTcPxrGoPKAdaqqUldtbkrYUg36BAX4UZFvkHPHX
ee8CSppsWo8sQgkfK3WgfmG13bdOrg00ZrUyjgswwNlGUbD3IsUmx/CBV8tt
zuOiBrSTLeUxYKSgXb/LTOUnPB5J4RtY9XsrhNEQwbh6dWjFaGw7abHYd7u1
Ma8ALYojb59lJccSG+N1WCTxeyO9zH+0Ph0TLrIGzdBJQQfhgHCCy/mZPe/P
1IEvCi0W/Ni7fuHl0cVPYQez2lJ/JNj0kEdtRxIjQ/KkyGOKFgtQ2PXVbwcm
7sZFpSL5Uo7pKy1mMIysYVj7Z7tmAkdKetKi+oXkuvH1zobJcmkYDQi4GScG
ToBbjWfCQ/mqWk6E3Y/f2dTojpd4R6tt8u3mzvjOukJDi2LDJsKF6lh35uZ0
WgOp84qD1IshsUAnurecH7JIMVoY0Adq1o53STWOcs8dy9/xXh+yhr2EgRfs
jJDFSgGoMvFvxZBRRODdmYQwJdi/l+epoyLs4RoZo3E8jyQ2D/9oBkh/7KU9
E/5k1qw4rO5jI3xhnm7Bd3boaSD+QHoZ0f1aMe2w9kWIJeDXVl9UV3Aq/G8f
h2D9Ld5UF2aJLXZnNFRP/734yzDCkbjiy1QBrMfCx8p/IYr3/riMeLMVlZUA
qTVOmlW4eXl+e/I3bCgk8qKADrH+JOotdjorHKD6qISE91lRjqQULhXJ/MHG
mwD0U3GVfYeRP9khEoCesuKTZe7VUGN2X6Qdx/Fslz/xJPGYZB2Fal9y4er8
zTz0EUXn29ExVtSXKa3hc6h+q+31wfCCad97x8YvvSD+Z48xdbJdbWe/AVAn
NUz8TojjhDBAjAJyUABY+apu+rWiAjokxuMIndZasnTJhHCYsm0CnB8NfRaC
pppiUndWuD/tzxb41kQL9QoX/MjHtWr94CnJ06Uh1KmrqNIJN59sLFZlOpPX
NavVB0YNQQYobrwjgtwVDbqjFI99vlLBC+k3GtrKR+CgNv8/yZliIISUeIzJ
BbuT0a4ZiGMQk5IpcKcKZGCYXtynu1FU0veKdSyw7sJtfsA/qJKTNiFe6S+z
0uXT6VzuWebWWSY9CSLC7sG/Vuop/qpjrrjJVLjUj/dbO33yHucbBwhQMmUz
sDF6GhLqCQFT2j6cbGmI84aOPDtGFh/Uf8Uvy4YEZypvHsSAZCIbk5F3bYli
v/kP2Ax1BB2BjaBGCFSU2hfc1XaPCVC6oRwUKYBBez3+LL2uGNZKH5VCcCMZ
iDroNam91JoVDEpdVkLLb6vM8aCBqkV/ME2guK731ifdsdoWP56bxFxHGbPh
LKpxpWhNSUqIK5ICSEiGHHQqbtqxtYUutgk19sttkzo0+aJ3JHj2m7nh96UR
S3OfQ3zdnMOLt40U/W/GUQL+PLCtp/9CDEXSOaHzpPVIgtDj37fFDiqxbF/V
ZVvLBiyGGW/b4X3wqeAZAX1+STAgdE2ArDF2S/ThTGLJtja6ZHXMZm6Ta4F7
+WKYecbd9w6ZsrQR5fAhnC24BypDJipDTHHP4K/pnLYRTCpFZkAxIMNl6UZL
2rChxVj1eaJcOQXecY+IRE2hvCQALqh2JYhGg2/+GMmfODSu1+EeU2GcTKxR
uENsK5pz6iZYzjleqlSm1MzCVy/qggiQMi2NMZaby3dnz/LqSSa8v8+Z64di
zYSjChBiU7ph8jWWsyXUkWka7dwzigRkxzE/RLDdHFQpQM6ZsAKuz5fd47C9
qsLX0nStEgheqVlsnLbgXiJVZt4ZiWbmX6RI71G5z1RCj8W/AT4/AwoBb467
/QKvXkGWP2T6dN98vSLyyNFhc5f/S8HD5UqIJDMG0joXKIh8pHtBeICrphB9
vdtOOgEDUZlH7HU5PIPr/AMNPrg/l4izz0AP0fPxO4Xfmgw3WF7wpEZKm2aD
40Wq+XrljfAKaz5H4JFqOxPdWYdzBOpMy0QSW1ek9Wy7IgLFjsZM3Xv/XfpZ
LJ7394A36LMn8oDf8qN02cM1XS1CJ5pQuqVEjHwVo8YIgCQLFSw+SxFEJSvW
7YEBOpB6XKy8YQnTzMGWJWhpU4LdxKTj3s8c3ARcgtz41JoonEecD1e9DNdX
nKfLlLrTx81ctA7BBdW3nes2sdapCfh0NhkleOv1Cs1f6oxVc4OGZtccVa5T
PNeeocJvsQFhrgYp8Cdvn4Qax6CbaHgO/KXMVcfzhoQoStapA8/fX5SwwxVN
IpH0lVcBAFqiusgic+TlfxR5NQ/0u5RpDbfeU3u5v5Ow+tRWT7wyjg5jNF04
skBiAxPXRhWiygd1MB7XsYYNpjiGdCv2s+EPC8fwDO1FmxvJAup+bIn6Jj+1
pQGofvYzXhe7VHvc+3QiwjfMuXye0r3rZaJocuc7vP4IS/KqFMt67IXrbvbr
fpGUEobZ5dFg0sNvKiXSFCJgdZ9orxg9drdRck/bkM5plYBHkUbVOaYnzfpo
WDbF8jAmUggl3ZRgCQ9AO3rWbB8tMPpLs3+RenZ9GkX6s7bR24WzOJjnqNWJ
HU0jAeH6b/DlwGarkgvb7sLjf9imYfYU2zag3jIz2210BozZdDhZvlEzVa43
Y/jYoBMcd1TFjOqPq4SsjNOAONTWjOFdT3e1ovk6seS+1HntQFTGBDFEJsHY
VexN7RvfNOdvjIFtt7nGBbUJIym7KoJs7KrIttr+JciTLHelm9IIVKWx8ZB2
tBDcfb4s0H2hTo5T0guD54qA3wsrHotJhVnQdSlv8VRJxRrJjqAzwKgsbdQ9
talDizjdZPMsBDloDWLBrqmV21aJ3LXYyra2coxkmdY3xaCLesESrSWFuKCv
ChnS8MAeL47RaLTjecFihX0zgJI9aBZ0Sw2m5zmknu81Ryvwqu9YRpC4Xdv6
IzyDWHvszgJac/+N07h9VOkLq//hjgcDwf/ejxMm7gBVK8axPVjFlJjw5LzG
TWhNTXWRo0++PaZFb/mYY68O8GJnlb+E4RB8tQeuU+1G9RuoZqfXsfRdWFEM
bZg968kM5i1ecXEM+ezva1hLa+lkMobF1TpOL7ceeftwcDW9Y3xMngl/DL4S
GWP+aaJe5AkK+2UhsyLiynTYKlR019VdRY8/jVgPFvydbYac8yvyA1shGiw7
uLdbEgA/d1WfzGS6YWRh1rrI/hBrAHWgsqC+lnRozhsBASKFxjL5tpSRz4sW
dUUWDvjVE6CYB1RKXt0VNmdDrCZfaLMIa/08MMThdAJRn/wzrGqT+PIIqZSJ
+pOWDk1TSdXF4MZiv1F9Xk2xVp4+ht/yWVCNiEVUWQcozNznU2ZAWm/MrJc7
GJSaH8DsAzGRYUx/JNup+91nVQMhMJ2DLD67c7mqaLdhV4mEPO1AFTOTdDP5
rS3oYjXjsJE/E1zzMTO2yiF0zgRDVImd8yC27xB/KTb9M7U7n7/4NbZm5tBC
LVIatsT7QAXH2F6Gz0muVbYHGK7LnG5tZn5DqfqZkaybFKbOUNtlATZCqvJH
kugZeq9a24tLwTaq3wHlO4KFRCAuV90WkBFdXvwnL4joxupFN14j7cJcAyLG
Pr6Gq3OpXHfEGzv6NtUUrGOLHz8JRRFZ3B0HOe7linwMfhtWmiT62VP0eNYk
CX8AfF1kEPlttD+u05Y98XgkxPUbRLiDyeHVuX4FTLsroIWIWW2PBvWbOoHT
SG7f2hBZvK16mhbRg2oni+3phDTL4SWJ6Yd4xOORtqzUBi6wRj4DH1vqfbel
qgVpz5N/IOjB1Tz3XYZLinJ/zP7J2JhX7qGCtM+Jf6OaR0Py2ka84Iy9yIZG
WV2Oh8KVX592CHC7L798DpSwDUC0ZUsGSsAHQqEz25Nth7zNpe6e3ebPjNCv
dSxrIIVyCf68p2eyWKNf5DgOv0cn2eB3zxKW1zpcs3dRJj1simZTPTedoQhL
riHo1b0p83Kg3rGPPIFoHvBURjJViPhpy9Yzh9sZHdx8bAFl/IAtS9szWIQn
+UKg2qsFd/Q5+aUKnzDgxPRFX/LsME6hE0XLpuKBKVv3hbdEtpIIneTqrATc
AHn83kuwWNTyiIiFuUmOv+HfYKYjIM8vwFeuOxS/rQzrdmwV8m4GOFI7bWnO
ikSFxpEfqzAqhO5hwSyZOMYFIH+qYo1rQk+Zk2ICrfFls1yG2Qb6oCcLA+sD
+xvRkchnxVbezzR5GnTwIFhLMqxgf06rYVVaKlbYNkNBlKFPsW7IAcvbcHrL
dAenkWYHmRRtQEeiTaRThSFSRIXjJZfIbhNUwL5GEwnYwoSV1p2HWTb+yJOe
PCqXZ+CjNu4ZcfkgSCGMkZKLssqAbtlO3rNgC2ZSqMdzadLSXhyVb1/qhvLj
RiOw6hgZUeFRuE0JyUKhwW2yVfkn4pFkwnLJ17dCsjC1Dx9Xv1PPm1bQFGAU
bfyC8RaxbyFTA6K+oHmRsNHZR4XwOgcOOJk6LioAcLXL2hQvIZbPGd8Xdo14
1Exdjcq/l7Gxc5xCjlLO/1ELOTIkAcyN9K57U2HrlQrTlZx2YIlHKFyx1sM8
kYfMHrCxgHrWgnJr4OhTDT7vEij0Y1ePzSad6uY3rQKA+7BJW885eN8Lgf97
uIJZj35A/pI7q8xvbUSQ+jSUsO2g5KYgizy8XTpbPmdzrgonyqV8b9vCb80U
bIIxV3y5/xIdaCgwEwVosYx2Yy47icUMOfMpPkuOTBhXUt+tJ2OAgqmMucfE
9ls9f0x2nNNh3/+AyPpfXvT5QQN8hCHqg9l3bZy3iJ9snADpgvdLYkhzSb4y
avfMgna6y6fxQleFs6R/P8MJ6NcA/MSEce+APRZyWz3J5Tu37RIzNjH7SIOC
5uRKhWWVNpj5PBb0uupWrH/M6WfLWj87FHknfTcRKoJWKoWKblXTG4AGU/cB
15HE5e/fV4DMt606IKbynctWNt6jbUTCRmY8bq77KAhJbrmXRhIXHKl36JgX
bF4KTBoX5jZBg+AuWoV+PhCCluEk+EdWfXGYoBq1TY6648+hzPbvPQsqM0xc
FDnGeqo1BX+WxP5WH8MOT/iiyl79Y5bDOarGnIFE66HTjJSKqxC96UumYfvB
F6VbM2FFR27k2jD2thM8p6XA7r2XdE61xDVFRzL6NbYG9Jbxry2GRtEdOZNE
cBpusv2rEv37jkkF1G9Dk5otuKsKyRl1FM2sCcv8jvD8mU3sd4Ct2oY1/EaC
52ws+IS/oBMK3Fl9epL555Agm+zPfRcGmSmaO0Y1uPNg/u64geBufmtgRRpc
fu/aaNj4KPKS/2KDjzm6wWhK8hr5ATZp5mITUFahMHY3dmEeV00iZgRWbw28
7d9sqxg1aWBp8ovKO40H00i01lFFIi0UkOW4RutdWDNPl+pqKpL4eUtd5sG9
zS2ywzgL4Yoq89eDtJTFDV9ZX3qdsDr7z50ksKsAZAS/kgh30LO9pS5oh6WH
3RlLqzi0+8x4gYBriFh1sVe8zxUbr9uCenpDj1X67Cgb8IySRO4IOL2jPfDH
dOAL0OhoRqoD2NP8baUKrcgRrdhRA7bZMGKU4cuN31CeMVcp2ME0IRGpu8ZF
uKP3LFwn49EThFwZL+0MxVf7ioDzsn8/vm8MQnMfq8GWfGXEBDtisSwQ6X+Z
Uw6KUcRy6g9+UAeH1qgvBZa6HDRPd5gvouF8J8w91MPWqY6sauIodp9LJLjv
pmW1ERneG0b5EKt4iG8UkyUlZmmOKfeH0rHa/tK6mVdIjlmrpObUGdaCHXBZ
n27PrcMxz/6fQGA+e13vp2NTARnOr/f+m7KKpkzG7U73/mRaP2jSoFHkAhwM
R5me+XVkBtDO+aq7jfA1tslwSh0zNQBNe2Nhf7Dh/VuhVlAyzp6+vPBV0faS
4v0KwYFwJzfE4nWLwlYT3UzBy9LpF6OZW7KnB2/2wvhjDzjC3rT7aF9kqrAz
2koXagq8lu3OEaVc9wwfD0G5k6KEHqQ3mAI46lRPFP9uSuw+yyrfEzwkdhas
3e+ijGSjz61imGH1vAx6k9JS/B6rXpnZ/u3WuBufvaRN02w3J1ZpELZAhaXJ
VoCEq3TWHU6xSucTYSBhZsMAKGj8ibPeJdkl8uCSjb4UD0S+qsYmvhsETkd3
FSQSbwFal/JbHwvYqG/ebr5V3vX6b/bqIVEH8tLDSwGAZ8CY8UasU1WOLZDe
5ljvzRtCDvd2sHE5HAJ123V7J5q4WCJmMINzbor8lxQWjYSJhtuFKTdjXSxl
2Euziug9iF+i95Vr0E3BGughw3FeAR4CNNxh/W4YGc9ewMgFl8GUTv0LNLeM
wOYX6UIhBSM+NanFan1i0cWm6Mj1D/dkx+4EU3/gqmyf/C+kaFM1gQgP4IGg
TaVdniDEMPtAHNUl6Wl7LBaGuLD014mXB7YEMz5a+tFDeKX51jSHYKXB3M+I
mqQdWT5kcvn0Z/d5ZIB9NvPy3oPuHS3JO12+9D6vU+j24VHZ+MAS25mSEXrl
Qa7iVTPAc6y5BNZJKOqqTa5ldhsqDvhcf7+T0OHTeut2FDVS5pJ2Lkd46G75
wQthrVILUoQfTqxUx8GWQUhEhQLKuqrpDddzIB4mYTNlED1f9kLK6q2HUHbz
+vrt3co8n9yQsfP8zGvd14EK7lGMl4MRjz+D4a/Fpi2aM4fEGnkBLUrc17Tq
wSvBhpZuWkEhEy4xHIvuGZSR6AxzXoUi5HnLzyiWFM35CThIilOlMN9H+0J1
YkGERLtwruAx1YZYJonBExQCs66p+Tt52Aj0nIdxvlQavjDmg80gJhd2CsXt
JQdiqgLHD3dWI2JurMHB76LLDEt3aGlsnsKF1btTLvEejr0svaCmoDLs16WW
BRhIcuumFHmxPri2FvCDocrMbgiS6e7S2rAGNjf0KRixB0JPHbmpMD/mfbMX
iRnvFq7cfEX/SJWSJan94OBCt54db0pbzQ4hE0egRoDNV8oTH99Hhg9BBBFT
7KBunYputX/VVavzNPt2PLFB9O5BhTqTf/1NdOXEkRG1EZG7TnRKwwL96HvO
ZBE7IIV6ODjKi7etUxBrBX8K6FLZj3bH5neCvpITHodO9a6jhe8aEwJmOrcw
Ig1EvTjM+vE1wyCndLhUkuGqIANf0umJHuxsEpDCLzluCUrgWBu6xsb8OQNb
711kRgHAsB7l81UcQXGxGdE1b+K9WFIOrw9300rMPPC2oQAOmw86xiEpGCJ4
QF9QVY0kCFN+z5zU2C9Z4zdJ/Jn8vAdglQLKDBWTJzQFMhsGCUGWXTvZdtOa
xf1cLN7DtPigU7UypYGvcx2L4lmPbn0s3FmeLjfDA/G8Kgf3Du8Cp4pMAdLu
cCdS0HwMeDkqZjmgaC3zQJZllodqy2AUjf0+Iy87g7WZ7w8xqeVCekvRN9Jl
/YDUKRTLp2Fzb539GX9FUbPoLotc05lp6VGpfCHKsEXjc52hV+XNGc4hcOWK
YUz+sSoKAjilhUkeUQhtJG8NNL4dNdDIzAOvoX5SkLqxJxYwdzbHv7X/VVM5
sx0k0BETWdoTZlcrBiqAoaw2PSaGzfGCtgm2vqlqMR2JSMPy9pBNQyQ9nf8b
D4U+rfsYYIXnAo+4h7mDXxaSnMXWa7f9KzkxU6jzCvSRr3Jd5pCGNMCUBAoG
54MC8BvWMbavoMU7UuZ/IgJpSp894IFrmMzVOGI1kXpS4W2u3QqhVeZ08FoJ
qjwjk2L1AWEWTuf+45Q8kVcLO2xn6C1lofRcAlup3BXYdurlKTU7kXyWDVr2
7sj9GXtym/uiHOYV37qMN5/JbeOJTSpAFHxx7j8BuaTI0wPyRMrqR5UZPHQ/
ued08qcEsmvddGhLKXdtwgtw7tXNmomOHXVr6i9x6CTk1g/bzjKkNK6jRY3V
M62JxPMP1TyIgZvDbvNTtlxWi4059z55nw4mCAw75I/8cWpsruihAoO6C4kA
CJ1SUQYUApbycGR1txt2pkYliB5tpGaxZGDoNu0jRTTXdb6wPzIpZ+AnGYkr
Vyyt9yreUIYqISJkqjvlgaVLDH5sXuCq8nHN8L/lGvKQlbjpopM+nsVCiaX4
mVJEETls2yMrbNs+PGpok8gtAX/XyDlvF8vskR3JxaIeWdCVP7OhTRaWgHvk
0v6WEUFNmNJUJEO8nMEPl3gzzrCCdKWBVMwL0DyiguXy3/CqkLd0WtGkh49/
fRZBzposqNuDARpOxD0TfkMrMbxPG2gHSiN0ajr13xi9p19n2PTzoDJ8sOFC
D2Yfw21zvh2tFWFqgam7N0Bb3SdqjqqX3IMO++XyMgDIWFJ0yAODwFy9zJof
F0LcisL9upIh7IbCX82Eef0fbD24vG4qf0OM9d7Ls1YdqIu5l86IGhyBg8Yd
xLojzxBlqHcFgA/LeNnrJR7gVpCpi4XerNEz9i/OdTR9MBUNavell5qnuleq
aerMu7Wf78cwlYXgNGast32C4DEdnbssLgv0bB6h8H56gzO8QeXu/7eTN9lP
D1rMe+Y7FoLKtJFZgIJrbHs7LHiLAymnPWWsHY5b08/vlNXuUe2w3PkeeetV
8M8mQ8dX/KbuH0prYY9VAdEttMT/3c+JCtn4KqdWV2h7g1WwVaSup27vLyhq
k5H+epEEMz2ZqXw3vOsygjtjzJfB7IZ5nWkzU8zenjljWrKk09LuT6WQV5eD
zEqAuKYjHwZC6dPiRruw7KVk9bVKOH0RwIdVYzfn+t+0SFDA8qtUKQd6QAJk
qtzqQ0mOA1HF8W0nHBIPVfd1IQFX/2FA//mgO7b+65jCq2AkrgOSBjsoeX0O
Vh5CKZP9ERdJPuAQDCwx0/ZgpIT5/2zb/kMmLrwXbVH63pDJECZfCl9VZjmC
xtxRnrh6+bk/WBUviNOPKOJcW0DvrZjsNmt/cvMA/jeOTjfkf6I9vUMmzZyS
6v2Py1qdmrRh8Q20AZH3J46h9J369dbFWUb89Vco0DM+Ll7CAT98jyANC3DP
7R+m4CC7ZCQTURtR2CKHDBYXTTAxsa4//aAk2DFjHzA99wzLAqR1wnE6lqoj
1uL2qG72Qo79/D1gHZz2fQ7IBvqntCUaERQ4UUqioUsnX/WF6p5bBk/SpSu+
AJ0FBJlixk9U/lMDkDpjNeJH53fMHT4t0R2WSIAVflASM435EMqEApTgiYNN
t2IFjAQHCgiGVfGvR4bWSGa/zt0lXEL2IBDkb1JuZEZ7YW8SFm3611JwSD5u
pNpsNS1aHhj5gXAQYhuMXnCzu2j6ihScZXAO2QOQ+GHQkFj/tLgFYN/HjeJl
bZhzfgZkat312kAeCQVb5h9TPC7NWMqe7e3yQNHb5qn7GUQ0QjDvhtjLPbyh
vcaEmS48uRK8rxQTu42uAwdaPUI38aL46twEdpesOryZJBcJ1SOURtC8ALDu
LbERx1Sp9KSZZAK7GIvwgSWqzLhC3WwhpHukb+cpZYq59B2HxFbyD7GtZU7l
eynUbfiY73B2GibcIt40xsEmu1QI8fvVqDpsOvpiB1kMhHxT9bRb8x+lbKI1
6XBnhgH66CrWBtAWcfbgoyrrPfv0yneiYOxc9yZpEfj1lgscrZDZmO6Ss3f9
EhKHW8XGJYU3mPQH5v7PSxLuW4Gc+ycjGvcF9PZipTLsxrkUxK4TsCAaE7+M
ZD7x9FjoEAFeSWSgBxSJsaC9gFQ3gsdKlZoRPBdnhL360SQ9y2redzAX7icN
3auL0Ho2q0uNF9gHJJJ5hpILcSa9oLJX4Dh8ytvGCJXHEz2W/facOFE61LBJ
5JZQ2+CPCuE4pLPXdGh0rlyyoWOz/8iZVIq1jzcWBBsgx0AXu2pwyr+EtE/F
4goamUft8aY1XHKOfZpq3JJpuQWthM4KGsatR4iaJ2whMeehIeAESnAfDLax
yKmzONOmdygrG/5mxhQ/qPvjXrfXzWaha8dBYSD+IlIf4s4a4EgvuaMUYRA9
p1KHSwjIIlG2v+nUUF54D208sfkjxrkj2nh7CG4MZcu8s0Rp0mKDeVrYAmcn
ilNV7HR5gdYqNQ56w/qvH9COW791148pdJbxHy97zql1TSgcifTW3slEGhmr
wEdDPmvquPfNbaRZj7g1wv0tvEnZBD+2FLmiP69IYNixWYV19FfXOoTCiqrH
0HNtyF2vyjCJq2iTMnPj6QYIn3+PjC+TpDEavGtQ0tgowWQfMF7klgzsu5JI
L8PvVyQq9bjotnTMXEfx2pKcIKyI29sra0AI8jfKOMOIiKSrH3BAD4Mx6Emt
lRliOjXcXnFxrc/El6/V0AyjBEd/c6tPpaxQqnvJzjlkxTZ6eb8QwjG/yZpD
aMKumfTK2YbyvYxEhs7F3A6U/vehvxOmaMAgS+YRNhNSK/lXtH3smBzD+3m0
2N+QZ4R6Ln72lGqyEv534Yt7fbszo3vJ8sn+PSxFWOvWcOCYpklmLngPWJrk
6qPvPGMN1okN/P0wCKqpEHH8hnbZHTEfBsoC10mFDKWSL+SgSTPRnaqTUPQS
bKjThmd+BM9DaFBfLauf/3nxBxmJH4PxBUJFZa/5QnMplzPsTZa8hHsyUc3Q
6zKtq0Nm+NLMZhOhnZp7QEMytf0rua4D4P9KBwhXrlM3Ak64jmVCM1LzpT1E
ig1XGVb+YtNZxc0jh9BHgOSny4R7hfp0m+/Hx89GvylL0dY3ijLT/OrLSRW7
MZL1AXnOiKUvjDwFJEIU1MQT/QpycVqEEvrxNgCbQC5TP+WbJJf9IQutrbV3
9/utYUMK/c8SJHL3Crj4gROqztem+QJk+3FdHte6h89LyJgDVprin5CVhmO/
Ah47BHq71SsgTjo+5W8mKDvZImXhHs+RbZaW3dfZAJJLucHLak2jeOq85hNM
1SONOfe9WbEmUBBLxJA4VW/B302IiZAnI1MfouKsRdKv2t9eWbh9GxMhEZ+d
pN4EkxaPXsZSvrlXx9FMuClVsa0jXMYtYlEhB9WqPr9DTVszyfhN3OKHys1X
j8mo9lDkY9N74/AK6yHsw913u/BZ5cZZA1rrQC7J8Z4lJVsVN/bN+XofZ97U
Qq9ZfXIxEcU1zz6QpC5CHRCJZ8t7wNf/4OhNH1ODlRkEUdx8bxR1rDEq0lxb
X4/dwkpdUCeBhuU0ojddGrn9Rt03JqR/moEDIvzYtXYaDsBDsyHG6wWf27tw
qII6SWE7uydA0tBdnTtO+WbcBvqTA42RGh2Ae/v45XYqbl1JVwJ37LcQVQb1
7GrJw1s3K1JudTn7IPDq8gvwFY0vpON8pir2QhoBfmh0MnfbuVZb3RlKE9Uh
dXT3RxNHk+iOXb8SV64repiepjd2h1Vj0Q3qW6IfCcf6udYfzSNu+lsn/aL7
n9NtXTuIBZeWfBU6dJ/dv4MSSE32+qMhUoJUzcLJn3GnkfDmuupHY0jINXiz
2ZlhSwbwAhY1f5RN9rcuI2cJRxIOh56nMwZMqqz3qWtfmf11WXrODd5kox3m
K7cmadV/QNqommnIrUkpsAykKu7X0gh2v2ClD21VxAoRfFf3sy4lVfV9avtj
Z2dv75ouucm7V1zweLtitNg86MYjVfMS5jAgbZfb7NrjANzzjyeTjwxBqocn
pMQprhZN9Mdg88Tjth2MQ5+bXMCWuWlCFJMLpdw/qr4GC4ff5Z/+sY2+DDao
qCy+ILBm7gAG3Bti8oIGFX3ZMSXT99gDA5ZC40MyAoW6Zzzolie5VVpY2D0s
Lrcw3+1cSUNg8HnINLpcDVo2gEEDdZHs9uKrnvPlNyJBvnxPQvOuWXargMGx
RmViDZSDv0moRrl2Bd8DmLyviyZg4aIwbkuwwnwkHtcYsndSX6ZdAMqQagcb
dkNocQVQYsm95kZm7gltVEhzmDqKeS5whLf99Kpy3C9mRrZTaJdQdneWT4W5
F3LPe2Cq1kgtYBcOROj9dkp9W3fZCdxEiS3zP235DTEOKgO7Se5c+ErjjjXC
0n5pF6aXDD4TFVnnx5g0QihvHJGSfjZGlY0o5b9IbxaFOYEP6X42KPmhKShH
1V/y4Sf7pV2qBAUPB90cSnuUWnTZh2E6VZPti3NTodPPdZ4/T9WnhsBVRulD
LFxGVKcrdsN5JNepzkci9sgFZxs/l89o9ZahhzPIxEzs9MhFdp9EribaC7kZ
zCR++fdjefy/Jd9JHUU4hDdHVS2J01UKqLRSpRUsRo9XWPtxznjhb+L4MCMV
+C5heeRj/lcMSFIg84VXlXikkKNK44+bWFScv3JRoDFigBlFdwFS5NfTUXgl
+ZzTbIH1dr4xj7NTJwLJVQ+3fnLu/VR+E+caRZDjhp0Fxk10U7eSJyBxOSR/
gffN9eNdAbDxnfW5hqlI8hRVphyFlBNjaU/DqnsNDZQAc9o2rQgzPP4LJgI8
ZgkdA/NRtLvS7nQaukBlYCrCvuK8K/cW4hFZjcIgOgqq296jD9WVbYcK5XHT
WrHmywAWJBb/gvjHoKwQEY3tsQkwTrHQipPkcv5erGbaq7NxR0tvJNT8yoe/
OZK83DjnFFCV8a6XE4Gqwq6b5S+x/7y7nPGisEMhKqXJ7Hnv7z2ioEfh9SCa
wNkpljdD8EF/jGAxBmuLvL+5F1q62sMRbavpsLIW0A69fdU8aL07Z6o+y+wQ
vCch5xJhiHCdKArUnFeEOBAlYHnNSJQKfin7Pu0frI/KUOZQWGOULeaQeZO7
YSLcvwIFJy2QzZyHG1GWhpX/79BKhfe7LkGJof0vUMWl61ngolAUqVTztwlS
3eeF/R/AlxEtPoMTX1CpIyI9D9KZJlaJ6gu0pULx4A3FnC0/FO21rOy2Z9jb
55bwBoIeENstfqte7JeunrIluTsRg57I/9+fHB7V9S59lh+MrVruCic1wtGz
n0TDwKpUkzrvVzVINUdMVk1RQzWxY28ZkPj/y6lhF4sBSfI+JH6HQgpQ9hkl
xc0KLxbmcYVNBiToyA7Oqe5bAx5jCrwPtiZl30uGWtEPLvwwI0JnpH+6G7nG
1dZNIxHHrLkzjvxn40cjn5gtzcwjXfA7Nhly9DmcJ/WNWNwr30qW6WyzZyVU
ukvMvQ0RVByVrr5l3UKhFS5zl+ne/O1DV4m2/TUhOwU44zLmdOT2mGM3kQMT
yAFALpXINBdCeRCJbt1faQzzv94D9BZkuO00jxwytvOaIE+yzgUdl68LspL1
FVY/VW6dL28k8SecaKhasqe2+cNZ7sbtPN/EaNnwHrtAenqdvEpJP+ewBxyw
kdSkB4UbjQRoDffy44ozEz8jDxZlCKUe4j/DnXGrLFpE+fa4bL7sj94PWfIH
4YiTxfORxrZcik+BruWhyzEFHFfn9jTIGBpP4T6sDJJcEN1RjgD5jURN5R/D
P3Z5G9LDZiFn1DnlII+Rhnx2z6853jjuTpnOwBOcWTGecgaocCYWaGnqM/fW
0kNIymL1mLO4suG7PxloO3LaBdmEz33nUmv3GlrElVcqa/iTslFDCMHYqFRj
w6E0oPQiR0s/gvMo68aG6lkiFdlZOgVn/p+mCwoLZuimMFfRdr5AEFOI777K
hD2+SwWIUl/LihKtccp1a7GQXq8SkSIEHGDnGFMWfKt0BKHP7ZwJhTqyKy0T
he3FufP26bzuzHGMr4bF5Ty2Tpy8gajZJNFzqBJ4WfEGwO4PKoxuVNSO1hQ1
fjzFGrcVKjlXWKxyLD+8x0RMdoUenpK09QElRcmAv8marZJCV2/0nsExOyGY
EmG4gnB0MdSPqkIXuWDkVV3CuDr5hRw30T49OFBBbMPTL5S+XJiVNYAfaz2y
Ha58XVScVDWdruVB7XtbsGT+EifWH0E3Gd0oHNOZuIcdvAPLGUw/VlMykE94
zCOTgKiQuIg2/zhUlphbM0n5rd8F1CXtzF6UU7smR9tr/sm9F+jbKCXdeSoA
jERbvbO5sPCLViXqAjfHaFz2XwY13lS4ZISNlhW/DJ/NSo+07dTGfSMu/lM3
k4f5KJ1KppdcWCKYIQEyjRQ87/ud14J74/vAS0aoDLP49bUU8xi/xZpbMGuY
nBxi2e4JjCakkhk+FgAlooj9etBFb9ZpXzF1QsrMNnOM/LiRny5NSJL8UtzB
DV3fRBzaZJbKvwN6YWsq6kfvfjQV1wmzT1f/Q9Jg3JYZVh/VVS/YLgU7hlQW
DYK8m45aIaQAcWb4xzjcDLFKEPApaeTIFTcdz+/Hx2JaGXBZ+/qS+eo0xM1j
ZjkjvIT7PoWUodx4uyWfwNOHyKFOmG6TsWGolXV+yinlRWiynS7eXslrOEfi
YF/IlsoimsiXRTspJ7mIjv/2zB5QVcFsHz+Qhlrz/EYCWaPzqF6rKT8H/zWq
u0JnhQS2FbPVyKke6SemSCmGvWm4+VVyyOZXuDTtffEDi3DhV60j+soh+nSg
rY/qMyQQVLHXmJ9U8jcyALL/1WfXrc5lDNz4T9DXc/nJ01JtvO9wd9ZmFrm/
5cI6mxaUeMfZ2kOPk/W/X21etmvId+d5xc5Tv9LzL/2wSixN+I7RfdrypHzI
H1E7AuFYpo5+SmNO0nwYJ0egCaF5NHBb8Zks5WLSf4spPBc77ksi2QGpnfGC
6MlezP5ofOJcfHH6SAoVgbh+JWNQ/PjIZC/D03dzm1o9mSI0it8acG2th8JB
WeeIWMi+qMu5QtA6WQQu9c9aTVPcqbB5aprn/W+woMVUVGxkwS/4EgZ7BXbr
hw428952Cspo3DRQKOdNeXJ9x8QxfaiSxLB7iqcmrJ5xDhP6gizQB35hwVjM
OOwEjPNveED5DfgjUTSbevwSZWO19CVGJIlF4jFK9Jbpwbvz7bfU19RjYXek
21Quk+TZiKSt82x6PEG/M7ASp0K9dZGjz0wCiHBHyjR6m59/e6TIkdCDvcy8
5/QbYNoNgLVcFCjIoDnNuDPIGNSzQV17iR6nSrHKmK//i4WOSVLid6UEpjUG
VXYOqYuU/FTScXzoJtrKxGdkbakLIcaSNVa1wUVXHJYUlDj58Tkd+DOQuT9I
h5OW50aeLcd/iCiy/0CWAmjRida5avq4UayVzNKetZeUwqQj+A3V2VwNfGFY
ggzjvwwm/K43JbsPFWGZr3uKgxw1buwmb5X8kDL8Udi1gGTh/Yp2dvGrAwPs
VKt50XsEjIxLGJ2VSWCWoB3A8E8fGMVXEqbSYODKdDlLFnJg3dIeux0Ai1wJ
QwUB6WpBqt9DFADLgp7JPyTMq2EjS1NCNUWrCHm17TLcrwYTJzaeljSWrEmZ
NZBFHVsluuTAyHIGjfRAkcmJ6XTA8JUBiETNCHKCebT8CJ+2auPEGkykOFKr
mMwLXv4AkFVnzJD9/zSKo5b+8+vIKAkLq+ATz+uKnpBMFzo37nJAoUN1AlFG
0vROKCOtLhMIfP6vKEayzNGnveQ0LBjDwocJwpGKFBE4Sup4wYbIi70kGj3J
EwSa3HlLddF1m1D/3BOBf2n1Zp12OLdCuA6MdXdMl+L6P2gL1TEYcUK2Gp9J
jDJnhVDgilmf72yuKDq8XrBbpK65ZpnkrtwHP0qraUiUI/4JZ5Q1/UdSbpAM
CetArjOSCjpxWo4PNSXDHMFQ31PrSzxrNHEb+6i3JjrZCfPuigOI+4xnfiC9
9CoFIIlwzsPQRchUpmNjfwbBEwQzFMp0hC1hWRgNAY6BgaIdz8KeZFZ6bOhs
vufvj9CTr6e0jnyfm0or6TZz5laf+BJ5FZrt1tahaRSHmLvm/mYOzQ8IFhEy
To30U/JRMWaV1uT9KKxZKdxTqrU5R/Jnx8D+KqF2TyG2zK4aqKEnCKiatlVU
x5WmpPzPKe2nLqz1Dr78dCM3u1++ExWMX5bO7ZqKWvv29xyxbygd5r6ANkuW
Gw8FHycHNTAKVdQs7YvYslnKKwzhG/z7ISkg8na8nIwuOh+6/TR7q2NbVO2P
xtVhMHd+xNARMbNNE9eU2DxSv0NUd7n+hMpfDc6Y9+pSi5zK77yd1WLo/36r
A4UWCuZ4GXxk00NxKRj0TaxKsqirrX875xJHp5CbPZnGT0qtX1HRY8V9Fg9i
XdKavU2wlGQi0CgpKM4F1+JTiT/D6OHm/pNIwdDAnpqXeomi4k3T3WYZLGc/
w9wS5fvw1kgy+g2vcxVuJfvZG70lpGjH/2U3H6wL8fGWbRU7NXNm1FqTdN/t
lVHUkMz/ybmMsUjp482sTPToEJKNKLUIRRQddNNi97iYNxvD2Xjs8O6RSAni
rFhVuq+3/Es0Nw7FGK0ZJ5Y5EOSsPxdkSszwv6Z6IX2ZSjlYwBUzdbOw5xsX
WR3uy5yoRWLinoxJ08BqlUegx4sXrgG9Kw6mgV3XRqgLO9HwKK1E8nRgVfmN
MAt/7yZNcL13n8Hed37MS4IXatm2E7Xpwyy9s4jYdBjsi0l0O/baC3LgQdZr
3feJyONEjWJHIngWtsk3J8iUC/I2E1V6qrg+Ya7jgx8Gninhnm79u0Fx43B5
ROMCJG/gyUTPbNXcrpfyulMxnUK9d7jR3prpAR384NpKMer+aBxDyQm0E1NE
KTadh26FJ7+SG+uYxYkWGP2JEvFqzkbF7A7YSqkrc/qWqvlhnVo7/WaBc0LB
FbxJ245evOonGomeboZ9mIL5QmZL/ALV66Qlgffv50TkkNYCLiIzrSvqZgfZ
8hqGtKaLQruxRfe6Dk8V2dRbsqugvUQa06/v1viv5XYkNiYF/U24qdtSBps6
uBA9WfIoO5f/R2Nip65n66/6bUCRCo9k/P0tf5D+QS14knkUPiymTQpf5S+F
624kwA2eVbkgF87Pxe5QJPlIWx9/wRf6nPBu0ZiFSutbVmssm/kFrvgtBxRg
sSKLwffiTvIWMDC+R8QjprhI7y4SZxVKBtwcTp4cj4FEmuflS6icbWMvJ6Q7
HMkJOaTRX1SHRS/mEFhwyaFetWPOgok6zf9ddSmSYIx28fd+JSWYvWwpUDM0
Y5vEbkJGX1bBqJx882GWwwlTAUVKaPtLzm2AS8WKrcjOqgtD1Ki5JdeF01RO
xUo9PQlXcbdm0q8rEWJzjqR3rfUPYOg2C2nQnGHX3l4htyKFd7yaEP3p7gKi
8to9hNRfY3+N4S4GhbDIS40mIinedYqR3aiB5YKora2P2whYoQlCTpq+PPV/
GMqhHI7NW+maEtaf6TtUpDkFjN7cOcMJUMpyxAC7N+RxFNaUcgFVPNcvgIyV
d/kRpjzhUsVyfOXjjtkwS3f1VN1MIeko5dQZ76DcuRgbf4YXpYBdie0GWAJe
TPbjgQw7QkOXcD++ZuzX0s5GkXhLNg0Uzh1ax558hzw9OnIYn5VYs6eB2nKF
ZwGAwfBPC/asw82QyNKyeUx+xfi0SzYK0JgFOksWzUSHydU06dYvstasGrht
KaUhfP14WPP/oTAExuA8o1jX0I5jGg6ej0CwOFlWo2xtaUriasS3hVyec+lG
h96esBmuH5BS1HJ3Ik/sdk40jeuEbmL3c8UGHRgv/ubniJLh/TdTbpJlEEAU
MhO7/ufz3G7u3yMcAJ3b12iB61WH+FWqcb/dd3ZanuMyKSflFCQDXiN4kJYt
SPJrVaKmfDp9EEwR6rX9RnSiUzh4PTbr5qqE54u+yCkW8bwHR80MkZNgVyxC
80HbRmXO1sBO9WgcKL8h4UUPfegKs50vxThkto0ZWUoXMnj+S4AR+k+Sz6mU
9/QOLNnmfwWwiHmaIoZ3fUuvpOM+M6bWVW3exrKzCg9wk5EwMcRDM1zfui6S
7KhuQqgvuJr5h+ZLKnZcZzEtxH3tWlr4wZ04pyWIr5eVvD4350vIA3pBNquY
Wgl/oStpeTGsjXss0E4A1YfAmuvq/Rv8Aft0gFm7ugq98Q7as/bF+8Kcjv/Q
p2Zdsivugi4GnDMiIYZRVjPSXRweitQugTsad+nNxhH842L2/Z2X1BhsYeWF
OWNzj6P9nrdW8Mhv+sv40DiLJ46fSp7sx4ykdazOvsVhrsSMImPviA/Lk1N9
t+ddoMoLNvuxa02sStFUL56zG3t/mx06cMMMnSa1zeG41RCUfZNY4cgG6SdS
neAW56Pe9CwTFZVVgrNZ2gtkxspCr8LLyTda1Cbls3QVSwiIYYrBQPTCAwYY
8MF57zvX93viLf0POSbwJz5wIIFL0bbw60FvEYWHsrq3hdhp1nYTVm6GOTuk
hOvNhgThvMJHhRFKmVJ4d2e6R3gNUdCws5kO2/3Jb6xjRggUEJ/SfL5XCt15
vZanzLLuSvR8Aoyi9IOIJr+27Iar/t0v3SUrKUuUt3CM+pjflNcm7sRIfoOs
T32TxkbEWmuSyQzC93kAHvZIkTR7qzy7VZDOnWXjJ+NS1WF1Q3LNlX9WWFwK
HgICvDFGtmbXuO42+lJKbhsYiTCTsQGCXGok2r7/jssEz7u3h7y3lzmsNq/t
8ECzI/tyD9tid5O4rJ6QAOZNKM91KEO5+jldUdCKmOrM6Hp/X8QBqwvH4VVV
ge/SmyWLosRmbKCZDnkVqrZecsPVRyyKhOKCwz1IB5R/N1IRtp89nDOzTbEu
dk2OHrqDWIj6X8K7ghkCOSRarIZmldAhACJJDd7Z+nWW/S2ouvzK5Rqiw0ox
+6lWaLTJ0WF41BrOBq+RGOsMKXHTDBasq9ShpcHufJdtU55BWgjXzUFQ/MPL
me2aBr1RN96O4qdJtCsRF6vLRtcIgaiqVwMaq05eiGFkXHDkYYRrVdQKZYCS
qnvyjil0ANzUGMjPXk9/rFTN+YaJ3h3zI5JdPQp8v43tysE+y3wdTeR5yC8H
fGBVShzm9nc77dy97EoVRjYyNUepwj/I3U+Ssn0sWF/th/XHbvfY//nORL9H
t3qARPXzTlE+9wk5LUKucHC8x0vlw+FwhLPR/U0Twfu80j8pdz+QmS7bL0H6
EoLq5U5Jo9erj3PIAYJlBQJ8URIkgjHQ9JrxTC9ty4jiTjpfyqhSfr28oMO9
GmrBVXKul+aQPvq6Af1tBl1AN0+DQQcQbIoxVvzgKVIXJ+++tei8OWDVQYLi
J/VM6zBorO6w6lftc5wGHB9i8VULZ4bS33FlwtLwQ90xokn32bp9p/paQvn2
nZBPy+y4mMA2lJQ7Drjb7t7hBYq3LG704wpjz62gurSCb6/VoClO4NbblinT
dRnauSM3t/uXecaR7301WDHZQ4Ju8t/o2S+22x7+5JlWibdSwBRJo/IrtQxT
a/Q6t+YZSrxI0FFG2ZU22wckGHM+SbSnzfEn52PYAXKHs9J1CkuqTcGFhI2s
1WnBRlsOQvkIJZEo+mMDkusdsIxcLZGOK7CGyvZfd1oVCoGja6egPLrS6oMt
zR7ejrSpOQIcbceAmEUF0Xf6mmvlnNiOLKbtSiphrjY8tDwDRnYJ5Fviw/2Q
arEDoKVej9WyqVsgTpCbZM93ktSHLuDRY4g5iPp3dzp/8bFcn7iJ0GvqHZXd
7xbmePnW7FWSZ1mfP5WW23ivDwh1QNtEHKd/RWtiNOapHpnqHXd+cnm5iPUm
3l/RtsH3bOJjW6GeEjs2iT04MmCJunM1S/zieIXuB8U0i2sww+uwavt0dcjm
arqDZFnru5Q1THRhqbwhbWdz7EuRdPYQLvYhi3gy4y3P1LxwlbfKJzjAT6ZH
8iUuHc1GXcbWJilQpmUkpdHqgINEGtrFB/bjx1uGkFtBiLVwCnmmH/XdZepQ
diWtHdWRzeVVha/ypt2luthD64RNie8xuAlGlnES8MBtKIaNa7XSEdPMhqic
5ibQUQPM448SkSO89HfdqGxjQACy48BFHO188bnicwiPoZPTRHFEWbxW+EQn
os+/BHIvZT+TdfCBX4mYk7u4ItrK++iFycufLyXVIg96u5764J2p+2dxEtaz
yI8tdz697pNkUeOpG4Owp1PGbct4scAK8fovLE22ogr9f8DzS+ftweczZZuk
HRuN8eMZxLwbUfxlqBRcMkIGNDEQymU0SvIftTkkJBr7uhlVwwojotmWg0UF
LJg3pdknuP7VR0cDIuPtM7MYEESAHFh5/circYaHZWstZDtdyYP0aUf7c9pr
hyYclW78jwytSDQpC+81TpEu4woUXz12n5tSct0nQXtR2Reuld9qjfKRsLet
cT0PyFhSUT5GbFiPYk4PPNV6ji8o66mhC68MUCtbQcV3jlcgMGvzRcrFPvz4
lUlMZQiWDBdjOpWq9Dy5f8uOQ7WYg+lJrUN95nYutdAfLKslprPTAAFC5Vn6
iaPY39A4a//W7rQMnC3qX64UXNHHklZxwbnDojMkuau8H9zBYDS1xZXzgocy
u2fW3FijGbHImqELnQEX0JTux79bVws99r8cVfJQW4Ozm6xNTOmeslOObQ/V
Q9TzVgZJontr1uSggGcvP0ElsPSQVTYcswhvuKdLGKU4uebHdw8cJj6HOptz
aHOG15nP+ksNiUtlr+1a27eRqZqoRGYyuTX+2iqEV6ovN+erpfy0oyDnemk/
T8WHvQXGMtxjwbiMv10wj8P3991JdJGQKMZhnKMvgvzG7MhAfm2BFaKm94Wh
sljgZ6rhQvUAMmAlYow3l14MhB/avFOOUHiBeyaxhYf4cCbkDRYAADiPL9SZ
v/xxREKmm1sgReTE3O/iMpVrV68l2+An1437/NmcGtCVob+GHCM1ZCbk5pFO
6BkLT9q9bTeHQuHeHU3t4JYoQ/aQgd4hFKiLbp5Ezvyfw5wk7K2aCDo0+AOS
Ukl/fLb6lF9eNy6sAbM6VZBrSJ5NKMicldA7MQHaJ61iSsMi1JZFtIJ7khoK
pBeC9I1fkQGkQWKXKRkwN8x0gP0SfrGf8qENjcUOgfIU5K3n/FUtHee4XeIm
Extd0Bu3OPptNBKPXa14zN8Nk1fIu4WRLSfUORJC0QqfAlX4qpgz6p43pc4j
hTqCwohxy50E0O2nT/GadeU5zQBoBE7GdsooUboFXLXDWsYI+SOU8nzldwBi
4iLEWwY4hxHmuPRWkYHq4OkZwWP4jj1hSwGriXxiYP6/fdKC+w0OzF3GMy8t
d5pbGF+GVI3723BJw1nwb0z5bxPbClFvLk0S9QOk5B9HgcEfV2Rj6gmn+3Px
Nf5hRYI0LOSGuX54ukR0R5U5ZkhAn8oRuRcKvAKs5+ho62CaTbsgaVw59F0h
BmzZ449Ff/S9JWZCqvZ+9qRlABZu/8iHycMIRX9ko8aVr2pHwgTgf8jQ5qGp
rUhIshtTkU3alq6qQlMKMY3f3LwAZXH3OR+IG7z52BzpO26YH1bxcyLcEdWL
GNt9dcmDjOhJXpHyChuIlYB99d+gvU19aHEfI+7s8mObjRuTnfGBvm5bN5Zb
KddIp1eykLzr9b5zCkDhwlOnSCr7+JWp7mkNcH/bjT8uW0aXkc5p4RWTW+Oe
Q/OtmqFORp0MO1PhsFIjf4KSeZL9pNa9xZIO6JbywyX4OH8bhsPTB0ypdYPH
mtSvWOM3+Sp6Cafz8QsqrRcuN4daRhbbXYevxQR3LroMgZH2+nVqLFqcB/SC
iuAwQIkEeqMMsnOV7fmUl5fcPK70dUnFBLs4a/5VEMctW+CEMpm0kQSwTZg5
Tm9yjnG5pwT0jDFQO+rejOqZN6yyejDH1bAMXqx4X7GzuIlyWSabfScCPM8J
c/zAbtkr/gNUYFHlNw7SDOYsS7cGtdBdbtKlz6ykS7x7wkLAZFE994RlFtl0
4zHCYPMbu45+2EkzVJPNTD0icEHVQuKTq3jV/cW/M64X1Rd+7O/s7ebYCeed
YeZJI5t4926GHgsuTlfU3LBp8kjbnH4rbSO/L6fwxlTqudSr0wcQkFgE5X86
crk2wfin103qrlpHuToS6xKsCLA+Sd5tB95z8K3bjziFbuZfTsS71fiUbmw0
xS+Xae/12h9EPmgadG6OtUtJ7AnZ99ijHO/7MJ/MYIhphNzLVkwjO0UtJQta
WSOWFZDP9KLWlAHP7y05hrlxdwfao26FdTWUxbuNGUv0avDd4aR3HDQLcB1C
BGvrfC/vE6HwaRZNT8DHDqBtbSZeRwnhMWlW4oafZtiz7j9nUE27SJtUCagH
iAOAf8tYFrtOE4vppHzS0C+mxdrkIWeVORvZCNfyjdusu+jshU9DKE/eJjv2
A5NQXdlzTIY6kT7hsmFIFtKkkH2UYOABRrhj+9HZLhCcz0LLFKMEkuOmv5Z9
hBIH933YKhHF5T3oQYL2o6kyqCWZL4XttiYoMEPXnDmkUxJqjuvU4ihr0PYS
yqkHwdJCg0gBRHxbt0REg137hy4a4uDdxLP2yDedCCv+AIoFgk8ea07C+ANV
/pfUWcx9I9WAdwToshBDbfo3+yCH5kqxgV5e0aAIxVumRgV+pulb1EfuF23V
RHh5mhjrWqNGzLVo+6x42SAs2jJ+5UFthy/Jj2NvZTUhX+kak57QN7cGmq/6
2l54fEgcxlu9HDZVvPjS6ed2eBEJCTO2jDuHQAOQfPG5IAkL7O/6fd+nwvfW
KR63OeWIPt5nt61KOtR64Si6wcWfGkPL6xLaZE+ZVcOcaasaWri0JtY2NZ15
zR5E6j0o+awhxq1K5IjQNm4MbGxaRuXbSKXgInnpNFJBj4ZxonkR2B52/qgB
y5N4Jhjlo4plSChyUzq9EIIPKTDdhPmZIgZ/n0r+ECKP9AcExHh2+/V/lbdT
HowuJWEMNYrfbsZfGLAXTBj3Er7zi/y/mXWMoI0hmTr/ot5f1HqoHHfxXMyy
NuFzGuV4984Rjs77qDRbCSpWFZFF9/5ip7vlDV3JoJBSWsIhBeTmlX2ty6eT
BEdpCup1QP4x2S3o1mWh/UhSFWtwKyGtsoBvjuUwYduDQgy3cfaHxcSm1QEQ
+iK6iwsd7MNS5doYKOc5q3wVN7Axri6PzzXKrFJd1fMmtsdGd2ePZnTfx2CD
Rys6DZDWZ6Rb7RCx9wjpHkZnp0Aqt5ThcQa4u9jK81cxGJymNzrhUiatw9Hk
MXPeEz82P8lYtKmAu3tpoTcqjPvFQNcG1qsd6NRxpw3BdLSpAY8YvLHdE8Ac
yyUddtAsm6Q8FqKm1OdgONElvIKyWBaqc1RwVcGN0kHEiH+1BIXah4Q88Yzp
eFwwJvZhCgz9pfcrGwCKKtRDry5Z943XTZZYCeOLDcCwuaF+70BXeM6AO79y
cXe6f9huMqInSn8lXraD88Okfct4fcUA/O9MRVCmInmysD08k8cGtT6ZwMiY
ke9QCXmytpebe1aIAzOwG4+t8mfrGQ0+XW3rDXQFtt2qtok9bi+vJw4o06wK
L1Lu/js1ohMiOzjI1Z+SRvkQSs3GD9U+UVELnXxLWybXudaOYbjN9zHUm+8u
NWEdnCA55jxFGqh+ITWYxRI+iLZF/A7dMjYY1+LfL0aenkbmrBdAtspsSKVc
PIaajXdQ0n5vTcLvHae3fbHq1gERBexkLkCPpLmE68BXVzWxKv57bY2gbWsT
fzyTQ3s3Au9nWEE9jUgcWfNppZB27LKiTo/ENMA3k52iloHKVqxAVTR/4XvQ
mNBnD40Xw7cEfMUU6Eh4XJzLT2G77NBXEAvhiOhXrqDA4q4qMHOkOlQdFjVs
S4AhCco27sQWN2g+Ee3dUQHl180GGmFI7Itqq3gtyBDDl4pdfvGeAdnbh8g/
QkVkk0jkLebVzNDX9IRJdWNzP3cT51AqWFljBmHm+4XZGQRDGABbaaY/JHCA
nAW/D289yoomPEmhw6M9mOWPsvQDMxuo1IR79gcCY7jaBAbhZo7UNObFPUw1
QpHOral+8AY3gmiM8vTe+nL958ORomC7LgmArW/ErxvjuryctRe17KKrLsmr
2bbV4uPfirHZNA71vwNlgKZ2kiKlstnd5WBaMEnlzx3nL5M8C8uvOiAyhcl3
lhMf2V7shtBNq7J52O+odHkBMj/24wIUg7aayj5xAsVijTJF60pUw+bCQyTN
NDi69BuXeUXGeG8kb/lxH/WuN2BFq7NDltKRvTjqrAA2Joa4rwqLAAI9VLkE
EJlMSnwMO3xabBM78tujxrIW+JDFlF+113KB2Ry8CvcZdOHW0CBcV1yyQzsU
nrMR4SPiF+3aoXS6o7dP5A3fMN10rJZY8lnESe5uktWz6DTjGhTU90/MAjYS
CY9rWIrMggM1ZTYb41utWCDDSYpGtftXd5Ig0xmC2vvrmRFGn5cyh0nzSDH7
t5BPQipjGSqs2yJCVA8koUelN3w4HE+87xHAqK9Z3AF2jA8dsiQuDbcS07n5
xwltCllx5N2CidrfD5w4HxTjEXWwemIs2B78zODuqqYdLU+naLTGJAfovk3i
L+2tu6uI0Dnu9vcOjpCtxOfH0mHtPhqljAeKywGt0bWzXGVQam7hT6Iu3Qdj
zQnWVpDl1eOxZ2AootFFzm29s00DZ4KmjAClxuMSxpdQrfE1qANCGB+eRLfU
2s7ztTBhUzoCRaQzXG02HZ5zJHvCJpQYYRg2FYkizuP6A8Pa4tcg0e4NG0fN
SC8eouq5VRBnS0qMLifhi7wynF2N0Z79Ean2OMff3B600tCFyYOMS1RshL/k
A/AaGcZd9eLMxnrsUfepVc9tHsddkyfeTUP4FemreR/nrcjrYvq9z8epGXIx
5GAi/xDhz2Z99eyXbyiWdYGdHols8Qdo/L6BpOYO1CusKCO/0SGCIYn5BzKx
e2/3xXm2BdfPXJGXZOTePGzluUfps4mSFXim/AP/98dlpYhB6npy2eI3CBhX
38Nnk32JqCe3yaJCLAhuFWETOBOxKDMaSQGoWw1ZWXKywH3pWQAlRZoRxOFM
t7eNNP7r65DaDcxMNOTK7iOBtOzhvgA2SpS01gjD0OIDUrXNYmwB8QSb01KP
wReBL/aHVueVEVzn/l8QQjV1CLTTV3p6zatQ1miII670JJURQHr7ZENq9Zo9
fRzo8TYDHGJWyxkAPw/PRjDOTF2+nZQsuV9b4ymJHH7tu+0mh2O4+9gXqsJu
P2F++quY49qGAqRoW2AO4LwS/IbfgYHMDC30KdbuBByDXmf4DwbpFWF9LD7E
ZQZF59F1U/F7xMqC/lwNgZ72fF4jEhWqarW7wDY4g/LvZlwe+taQrY6EqoeH
At1lf7/SvAID+QHSV1jvkmsONLZkhDt/6b9PU/ghwL37mXAgYID0YM7OTsvP
a7ydytcYXvI6V44Xz4YpZRvPPudfPEIlxfiYbcWQVBwbtt2pmhUF5Yoy9S2S
zqfuG9C1uGAbu7SCicAwYQpn/kgl3D3OclYdHe+vIOVFxFKkGWby/kpSEcCK
X6rl5PmJfeIlfCFn1d/fGn8TY0AxFCzo43sq5CRzI7NVvn5qsbhjIbqLgapn
09QBfgSar0H46Nzlpxf1ihEpXqgZ7QwSr2OngF89jVch192SdMf7Iq201inP
TrBocV9g2rQAMUPJsayuD0MKnSr0vbd/HpD/7he/y2oylEbh8Bk4O3xC8v4/
2yJm5f/7Zxm+J3UZxnRebczqrA8ixSvOdzBGpIJnAGKvwrPQD85D/uaACNsh
IIMIgLj5cg6zMzriH76lL5NO9mPAJk5HZlpG4xzRbA5REDWwn36KJ1AgNCLs
pZqJQDqeCIMCfqbprkibG/BndJsMWHvk70kbUIuAZuf4C7Ai5sn0RqNKRW9w
U8Bv08HwuBL7SacRKLDr/jm/tkfdu1mznYvB7SMJEc7TV4LEHdIYVHpLgA5w
ZXeeMWFkC0Y4HkH/gQdG1W9wihxgHfMUXhr2KpRAh6f7DwiUZT3q5dBS6XlO
pxSXTIf076bklLNfyNUaS8pvDldUMuNmD1A1lfuf9vqubqNXI+q6WJbzYWSP
M4WOyiqwxKognBoqBJ5yguGJ5I3FtzkKY1GZWNxHyoRMaI/r0sS5knPcus1q
YeGz6R5xh02FvgP+uP/TsV1BWy//3AiERjlLPl8SylGrRgnRc0DAHEjxAgYu
3mYWeM9eRptNF5zHwextSjmmLAck49GVBFTRTyOeAaq2QpHNoPSwTB+WwH17
HM8cbudUvXhIDRhdRCY1897dH9MDcGsHZzWih3cwMv/a3yOXhm4KAMUTTr2e
aihUVpeDm3P6cPMG9Kcvrnag1t7z4zRSxbieH/ZwMLioiZgFdFld1tgQOJYx
7QFk8+2t73kfDjNEs2dPDBtBdu0pc3Up7OLXbfba/or0GcWqxcaHfKRr+8MA
NMR0dfFAJ5G1+No3OBTL+Wspqq1bfUgHh38gDfQaloF5NbJQWnodXUK6TnpM
iVIRk+v/HBn6zL24qspNSPxXMJcEO6A1uCSNsFSEDhEHAEVeBk9e/VnTYm7/
idiaTnydDF4PfzUUeGQlxtcIYW89yew4ky0Dck7w8z+3AJ4DrWtmfgnlfo5Y
0L9U2xT4pyUM7f4PDbpYRHiXwGQsKONlde8FjBAb8ziJ2nVPjxogb/RxTZ4c
LrB5MAWtSIqxyLKaaSMAamr7WJfD/afHLzeoHY8j1sLOI8c+CYuk248zrmTD
hCjsAZ6Xyq72GymlvGBt5SnP8Xlv/b1sXoP1nSF1kDD2SKhbJ7WrJz+VabG2
MGbq7kd9TZ2p9uGHZ1/8r+hIVvmkuVzwVN2sCXBQ32XkdhEZguhEePeNEFaX
N6vKytwwB5h/DpfQVRF6DtlhTDiIh7verhcO2upTf3GMWLE9iI0yQs6iQrAU
16eFJ3Ert+tah9m13O9D1Yirc+H6DrX9aSLTwqcnMdm2hha3eRfXIvO/GYnR
0P/ZIjpQUa5bad+mzAWk/gV+rpNVT7JmqWnz1ZXlpv1mBORI1rIG2wdGRpiH
vc7zEiVPSMv0l35dbRmpW2jd3jcmrwx2FoWn65cUc5vfvrm5/7hkiqRk4nE4
suMhlbGoqwCDaGZkWFyJZ55+ukSR/1X3JhR1HzbO9YYwpaBJM4BilPAoDLWp
jRp8cM+gQjKRxlW+0QqMj2yKNyllbGF07LpywiXvTMlKqKNz5UMqRSjFszsi
6cpN20AMgX2lK118qMO0p/MjG+6ESLP+4xFxXpGq/jP2wVsmKxEUF11VJxEy
Z3DbT1BJ765XLBr0PQvWr3WDpRF28lExnMLdA7iYyTCg/ZltY4Bxf/sK6B1C
R6i6RS0t8x7jyMePGphnU/N1H7Wymupte9f6UAEHN9/SjPTJn7IuXAwRvJDf
+FSdaWXS4hl3I9FFpP7aBZcqjKzCU78CvhkQmvslWBE2m8CRWvYEotWN3poJ
6PERPU/6mSMusvkbn2t2RBSw2M/yf0EJElGNjF5qVRs9KfyjTKl2RrlmQ8Di
kctryr0dfm61Zu6g3ST7NFcGA+6k84iCSNPFaf3acY3klRMH/YlDjiWYvupb
EtFTWRzdv7z5EWiU5c3rs3T9u+X4Us4TzSlGP8ujq2ZgmNC20f4LxM44FkFI
8ecgfhZ0QkMnF/HzxP7W7U80xOeXrdRhUlQLvJ2tawjcoE/Vdg6DSk+mZxIf
llxhaOPJWM71iFvZzKAoEqNrjPrtWRSuTarNBdZyWfjdEafDn/4ONllzLndG
5wNNY2ZbGdg1ab8vl5shdSmhGVq+PFgobw+suEU4JS+scbyJk3MTOD92QtXm
dJG4Zyd4c0ZrfDrSuUeNX7B5+V0SceyJkq1c54vBkxGyzfJcmjIz/5QRI0ix
OzwQb4K812dJ+p0D2b7MqEe02sZSOU2pQV3FuHD9FiEnq6C+ze981vwVEIRt
omCfDoeqTJKkGeX7dlodsJXor4kjI7ur5tgD7OUX96Imo4+/LE8aBkzQ7INq
C8/VxvG17AV3V56rFBCI0zCymEiF84pj4naQgKI/C/+/EK9DvDI+zyQZapBP
wH7TapqWW4oCI6BOwAJt4wkfj/iI6wjbvdkb9RqL6EfynkYBOHrc1U0jJfdh
8hipJz1BfATR/iOWw/UqRovnsGSojsTXHn3x3DSqC6qC9k0U25x+TAg45iQz
StBBAOAkCLxdijwEC2xkFhG8zPkbH7eOPl/vgtGUvEYZbKoL1xS+/g3HT6/T
Qa/XqpCnudBr0WMeLYS5msVgDv1sY4bcLHVu8GxkPssjCejTiOhJgUUaD8oY
xArQ1ECpuYun+ZvC+2YC7TXxR1BuJXmZzvu61oXDZhAxR3tbQ8pFELQOuK1R
ygAFZ2w8JIMICe+LyAUUjUMTxexvTnj5lEawlGQtnC0iqXq9QxaXL24kWMBC
mlk5zYB4mNrmAnHF08yao2+JNf4PG9XW9VJQM5yraR+ImBiDp8ZeT6qyZ8fx
OQYhjssxBPb4w5oUa7W7wnXLLH+A7eZg02tcCcxerl1CzlIMSbJ//oAo9emF
8yyTMltu6CvInt7UHFCyAbv8Pu6THvw11FByZto6eun9iqZJsTFZXfjinKcF
FllZ7+LV5u2fA/YhY74WBpI5DBNyIuxj50JmpOWx4shZL77UmWN2DKDGJ6zi
tsglrWryUnoTBP4ixwBMl7GCC4THbr2gGWcWE5cE1QbVQ1TmTGAF07/a3am4
+dkAdOOLLCvyvxbWbx+BuIXf06xwcUrW84QaRn/ZwV7L5ZF1J0kYjWzOG6BJ
C82hR0WjHnyD8J6hiykxj94DavZPOMqGPBsXF1BrVw8J1VYeVV1Om6xQmamu
KPgmd6Koi2HRyeh7qJYcvKPstVkTWwu0PmzQh7upJcZV0P4mxahBQFujJ89n
hbgP+HOnTXF9sExs3vBe2Aw+lccD2rn4FUlUhtkwDpfO4H+JZ2avMU43B3wh
Erqmwm8n5BHY8+cBMiISBQUj5cZKcQRzmHVvWVg7KhzkHLFBI9ExGG/bpG6u
4KTqUIhx0aUScypYOWHiuJD7Ybdly6gBbjligQW8r3Bgpej74cT/F0nQWlKn
VFKYw8HC/cjPdG/2SmlHkOkcUOwc8q6JxCma03kqYRouhH4G7ZiERYGTlSHi
ls76GVz+vhb/nDS/9kzmlY80POmpnQh6SjS6rHgzFvOzYtHR2YSoj950ROJM
oMopqaTonTzkSm7dayjP8ur2jYbPzZKVWwb/IfawxS4pUY4z0H7CVnPjMP6g
SwzW7fxNrB/GxMcvryygS83BHp6dJ9LI8ZH9He4PQrJ1/v6UsFwZ6wGkfnLn
MPNhgjxEo2HC813X+Rhu9MbAjDSYrpQvHoi9hbFFkviMgqApO0DL3Y19AKcQ
OhSNRR2Nr+rdWanQoxbCz41Ee9eWUg1HccxQoJ+InmBYlYfLsGS3yCZ6f7d3
XiIhFiJMliJZkIM+oDGi4QRfnddC9q6R4TWk2raR/H0oM+w3Em1Xi7cSQEYU
ygkzgLq7BExnsCVB1Ira5Jl6Rbre0IZiHX9v+nsCov/Gt4Ack9CkidyA5lt9
eqk3jjHfkTskGCDTtNZ3SxOkWaUkzshGAY/OnN505RLrpqfIhtYKCcgXsCST
mnYvOnoeJrazU5cwzPf3TQitGJ6RANWeZzjriU1Syoyjw9kHAyyNDzC5Si4a
A3fDxXDXwQyASEw11NJ/itD3O/aJ96Penhctu68buhoAU+ubQQCMx1uS8jMR
6CSjF/l4aYJu1nQsBq4MH9lZ7RdynjA1BLMcNmGZh37wgiwkWg8SgHOc8VGX
cE2iteJrww48RVtXlWJ2JzsVUwuu/nTy70wOdMu2t6tvth0jKwnMv4m3pVUl
CsZcJ3hzAY1l6OuP/n/2hXKT/me5P8jf4DLB2uSazJP8lCs8VGn8P1Webnus
blbxkWGzoUnZg3FFaEs02yachYh1jlXSDrY3nijOe5j9zcH4nxN1j0vYHeZo
5RPy/zv2HPvyM0C9ZBbQsC7XZivQeDN5UoSGjhYE+B+MdLrb4SvM/vkk4bpZ
jiiDpptp9z/K/WaA

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "yaY7fTVF6k4Rtianf8DVUAtk7LLjwgb2LeGkSIY3RRnpf21DVI9tSyTJ6QspuU3UyB72ydnkhVhYU9ymDaPK8JFs47feqoSvWsGdNY2pMwlsIUHf5K2ml+QYbJMDDkjbDV+LbZsIBCHwzYU28ISwleUnMnNHYFQfv64JlmYCmnlRoX7xxKJjXhmboPQZRacCw7xR1isFiRsXGHfMl3v7A81l2rNEzQbeI1c6FUAWH1J7dB3y/4dHgvE3iqrIYSXPzkJ1Ox5QKcFT5i9mjSzbzpc8vNPsMwH+Ki8+Xnt//CLCQdj4H47O5nKMvrnbqdEhK8uDILkLwyarHymsBaNSFeKQQSj9Z2LgAqkJgRzJwjai5H9sRfzf5KFxyP/UrNo5u/6KhCbqAdP4EvWO98iv5+w9CNHkLWXt07kM9clRCyuTD7JffFdmt4Z16xWx/pfa0T1bJa3BftPz0u0hupv4vL8lRntHmsZU7NwlJeVMBoQsdrubbVaOC7evPdV2P9bS8jAKxOCp//9wdFklsCif6I2hdouca2Ioh02ZugWo3CRe2nhFtGQSQcMMeYYY12OTWNmukhn3btCEv+yNQAkqgyLjr0rg4RLKR0EBTI0EjRzWmpF17kNCHJNPip+Etkd20FIxbGuE8pkO/ypXiBss2YKBVpo9V0To79N/0twq8JYfFh2hyIF/ZKEHhBc9rJROHwV7bVypDHA0wYDcvH/NQJFL0BroVZPTXGs78PpM6L2L7xUT8sQ9MONAaQfP56e6o9A+dCln+lxv3f1VpoGsY7Pwq8aWm21x5xfEV9bUtp6oW6q5AU1CXn0RsxAxwQrJjfTBcxRMUxZx0oJKM1u4Xf15ltT2hw/oDTOmh8rsoN39vu83aS9ItC/xeqDM6WmFmM6f5C0wgF9XcaLEsRYacbjVljK3BjIVnIWT9iSGkygkLbCUBYnpuo+BJIvxkyvJhrat5Bh518rtbff0uO6oRIGqy7xiaRcdiI9AHOE5M33z4LNKU3/Lm5tJnScUsKYo"
`endif