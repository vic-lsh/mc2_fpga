// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
liVu8kDtp8UejNuqdSf+22/ssRBZXsHML6JfGyT85v8Vxw4+wwd+fjDytXLx
UQrX82ug/vKZlBZWXQsqwsp82nvAlvqGv+XVVsxPJtsfR5c8NnvcF5vSkZX4
SlwWLKc3QRt11NRd6niBgE6zaP4tPQobHZSmjJZ1KQOYe2vU6WXAQ7ErzfoV
TUl1dHLMQLwCXtn9pq6mS7lELTga7IMpp4AQrAdwWqjvYPPDAEF6+Kz8lDYi
DJPrXT31bZiKjiDiPk4Au8nQaLS0PDeYxsCVbKWfr5LnizxCkaZtjmtQZqb2
MSa3bocAwGzTZys3iTWuuOBX96L2lpZ1n5hzxOR4Mg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IOfCzWwlp938/c2hJM+FQGbuSIq8APKtg+Q+laaYnWk4BTAMT9G61jP9Yojv
UBTgcZJOMpBvF9Ei7YuZt381RW79D4Fzn/txmODFxgt82ueHV77S1B3ZoJmi
xTd3X+LZXgPvnTn5GxRENTmJGNjf40sd8FJZS8LN+vVqCtGY8R+XtSh3nVJ6
Tbwhwe8wtBL+ATXvn/QaGGOrTk0RSO4MNM0u7vWj9/mNTlK3cGpHCMXDK9Wf
PHKNfTusTnVEysX9/mnF+xFV88hMS4peVQAuRBLZw1XicgjGwSY/JRctH6at
1ubX2/KRRQsDzFfBrFZ1pBkSv9+CxePwfQlZXeI1Pw==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qQkHCGUq/LnCYvNl21DcuM6g6saKt6x4WnoVmx1HmfFGdMW2WFgHl1Ry6/Zy
F5Zj9ysXYWbEE23/ANIpcRGhj5p8y6ikLh8zGvWbGJtk05rioa9uz94JSxfZ
3n06EA0sGNOuZPx7I8uIPSTZYcCTxsGEkzJNHhy8Orhqz7qLZz1yYjWZNsrt
WAdTNUxO05ZM/GfVpFrCxfYkV9yin309EEyDFK7QfLB0FhkRQFmx2ZlTwM7V
nbOxJRZVHb8YB/YuehFPJ7E5c3mWIrWPVndoBS5fuorYeTb93kNJwj4f/XLl
Xuo8fA4LbjDkSTlE4LMiLnxAQAs/3Nsl/0HkoffLqw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E72d8zY9HuOh26cki2mNbXrta8wJKEhxjh/W2Ow/dKH6bEJgcYAFZ/tqazZy
CAJE3f+m6tWilzqCGdCT6IAU9DX9gyRgie/azZQjxMoQseXW+UD4KCd1g1Xt
fI17yZRD3gMwtMM1QLmU/WD1C7+GZYu4wpZ/Db2vucVTBbZVtjNwGlB50F2M
Bj36yZPPdwscTHDvT1W02tUyTnF2Cx/lftBITLO1cjB4BLXyeyT0Bj4B40x8
brg4p5mIgQ5Pu70aP+QD1E7/eP0g5/JgjwFTuukw7HrMh+TinooA3z29vYrL
WDq3BJykGqwFY5BGyLXzWwX/0kbFfYioN9FnsB2jsg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LnZ+lUh3tFhgdmHVj60XT4vRf0EtZRdBJBWN6/so4fjsHhtLaEe9jiVM0hc9
tonXsPpfn0km11KyzyeM/1987y6dLicvqxsgIbrEGfc8pxsFdn92XI4kRmJw
I+ph3pFVCNluQ56UDyLL0GL1+s3OoD68MUFtiPP+zWP6HhNOo0Q=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
qJeZRK2dRIw/bIKSuso2HNcjcRKIOVtdenrivcMUhTVumxZMN8ov4PODuwXe
bPl5YGkkkiO5mQSuCxgyllVee0dHcAFNv+TF/xLFv2pZUJhD+IhmlLPtYkkC
i/F6e0DOCflf6XrjdrU/Pahpk/SjzmLZuNIcpZNSEkHjOclNAILNZsOrEwYe
/pVm0iseIcx6voRw88JKImw4NYQTryCMyy9ogG93PaGQRBOb905KR6BSon7F
KtSiQV5dwJCuWAXpcsWmvTYlXxHrJ5y3heVDZCisE0r5wk+u0CEq1QRBbxRB
lb+AZQJoGSixk0VUg4tCXYOQazAuazrp/ltkbZzE7ke9n20EwXIRx9Yq51f6
HgAhNwPSdy6Pljt4HXQsd2/OW2WhkBiYXzF9RCPsa8WimEu1phU+oUqxsb13
1OqCksYiM3dJ5epdGRGJRSNQDXSeOXeFPKH9lvNHE9vnepirA9ZK6nqScHOE
ovnN7TFA8/+FF0Dqk42z3mWogmuFe3o3


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
A2x/Hkp9Jleyt3X77J/kKc30sJGB7RhV3fx9fAuLIzUpb8NXQpLIvbUd/GZT
nvaHwfyojF9fxBXRTN60oxnQyW/SiHuoP+dIoDRLX8vpgKVsEGNfaqXIg8u8
MnRdyN1PV/35D7YzCMoVGP80eriyH7ROpHCR8mawFVTGma+dioU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bIeYf40p3jXRwZ8zPizDilcTf0F003gFzOJ5iEf5HFUOJRC6x0MKBzgDjffp
oBRiv0JVI+wvZzPfDJ7/hxU9aMdtQKDBmCNReq2K1BhYuHHtrrSARuNkAhFT
laZL5BfqX1oU8vx80tE3USWaP4kvhm3vf5cDQoqvzyYj197k2+A=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3264)
`pragma protect data_block
boCqBWNt83VIxmcyMtwN0qwpRgvtn0rzmz6UvjgBVgMlx3vg+KwlA7LdclF4
KOS4FHfUpjz/8UnXIVcBAUsDWqC9iB3onWRCEVtxBKYRfZ2dy/mKspvbeM0M
vL5xFGG6++p/7lwm9dB/zUt2hXtPU/VXLg9AjV2Jo3JFL7nrsh5BZsBlIQyD
qOgHpyKdQuQb/t/QgxXxAbZ6BAIsQ/nV2VDOd2mf+0OnnowKHErPxQwR8F1L
ucAzF5OgaI7CS2ZuIl9fKGACb1qQ4q6rM4OAUEkSI5j6eJQOUdhvL1AlYNa5
2yQ7dxDok6xSLB7u2HItwZF17m20IKUipbaInetAbq1uVgFrHBAu0f4N3Xw/
BGi96IucOqsnc60fI0KCgdD1g3BXvx2KlMGBlG7DRyGMfz1B+zRnZ64MJ8xH
2w7dowmj1XXl8p1hsf1O/WEcWDrb7ErJMACWByyp1Y+3hanVwLewp2LuJgWk
+VAlP3WnxyF5i622KUs2ElMHMs0y/QbiN5+HC0SEGe3MMc4E2G8z7mRkaV8M
PI0xR5uqj3i2grphSO7NlYLash7XhtkkgZoHtBUDhYcChCkqgeesbENpGAir
OM/ycHz8U3mXqRq4e/NgoLK9Lz1hf6qShFttM0/D0NH1qDQKP1lbcTQEymS5
hOwOk2Pig3ofq3tfaokkSCwu08TsFsJNvbq8IwTlXPJlHnlph3oxeeV5jTCJ
u4kFqNzc2JTiiaYRamX/7zkzVLhgjjh9AB7oxkx3jW9nzxnZeCb7HFlqrawN
ATGbzncJhLGfIkmSeuG2p7zJYQQ7Wj1Jde0UNqzBCynrHq5sxQ0NuDSl+fHh
Ms08uUXHAFING6rK2uXJwNt2GeiIBlObIromysmj635PReEBYDWxnJ29L3ol
Uq4f+TfnEJLq+vDWXhiniPyBWEiUPyDCwNdvFDr8MDszDaaxww1FttzUIysB
UBTyColBX5C7ik1sm8pabBNSsc2KretWoM3RxvumigW81SFv168Dae+j3bQZ
FCz1FxB+ppv0BG0LFbexiwivUdfGF0Gq6ldAWe4wwvk3EzPrX3Qdc+DxmtaT
Rm1cS202g+NKisqc3cj/jKr2wPYFQnLbg2cVG59pqozDqDBw6ghXEiBaVBqT
wV75bXqZug2K4Jhmszi/cMoWImuWzdAJICi+xMfS5jd7mBIOje4lBCIve2Yl
gqT2R8CG7d9MJR0RkD3eCJ7TziyBMFc/y/IyJGoqGVi04dSQDkYvc49fOxlZ
e2F1jM4zTNquzah57svZ4d4zCUjkQwe9fEZtitEyw98w/wLOz1ERQ1gZ2dyj
ZMPrxqXB7PE85JXKG0qiw9FA4XArOLgEpRy2Lzo9/xWpP1ENfslvRoR7qh+g
6B3n6CLPLi4adQowkcdGKA3NfdEG6Uoh+XkaIMTovI8pqRShNx212p+LqBix
rdXeUTMJc9iEZqSjApdgjemqw4hkw7IfdUXb9CvTLl8CVfj2MwH+wDF2YYS8
GOcKNiFcTnWdIgiE34GpmwtllKrXJft/aMY5hpLjcMifVNPpbOi2ulalq499
R5vurue7/J6G7jMVNaMWfM2Rfz4XRH2dj6JIpKIvq9kEzcFNe9rptC9Sn66U
xVpBgy18HpuxsNhBE38UtivurmgHZXZ3YXthjaZN5/grK526GAsX+kJy09Bn
QSF/SMmyAOb3j4gUOZCQfQrVcq3wW9YIn+oem2b5jcDNGQKO3sjX2Opk180D
oYWpfAChHsZMewHNe5QkwjKnvWUqwi5J9yMCWM9Kwgqqckm0V50HNbYZoLye
c+vThTma1ZP5dVClNA94Ri+mRlvChtSFSayPYpnIUR+Ui5wuI66px7SuoUdj
GQb04NKVjJgYRDsGb/jUCb7IlONwe8/a2XmfXDIKzTxICt1DJ4Q5a3Q2ZIKq
JoYLHBpzvBdAYBf8IdhSdLFfMDr3Mju2zEsrEx3SvfR6XUmeM3XS//dHE5vA
3auQTjRa5fsGjOEiYvl4ITlrn8IE7/dT3Mwp0yTUGlWsvdUrCH7eX41TdXs/
IwM0LZ7FrLndod1f6yu9G24yhwnFzt5V9Kg4uGKP04cgdSR/Sro9+4sfzcV/
ZyT2xHQ0+VuWvLWDm+Nhm1Z+wdNCHCgPpoVZxj9K5DmMNcRrdi7UIkHHPmRi
PCDlpqCVPMr70YcqRQh2KPkScAUDLbJpPu+fKrfSJ1ba5KXKgKmzTdIiakjC
Srqg+FDV/TCu+N3q6obbtXRAuJf30SXHH+s1/qaZUCNUVyAEziO3PH04yAmJ
0wCkyFgVJ0h85FhcrKOxAV3++rsifJ7rLTJRfoNgqvo6b0Mz1M6OKwjqCaES
4lwYAmZt9mlR6KnL1r5nmo2Cg2IyS+IDSVYxK6dr9aK6Eol2wYZyhN9vYTom
91nH8lo1IgaU6TYrlX09oO8NxrNqa2MhiX1VoIg9HLg73EsWx1qm78f5AC8M
aQkwpW6cHaAgdMbvuUr2LiYbEIym9Z4+fwWx3uSEfpmotr0X7Lm7VQqqFBOq
C4llysEfjw/OMPxkCbbprFy/ZJdG0Y37hA7NryYwGdM+m/kRviKHX0p39A8w
DyP5aVW4QUK2+GHnjsQ4nI/DQzGyM+551h71F4X9ClI+kKdu8yDAgoVqR8ir
csRK8r/Rn0FiaAjvzPxCBWd9OWRSW3er01wSiYxa9L3JGj52YPu/X5VVKlcx
Ke9azVPZwLfCSWwkWaprRtdetOWbMS9se9BSt5tmog8yHkf66lpY3eacC62i
1Of9w/pKF80LzyhxqLQMvdwPer7tg5BrcF1I616RrkKqSnvvCRG15rcIfFek
DYcSNYZU5xMQRo0mKUt9m/I3qWUjc+YCZZgrmionbOEvIn38JsGm78scP/is
v0KcZI5lFL42OUmzzoYQudyMWY0OOz/nCCkjZF4g5LwzZGrSZDE0C3FgzIr7
UhMD8VHsbStcOxzLdA+w69H/qNd3q00JsvbDDbaOcVeR1DmUGkDMvXXv4prO
Wwrd+oEfBpuT6Fr5oZMnL4yV4oOmv/PcJU6qm1lFASUGOM2EGL6g1u+BO9dn
VNskYH9gkArZwGK5TZWl/hbnYjGZMrAcC7FnokO8LzQX56U9WChvj44DyN7m
ah/MxqlQChrIJol3OVpQahaereKld/d5uuLNncQMrwMrLAdu+etj5DZsK/BI
rXW/S9fmPGj3/UsxLp1cTRIPtAQ56YYFfwi31wRUM21XFEBY/+UFtCjIdZya
lxkA7omCMm9BW30+zNmyYjNvfGSS0aETcHzw7eTU73rUnJypsMLfX0kZQK1Z
2dsHQNNLiUeysMr4p3QP1CS+lKgU8wuQKmlMvn5ShQ3e0K/qUqJSED8sfpMO
FbgDr3PoD/8q6Y1a4aM2XppeeAhbELl82Kgf52c/vSyUMzPmY7jW8Ju4xXmf
7iRDsNNUSyJ5mOsvVHbUa1jGuTkNn/6tVZgYBWwsk9vvCmYcBntnJ7pVqz/g
fLv7WpRliwjwpyzDVhALIGeMbqiTyNskySLMnAFPe5vlTWK2eRHoghs3bapN
JTWUtRHuzhdCIWqn4R6JuVgd1Mi+jxR1wLY0hHlv29p22X1Umpzc2R5PpCNH
tMINgu2PbsWefGkiG7uXY6ke5zOq5sxEwAW1QhYWTbTZh24fl/n9SE2PaHaj
wFSk2Es7eb7bzqwQZWOWxiWLQSvBvnVOyc22KufbkaUzKXSHSPM9QE5rHsJR
pKY1V0Fk0EY4XgVVPohbqLMwNE8u7OgrQZZ3Bz6r5Pmwr2Kk+WqNnNxy0e40
TB+tfmfwzHlNgMmoYa5cDydBlyufxz8WO66TN2yfiWCWqtswSyVKOSajMcC/
H67Ai7Tsfk6JjF57G3InWa6rvqq/VV3KcFMGPn+HP9XmcHcErHHRGSG2QRXT
CKekD7HuqjjA9W6u6o718WA8cuuDkWnl33zKULEjKyz+afiAemHpvADa+sTu
jaSmvPE9VPM2nhJlMTuGnv+PKPT/J7wL5HL+hOXsogDDYTX1sHBJMi4v0D3M
gRHNJ7drGLaDM044TcxjEF08LsXB/rTMiz4mPIz6ddwXtCWTwXM/jekw29gc
Fj1Ik7C/Gn2Q6/DRSeTdz3uN1e6vzrdkh97D8JU222IWpl7JljRfoKIPZfPp
b4IFIKGQiayGDJ0EvU8gr1hXqlWGGksPhCwfWwoZHDxhhDey2hWFTs07uKuJ
OJ7BXSe9nMHmQcawW+Jw8UVL2RfDkjyicJ3x6LHKx2xCc8abC/jrSjvpQPGx
fwEEobEohuXU862RwZxcZ10DwJjl/HXnxA88M9kMK5yRJk9+C9adgaCbPAQ1
PATsfxhxf7oJxEi7OXEWbL7pPD2yOqet

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "dlqcmJx9Qhyx4I7awZaUP6WRSv8nfkoLmgEhCASpkeIHA4CtESUb8gmFSOphz1tpweHgKgEhVY3NDxZs9BPPqKGftfW+o/FmAO1kFkRP3v/8+n0jV44sgzhLFVje+nZmIhlpd9GWW0QF8qOgKtusK4VeL9ZPuxX31vWE7Pf7/oyzI5BKGkYSwQrtrs1aukEDDDFamxx3mdAUuVEXQ0W7N398UWRq97SKxYWZ5u5Mpejgp1VDpe91/zwj35UpPwJh7W3+hqCKJLId/TaYr4XaUwY0jWxJzcbuUYFxkgWDJaV5SeoPN5Rc0vIFOUxb4zZaiVS2w9rTy3yFg4IDAVxy9wIhbS3mpWIrr9kk960sUDD7u0yhnq/B5gfgJO9OqeXTG4P2JbecrT6wm/y6FGDtMz7SQZ/Bk+9jxOD/YIXa2XBUHqybCHfsZd0sCrJnlL6ndF3q+oAn5hmCYTEABgIeEtS3QGwZXwnqog6TCE/cbgMUXUAFbD8+/uffhW72oUc7+rblV7o2MOzVX6Y5LHc3BZ7gp01VCJ/I0UrwOhR448FkhsuWdkeH2KUN78PhN7dsV+l+X3rfGh63fpQwFgI/u6nmfijiZPF/rBLaz08JIpQKVEZlobyZyBKv512Qz9apD+U5yX9dVZjvWYDyEj3bCgiAhi3AN+p1vVYPC2zo1vNppSrFqLqv5n1rJeTOY+Qv6ce23ph/4fKrpnQD5r7FwM0f1nD0mpXLcsvstssb1i+4xnmYoxjNNfua9NvXhSSknWckeu3dOVf+PKLZsz+yw+VkOo9nF5j23FnO8yfQu/0/rYa6uXll2uSaYm7n7+8Y67Lu1Dso/a16stygt6Jl1eT5VWH+m9CkGLasX+i3aCdiPcs126/XAKT63v3EloPI85JebgG7FLQPYLxzNWNGkqTSbQwBqg8+JJmFRXedOSQ+g6LvhWlVtvjJSsowDwlM0JwdUwrmJcErRqUjP5jPxYQI69gNWoT1KhMzEffZQ6nmzJ6dzi/kntpFjrydHx+z"
`endif