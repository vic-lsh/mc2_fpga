// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
h/8KDKr2rt7ymhJSq8fwDh3/+7UfiPQMVAOynkPjtDYpg3KOdck45EWJKvmb
tHoSZMR17hW6kG2UtPolfxxMNWE8GApx9AC7C+FrJrk9WviYcglAZUW56EQ8
6WjAVIhrefR/VYaqszADM1FC3S1PTy1M/q8tkK7tPgG7AwwhRFm16fkGmVFh
oRiNwM1igMzF8P+L4xAy8/yWzFWbPeMwgyxsZsKLtPLsAAYz6eWXcgpH+PQg
0R1D4NpZlsm+j4LOFIjWM2x7fuBVoeXNiY08n+c5OuBSxHOImFFGSutV/X8u
9lqQdkGQXRHfyHGKRzEqlRbWa0bGV2Czh2HfaVzylA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pjgn+rZKPIFaMUmGmm+UB7JBYjijXsurS6HiJleQZCDViLgzK9haZ0ZE9ahr
bdOczpa5NDTvxznITxK48uUK8GcNHYamded5tO6Lcpdfc3I7J4JgkIxsxTdS
J1kuGFCR9nP7q9iR/BCHB2R1R/RWE0p8e7vskWqVlUHxslJoQbZcafaXIeg/
DUhg6PqodC4JAr6K35r9Lb4cVmPiqqIvCTvOq1Gz9uWfi5NZLOZ9o2AbBL/t
DgHAeAxQBm5udrLoSiZ2rfPGwjIXojy56SmpDzowYuWanpGIxQ4PkrvsZqiY
bDemcGSw4NLH34vtaKvi1sk60qfETp2GZMOqdOPzgQ==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UzkICwNFFariHNI0W36twNF3Zin/pCFYOMC9o3iXHJqTobCT251rEVDQs7bJ
gXHz24o9OzQM5+zey461X5cByO8dpeIcPR6xeyGgN3Jr21TCMrplxj06g6o/
lWVTiR+A+1jTaxdyc3zJQBFYZ4odfM3qZYfNZcSymjLLTGD7PWF/1DXT7HnF
IrSCu5Ayn3FZlh3JxM2l36DZwHmeslyQyJF266BGeWv0pZn86fh1xA2j9lfx
WqIBdiOaouZ01jaF++QAnMMWdpqL8y1Jo/Z+om3NmsBAbwo3iLbd/LOc25BZ
uGMlIUPV77Pe2Cd2GqGx04zuWMqRCjfJXYT765Txhw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kQkNvToKR0HVmg+iu9ck9dFClsR4A43dLVfNpBYdy+Q4XUxduWb3Yq+GLR3f
ga9D4XB1qXFxEXjJakfjdzfTNTWEFI7fnF+abmzROmP1yJ2zHHP6Pv15+j8w
l5QX79VimfzojO6UGTiNbHpXhbFZ6iblwOFzvjaAkp0SJz2ZiUJW5VAvaEdn
EH0p/x7WchLDPNRlg7dRwaXOiwR54E4tLGgjX3ufJmHkY+7r3ROgFEO8PYMZ
SkolxvS3DFjlIFFRoF/d16oIn0SjPf7ncArM9T3RvBQrAyr9ILlIWIRlwWGn
tjM9S0xGwoeZSFtFiEIk6JhFQSfm/xAccn1pmconsw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
W+X1k2DZHoCcagADjN/kf2I/o1WHvd0Z8Alx+b6ysJ7a9lxZG+RxJpmfjagp
Fd8Y4FpoRbSCovyqyNkag0Td26j+apVyB7se7dxxYpNhr6dCnJ59L1lBe+GL
UE6WXYQfm5MnQU63yTkbywfdTs0nB3tr/x3rGcV1OCug8EpnGbY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
fJsP85yO9/O5uTlLa5PlNmwgpPNaT7dqNlgi+veDmKoXW1qbNk8Vam7kEiFv
Rk0Vt9DT0LzTE5RvhhxoWJ5ZvEwQTY3iW9TpPQmVnN5MiLUcxesOeSpEY3Tu
kgsh91UWqtHzqAS995+6liLSyI76mZ4vteH0Dv5Uf1xTMVN7aK7nJPB1p2lq
de+1scgdhur8n4J29MUHZ6gjc5TlSYeyl+WDr00XfTBDlIOhSZqNQCBjzKRC
fkLojacZU4VSuRQnIj1yFuIRouaBvvY+ipxEX0Rh6bZ5I/T3n7/0Zs8isCka
ETxpvO6CyVTkmlP5hN7+CeS8ubXl3LeGHPlDLqeZ2SN1CPEykrXC5zSgo3hy
h/dKtQMwfqndjFO2leMcmsWQ2+X6qaMrK5mdIaqeFiCJ9+yeafyYzJeWbcRx
EcA1WoFR+dzu9XRv7MqQDfitklg3LwhVxgJJbMTpkTP1i/TAgtv1lC6/up8p
cVc3vNFCQ4jFb2NKw3NN/3ukZku7pecI


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
E627ymZNskmB+w54KtE+A/MHI+YDAIOhyOux2NETI77egmKRRfxWuCmSzmgA
KAFgfMXzWgKG3O5QUhEvDiduqHqYVou11FU6QW7J2+b8MDvap6gMKAekJqP7
HPSLLJaCsAJe7r6SMAx2NV8ECdcJffhVa//BAY8lpK5dkbKheig=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HzLDL2ep3UKqlfxleQvHxN4EMeOgIJonlyPxY15jWcaKENgR//S3FxF1g5AF
GTjMkqRsGZZwmDjILwEFbrvokfQuY+I4MgpHTZZX1mpqXujjdcTg30jG9fN4
fsncJSFUy1zXSIiEs5uECf1CuhV2f2QnDROnPs29vvBV74HyFXk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1984)
`pragma protect data_block
s3pJWjIWKROP+YJ9weqJB6knVU0d734vhyQP/Zkjx39HGIH5KIZmxiJB+SOn
FjIKkZMya7CG3Zb4zTR6OpqTJmNfx8EpI5DW/LMSHiK3Gq0/3B1AfrXFBBN8
8MD+R4EAw9VcfgAWkxL+bsw2Aa3poWauJebG69SZxMDeDIgnKlQ4nEyzXpKw
noS/lAwa8V0PqhPQAQ5Ca/kd4C7t0vFOT0ePgcyqcFY73U8IbApnYugFxqlB
BGCOcZ3hJbTUQLdCfp99IE1C8s4AUT3H9EYeGkBnb/N1ZjL311SbEHdgl+u9
Ab4EyqPC4jGQ6WgLZkdOe45bExedyLQl1YLNcrxQSl2AijWIEuEfan4iLDIT
tm1r/gKhVf/G1IfiVPoOcbU74w2HFhXnamGepcIM8zNUYoh+cvC5SNA91SH1
309POwomBcgomW/AMONx1lNMavAcNwKxJIZkzEnmYfrZoybmqTY1tvpIatAC
F/hDioY7+V3vaUFgf9sjkIu62BHcfaQyq6Y110tBeR/0y9pemjE78zCS5L7p
lBK5NkfVul6SRPTo12bGxl1JTc7R5rAb4E9sjsa1xEUhk/hRAdWk4CMuafV4
Xu6auCTJ8L0wr5IcVqPnPmP6zzZfLWMo6wE7garEYEHhPFazCo4Z+chWlQdm
zpuhQpiPVQft1nBgAey/jVDNiarwLqWC7Tq+ZB/xACLrVF3Bx2gTxAULrMxP
21bmNXURZfB8pz0MltorWGZk/S6lgBTsfwL9JfmTHvwt1DcZ+g71GmYcqbDU
bSRlDiUkpUFHYHt9JY3nkTKfMFFAvkcSeOaRd0MfS4j0i127N5ictZZHzsvu
54HXz9aVKEimx2Zp4ynKAfgAkdyYIE9VTsJNgIqat2yrj9czwpsEQDX6DGzH
xq9qgD45N1b6UFNFSZlN3Kk94ZuZX9CRkhliO9SvamFnyzeeyT+8MQHrWYG6
ihdvH4EtNhFSgNaDkJ4tMxz6CUswnx95C9TlAiGyWX/7LKxFAKy4eQtp5tJy
byMihKRM5Xo1JE27bzeO0N8xSWOttmuchgcMgoGfWXEkPr2QNKeG9awj/vxA
CKGE2PQFWbPd1JITSL/uPfZv21mY4SHpFMp/uweF8lA2c96xmkiefRUsUwVE
2f4AMloD+D+iwBUFooydVF+3PCCjoHcBSr2f1gKDwc6oOL1ZhKXEue121O9L
/7/5fgkinRZZ6I9IQ2kduhrOnMTuRz6CFl5ST5hzK4SzNBGcn9uDgKo8F0Ke
8Pon3pysfQVUiBRX+OH/LaCNmXRhU5AB92S/XHoQuF/IuX+Cj9enmKb5hk0T
g5NBY/MJhrImzAKVrhr7YUndLtjZBZSupoNKghTFZ93FroPRS+MLnsMf58/S
wEvhxcbGKsze34k8tUxSUa8pMKHNTCOu+71CpdMJhmml/kzPVr0X3GmUNLbe
0lQcUl42QdTgSgLlypjfYtrLZ7WT2TpG7UE27JaAGKbWp7ZiMqDc4IufnFyD
fElfLwrkgipM4rt3JLjPs/S5hjBn24OoIWI4216VF41onLPayCMO4YdApPtp
UHlO7TKcsgw/tVHzRDT8uLMKa0vnuSuVCa2y0bpY8nX+hIS0QeqE/+O7XGFA
bhnRYLCuJBFqGGxK9mq/surQi5WjP/vEpljMOUvgTX/XVM1eBALZGjk5YDoh
smemCgmTbnlP377cphonn+Ymti5VbnCICtpGyTgso5UqqOw40AJ+DIluk1Sd
qNI+qNY5RXLlPoyaMye2L66fHacAqnmcAEj295bEkl5lOsCku8n0hlQW49hO
rh9M4I4RzmgFeJft/ii+VGHetlb6+NgcwbSd6L3Jc/D1AjLIPYBMeOg7GyLc
BgmJCxgt2LtZ3Ckj2pfrhH5DuUMydOnM3duSXgMdBcGqpWZqWhmrk0PPUd5X
AO4GDMA0P0iiKLHnJqCkRZEp1celYZnlCGYT3XbaMCz1n5YcRxggs9FIhjkF
HYLKlXLJKlLQWDjQk1SrGG2QAGOWGr71sW/DyiKz9Km5SkjqI/pr49Vyx3c9
K8dwHzj4Pb3naguwprJoOMiXaWfPe9GbELtZuvdXX55PR+vRkyOV3Ro8s4Il
Hw4IgC6vXpDtmEZMO2PVSRtZzmshptL0bkzpijd/n0UP/qwUHLa42k87oT3K
xjLiDalov0UP4MPRz05NxvdswwZOLwt2ZSZ621/ORNwIJZMq7iewX/iyWlgg
3UeHU7GLj8OAYa0fu5w/gRVOqOcWWdCwqzcL1YhlH+eiTkJW6rHZJrSqKRQK
b3Rl7z66hT0TVkPSTm3Ed/AsDhIFFGN+++bK+GQN0DKOMocN3jiBl21Yy5R+
FdU/QPNuAEwTbln0QRT7j6gEwweBRbTKwJsCCwQEQ6b6aiJTmS9iFBhu7y0G
fdyOobcfWN9lKWE8e7cHaCuRFafA53Lsd54n/wIbs1GMrOc/JcXHn4Ehk2n/
0NrC88ej8rTxa+FZ+YipHFOmfzSQSw/qfeK1pYwGVPmrms8+ESeqEDO62sjM
cnsK/dZNaUav1a+nbKd0o0CO8WIRyLpLv4pX+cNhpyYBtP3gVxpeWl/qpRu/
yQPNZ/He/qjMa+wX4IyBh/KoAmKSheHJEQUbEQZOkHZXM3KvoelWIvOOMfro
0+XZwA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Kttctzi5aPKQ6vg9w+1g45z6Da0UaxXtt50QPmQzmLiVao+5Qg/yS2eSRK3c1uFoxS+G6ngDcAKHm0LGGibx4soakCOjaaRTqJmqblCXBo4qigRRJU5sOpNJWGKfxZC9LZLfFjqN04HCQ8ah5FN3P2yNU1iObRgi2dEkx758LbIsGmsSUmn36d6MTHQGWCnH/AC+2pgOY84Iul0q5eg7DNO6RSxNOih+2JmnF8szbMML55J09CbsvunyySvVbq1k2zLZi/VVeM2qUq/ia3pHCcC9t4EcobWVpg7RqPjYZ9LDvZkizaayUrY3bY4FPFaiBHSzDM/fuZlyIQdTNlr8+rjEVPo0F2cW343TOplNIARyl0MCJGjWuqTn/Rcgq1EVb7UwFZzB4b1Tw4ZSOvh0C1lQUFgSgadhsrDsXGK/YVy23k6olGsUf5qhH851p7Vw1rMcckXveLrWTBEd7xg1zx2XHZ/Z1bSYgFSQbK7+e1Y7z0LJLRb6yfzygNswBW4jjrLcnlB7qruJ6lk5Kbq1lr2/RV7BENM4lXaWllClCG1x5wQZjMQ/rn3ZFgaZnwgfxyG4KCMPBuHHE1lqJFLQ39jWEId0pGmdUPt3aTxrdC9EDNFP8VQzlyIRJFvboBAmnq+298TmsIOcefQFUrHsqO9nx8UMR4SYyesEcE9jK0GuxaFilBecsn0NtnlWp1geb6f5enPdxSgszdlkcP9vPREMG3xghfAWAwkH4TYnu+2qtJdndxOecfnV5JCa6JbyYsu0S8w/2GdTUn+zcHgwVnx3UUc6DhEiHdd76wC7vCY+5Fxk5f591BlNj2NYGguql+zAbkTsqIesPir8tK0p6fQqLq/3dThj2d1V42FlcZgmHHQRcG+SxWCo+gVvvCQZHYfMHkXfOEoi8hJDcWMORSKojIxPDaNLFlAEHa3717+FVABlDgcwkI9Lw6MdyeAysz5S4KVOIIU2B9ahtV+4gSXw+sXeLR5zYB99fXFycZqVRsDjoGX104PMl0rlcIvG"
`endif