// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="24.1"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RVwf2pMX28oJgcu5rDsNzCLiJBQRFjR7cV3M1CeLQIFTKBABs36JVFpUJS16
Vd9sE5hJHVLj2HZh4SyL+rbGFBIa5pr/e13ccV1eI0wesqCxodcx6DmCJAB+
YEWreRXJb3d06WrjFuiUoVbTYWScbhYU3CKJCLTHORqeazYxRRM9J2wKvrZd
5kckA53FGEY68iDS+XpHwAqNY/4GG0pliL3TJVgNkJNGPIfRgoz9kg5V+gr2
89PGQ/HI514pbBMzodDvyAf562Gf57+H9TuBLN7nTg7leYrdViQNhsLa27YK
BnfN/xW7QHsFBh7YwU1EJJWBYsr8iQvWSsmhP7hkrQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
l8NqcBspS41D+D1gVR2egkU5Jacqn1AVsHluTweNvm6xoLxOQr+NuHaK72XQ
6121qgdZ1B5MftjPgb9/9yEJEqJrCOTv4B1t3Dj6368quJ9MuU4D7+/97Inp
Pmn44mz8TRZ1wRTaP7nLNANjCbHMu1UVEn04c8wZmiMnM3IxMujj0fqZOW18
p79boC0jlljNo3eE65+wTYuqdITDPOpgUeYkIQ7DFsLImLusktjOyMKBnp2g
zyfWJ7bKFE6o7qQxQT6lGQhz352nwkepZLj42cWIsr2wpHmAn8qgeAj4ZnIK
Rxn73vmAvjqFBf1c/DeOhX3M0/KVVpUeq1dWastsGA==


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-SYN-EC-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hS36nh7HOqeJdABDjJw404c6hA9P7XFztGRgkeuj9xPINLbSXeZ4rvpT/UZF
x1eo0Bvxkrq6q2qDZbQYhqHGKnhPtl9d9SQxXf+WEbciYjUw2wAf60+7i+8J
DsGxKrmKo5dd3/eefsnM0/RtoYArgnk5ys69Zp+78m5rvGBkXOzOlGgtxCBQ
J9fs0eWe3f44yRC71JQh2oxCr5+Q6rwEGUbkMVBTKjwg+a1Buw2mUzv/p96I
SU/1UD3kzDmA3S5mLeQ3meFeM3cw/rNBoE2sxxqXipFL+xOu9kA6MwpAZ6/y
MAPv5TWj6WyK+evQXRtZ3mYr5U9+PEAgpz/B/WqneA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bQJbYy2AmGpsZHCaJJCnKBzpBLwWgi6+5Q1zEjdHEoajqU4zJi5mIRQ6ALib
SgBlR2t+QGJzlykY4xzBo/iLYp1BHGwD5BZULy8kRL9JLX9a6smyP3jRaHpF
3nbAG+g6cCnOyBLVZQxXBSiSTDHU7K0aeDJi6ylWCL3QIGLtdFPyFVaJPNmk
b5qpISt3NuwpEPKjckIKDPth4G9qiG2m8/6goJ6wGUvfkn6KHRIZnWpCKwS4
cmHn22PU4eAfLlRgYXDxeMG7qplNm1SZ7U7kiqZJ3qbXGBoWpXAOssgJfLK1
48mHMQACxr1Y2CPeL58KXlQJMWypEbsZTqhOTzo8Lw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
r/eTfH+jmqzntBjVsB6skxYmktZtmTwGaQhrbf//hy3RuG87IG85W0u92VY2
xk9RdaJUYVI4URVhwyMRvRrH/O5ffU5KUFS1CpDHQNndJkn/o+v/rvDz88Um
Ik/jGnUB9rhn5o7mZmyAcWogC7S7bcZDAmhCUcC8INO11klW/w0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
A8H3l3guDLFzlrulvfzPX3761XMZjWZ3aNPRkzk17L4FkUuHET3V5pXbvbUR
a/cCaNa8f/Mc9tYf90cRsAI9819vDjRyHQskr614cAB/wLeiRRfus4TrxmoQ
q1T28GxC2w+v4j2NCFY3ryHBu+/5X6fe9GqQyV/5rgBeyCjaMfdYoPPl8EwZ
i+ql+4SIJTlYg3MwZe73pmPjRIRkKs7+TuYC7jZhdY8o+nTsBbr4GH9VuL8r
DrnNdqWNkDlegDE/y4EYpTronFGGS+cqHHwiZb7JX5vexfZ01YEkZH/W0sqx
kYz+PaBJVmo3+5+4vIkKOy50IJXwvSBvdYqzpV9SUZAV0SvXsHw6ex9U69Tf
5MeDMDntsbzxxEtM0aUWXdQIx7nheu6C+aAX9A7b0wMJKJ/16dXyZdNLV9g2
bFrdbmOhNG6b83MZEn4082dp4L3Fs5Tw1wR5lQj04nyj6Fxm8zFQye9sSOEx
+tlZLOdw2QDEevamyxd5aZAlMmpNbNuQ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fbqy/VpckEc2x+PAJL3mMl2geGaGNMvykIBvQpoqEkEECMrr/Q5Iir0PWMn0
wJ+5EWsZBjSkRfuZSUamp0MjVk7ACe0Gx4Nc7lMvVROyPZfG7BSZm2k0JLkN
gbI/PhluaVEhVmsqzRa1tm7Tmv8jt6tP7zYhD2jm+efasgR1BaU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gldjR0JvpQ7a95tUukVotg3ZJIWxaJXdywFUBYMx1/AZfSHCDhTChLNBcEL1
bLhl6rOIYmdh263Bq9RPdUijsT2jdCjnA5gM2mDOAlz5vFVMywSVZWh+TD0U
sUJ5p0VpQOX+9x5BZwk35VUmDgTAgPMu7cy2GleadBZ2bzB1c7k=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 49392)
`pragma protect data_block
rqmjNX8dUFiYv4kYLocVOchnhGXDSKVCNB5OosWfTvvcSsifwAtRWqHTdjKv
zM04w5rm5oB5RPJsbOpa4hSHUo/5rSH41Xflj2yAPhUSzfZVohBfYCTds93T
USCGYdoryL8epuCBfwhuXmu0mkgQblLr2uK4tMbbyF/R2BK7rMlecfNIV+QG
z6a+ausZj4agBuxmPGrgBbL72kc94PVr5/zNWw8EONTY5+3ZLtsRcrWmzuoC
XXYMRNFImk0SKSudjkUFMZZPY73gPTdGbt/BxDH2rkgaaPzAI4/HsV09Q5Uy
CBzu3InZ16oSrRJC+24Asj+6947JY5ILAdwPqKq1fMCfbhzyo20jveT7n+6a
FHOi9D4PxIs4qTNIezbI5pvbr4ivsYcoGVaIxxxxXuiRnMqJAZVWSEcuaTzX
QkFSjR2n5rgoehoNqKLk79W44fr9plbucKKOYs2CEIXZKz6SS3pYitTE7Ysj
5F3rkZLZikdQvJ8S7cu8rt/ZhnOgSdEKtQDB9UHZSEV+pPrD71wmO3Nqo5YS
af523hJcCrBuyVgSuODFSlKYPEQ7mD96jVusqOLZKDcTSka+fqhLShwgWf1R
vlf4Kc/fjsXc8n7qrMXM2ErZRIMB0R53IIqmPPE2Jx3Ci/jHm5y7lkVLaJte
H32YRh2+I3Iw73+h85xMmqvdDBhqqk6JHxmIIjfiIXgch2pjB3Y4Rol8Q2tt
uPnTXyuaj5W1a632pQHt4MMFMjypn15cCljKVR0yl+/U1kNCqNB/cj3NuNV2
6bh9/gjhEBkB9g8rPIV0Nl+niQAsggZNXfrnBEzMcb7jPOU4hqLNlAsGURNP
O/TiEtMPUN0ZOT/i+Z1lhwcVcx4Lyzkf7Uhh69Vest4P4mTHtBt1gln3q7Ip
F++bw2NMRaUK6FqfOTzNEabSxm527WBMkmfBkWS3To6lWCzq/0KZSt/AhDl0
LdG7K5gUe2ulug0+FdJlqvjdaJSVO9xSzzYWcgw23nun0dEn/ZulUWFQgWN8
hwKL0U6J5JVGk9qldhYHkQIBNQ32yQ7VSXn6NdslVJIhGInvQKe7wbxYcHEI
9jSSA34LGQXcBFakLSU1mXLODWqJbCjLNwVnNYGe0kxjcgzCdBA3oeoBjtl1
qBuRy7hUQXYud4vJbYx4M5RGuojj4PoCUAnMRTsz0Pl4RLOjZ3qd0qK81ak6
3wnNX6lQt9mKr1N6YKLUELq+PT/GFY371P7y6hwDxZoX3GqtU537Qh0X12j1
4WOlKITDYiQc+roiPBu5jht1wB4ZO3tDQnkEvp+sGqP/EwBt1V5W1bNwNkHp
JMN4hbyPlXH23AE3lOO6S1om4c1rsjiN1RguxpymjruVELrTfhd8gfcyhIXN
P3z5kwpgVc5QA9tK5Yd/kkTe9QEgtIhM+aHTVyM0YBz3jFiudR3FTcMoPKOq
cHoIHhdnWn4IDqa6cz0zARp37lL+4ojsWuR6nTNfIefvk+2PIUy8x+criGHH
RY7cWGJdYI5hJ6wdOHcmwsj8ZmJ0EvAlVUHWFJ3R1o6IDVlGi3BLhKa5SeI+
L6ISKf6HzGGEFLZJc0w5d+zH1yajrGshou2QTyZylAsssfF2HEE/Z/ZnWLJn
0g8tbqzOmlMbGKLGeKUek+xDkmlj5Bhv3OrTNX2edoFNlvwjupRNJzsEfzCC
l9ISFK1hYM9kYr7mdK9X5PyVbZMIfZCyUStsnQEIpzATYOT37h9i23/H41Om
4p6XMFnZn3JMon6oyidHssFers9dzbL1AgkexBY8goIxPBVZqzJt7ULU+6AO
O/Ke7jpk93PnQnNXrPxmcSaM/R0OGqOxvn9iu/MDFnAcdPwilZ3ZH14loGzm
aLkY08QEnCwcXVqw6nSiVMMI4Faq47nuQn8oPON1s4NOs5FFzAnQbBdUofpX
xF9i6go9GcbN2Eq61z3VNc/7+R6+jLA9KQNWBN5lgufvIp7uiJKjkbfqsas5
A2ZEi4cwRDIrh/JozFN03fu2LMzRIqhDbEY3voiaB6Ckq4hd+SkkAgPy0USB
m4IOPl+EN+T2FECPoJTAmCmRnjtwZLNjIqV3EtA/KpMbZpYvuO4Pa3u6W6Ro
6A5Ft09q2d81rbSFBsDjPemtsmFANmmMWBO5Pmj88IIk3AdLHDjgbc3LSVoV
SzKdXn7F9qVJPfLv4RcxroavGJvGkHhBlWZ/01Ql9r++dy1dGRidicwHfm0O
RWGINcxNwSPNqrOPKb5FlUE40hjtXcQpTgeLDrWO/7Qe44GsppyAbCixHWcC
tbt+kGygj4HEbh1oRkh0QD0mvMFjE7ZhAHYu6NBkatuc+TPRLVbmB3FgHh/p
WqXVMJlob62J4FLKezArdJe4UpUc8GvKybpcGqDHepXmNAdzV4n+slltbtqY
0K4vj4PIt8GmBRVbcgH5E3G3LUkMMzH14yTI6zXB2vRWeR0oQzhObIDGpSMg
nfzg9OhkGnnwjkd0aYESWPcRr6IZVjEBAL1ry+jbV4JX8Vu9p0HgdpH4HtZ5
GsvkBpdsclu7lhWCEwsz5ehCjT3qenkXbqtdZzmcw4vHLSRQsiQpV7CIdz2X
RPO2lwadjbCDUd6mnkdrMDSYzsAO1jPEMKNQv9mb8T9Oag0CWznm8NKyaitd
ctDZVkWHKm3EZya51A0IyphAPHMlv6IHgZGKPVqIrzrtMOMqpuBJNaur+lNk
tGiwa+OfSJMzlK1Pe2p17fXPkik3IMq4TQCpAu1AYrwhqXZwblvqgqC93/9i
P1+yN8dNYFlw/dq/Rq9eQhPSNA93e5lMWWYVCq8cA7zrHNzLRwiF26rHpaWc
YA62PhbCPam7JmFplDisQxP+3NFfhWBlWoQskUlpq7SFjWsve9/2EEjEjdVn
G/00EA84mcFl4gK8+e+B1WG9eXVhNHlgNGrleQKlv3PaFYmILdnQ6HDIGHOK
OdBxoRLqYUHbGEL5i9EG3J7SKPgT0wdEdeWdtUGxONwlejwibqgnGk0JxGRG
8fxZE6Fo+juetKHGQNhOLFOQDJj6+zx/WZpW2olZ264U4aqPM47gHK49gdT2
4iU88usnScEAAVzjKkfr7QLztwy8c237okaAI5asxo2FSf7VoHVwdfLTfHLt
UJoWPt9vU6nJjsjYAUFA2g52oFwFnPcQLnYUvBAE4Y5XTzsjFRYZ5mVuX24a
BbFPZoMq5PVP4dtzl5KBqxJRW2gf9i0Ps6AyXmrBAf+bfnngmxX9btLD14Nj
zOY5VG+5qDoMh0BlrHbr+Gzlsj1yW2iIAc6if7jC4rZjghWF4y9MpBC+qhe4
pKVlxtgmqI66HgskrvMHl5XkjubOalBkxtfobazwmiUySjGhXAO8hVvgwOPI
P/CxhiUulpJhsFYQ2cyBj8wii1/nedV5XSjMFNpVLsqhb8d9RzpixqSk7KO1
JhBwarHObZpN15VZD0UxPKjaEj9vcQgCVh6I75KCuF8Sw46Nf121De5/5JvL
rwgoj5FoiMGiDMFQ195lFnE9ZpyHegZ2f8OTdg9zEbmAidlIL6RCSjWuWDe8
oWA2t5yc/SUiZjEQRL46ZnUonnVEdZ1IT/6icnwDYk7YlB6/YkXljkT3KHtN
r2C8XmfbV6bKIdapbQP5WH3k4dc4cHhfmAAyD0S3asHQfrzLQTPm+/2cDfBU
FnH+6X2E/u/6f7rxNfqWT9uaInWnNlSGZy/W2I0LMAXuWYKO8uynov/ZwMCG
UOae3FGXlYsFcu/tKc/GiygRvnHNBufWP/ssztQ7H4t54AdI6E6zSM2QqpIq
JAy3Bkdsi5GBZHmonRO3DhKhAezIakykxafKVp/EijTrnpGOeueWibdHny+C
1UImcZFxdUnbWxR7jheWGVfP9fpsJQ2M71V/cbYtv86uw4L0LYZCvjEHrix9
zBrhjF9ZdR0us2QvcEkW9035ieZXjJkYxHh2pOHb/8A1XMEC+TUYTUnmy1gj
0yVrz0Lla2Mgs3DZs0KkCju07nxKwWAY4wqdl08xAO9lFl1y0GXFdMBI0YEs
dFtqwF8trq51jPKfB2o0Pjk4Iw2mmemtinfZne32zYvAl9fsz15Mh3LAmr0i
tKH/1EnpXaZXGTwnos6hg+vfh4PaDVdAaVdgbqJlPcymEFve/E2h/NulNsN1
gdyrYLRshqhWeLZbALLVfXazCgq6MRA401K7meE4Q2Bwz9bPHjPRlkI7EoI5
Y9I6qPDg7XYg1H3BNYYMcvCv5PtbYfOotr4Hxw4jEjWK989JT8sXu7MGonKp
nUrHSVJvbXQ7HVZl9CFJyWIhk9XKde0Laxn4Xpwkd0Ot2gvnxfNst6a1ivMG
VIwnPY2xQV5EtaVWOjm/ZIHZw+FEPQCP0CX4YA5niCKbH3NMH0F+pjlMOfjs
vJF1ptg5qwwmfaCXf9m8FtONUZS2qEEp4mXNKPELupBpxghkW0Vtb/I39hth
cRpOiLbipfbG9fDHvNNO6pHgfa6aywlcc5gjuwM8+v6+/n1mSV9VfVTEzKbC
XXk1GPPAUSggIjLiJGp6GblmhU+3dERQVKPKEzxQlugelfm0rHC+nhavM+KO
w76TeDpYkQP9xsn3j7TTg6dDEhQoVDY9MhfIm89dop4pXDX/EsArfIe8YfDx
KaqdgGZhQbpszWYqFSz4hikO8eapuOvgpPw+L1+gvhhu6dUs8MrsZW7yxy0Y
49U+OL0+2/m2hABidOUGZaEUo77l/3RasfUwBTzVmC2fZ9lgHulySErnNM1f
UiablfFat8P6n8CQXuS2Xu6/T3+148SH1ZiAq+Myh6mKOT3TMvW6T2xGV8BV
qi6/ZfggSZLgGyz7KsrxUrGeQRa1Pp6QfTWsLWkjviUoEHOcDHoEqRO0eKJ9
4vO45/TeJ/+lgUNiCcj2TUEP7B7MzWhyR4cVCARPRgrBUvBNOaKZRWK4nJ9+
34Cm1UVMQlicnr69HDDHF48fD+KwxObbfBv4N1bRR3+kJzFfFvjW1/2zA9sh
cKLS+h+9O3JbGxBCreTVopYcnJwgDOqtI7NiNW15fCE4l4Gylz/lMJy0VsJ0
TS74VniTEl+AA4HGxk5eCSTC/p/v0qA1yDFHlt7ZZm8tRFDGq+hVhAouW8HT
9ET/7YiFNOJylR2XU99YmkiNimQiNMF7fNlBeshyUEaB94ZmmRAOJbqbiP0+
RvUsPPHvrvMd+eGdmeXssynx4coFsjjZ08Py3VEnc5C55HSegw5Kv0YGMfmF
GRQoiZf7yedhQ6WiNJhtWODQeuAU/ZvF/QUVqVFCrkeTChNs3Xc7m5yKgCfT
LYRaZFhpuGdygRKrPCjRhswfp4VmIJW2hd+j1ijPVSBVd30QIoRKR+vOCGgR
GlJBvj84XGEmWpLX8EomTCZ5JfxJomjY/W4xAQcdccL5qt+1VmmdSZoJUiEC
D3+m1UGsOydhXVA573hL+hBCKnQlmq/Mcpi/3q5hwH1ViPs8Uys2JaMZuH15
HWFXfgDrKiGTQVA5rbShmo1cl0U899VfrhlB4Ho8wfp1BhOnB8ilQAzhE8uy
ML4ot9r8R6ngyyltIFeD6aIOavzrTq5gl0innsnITG7ccJ3Iwj47mxv12A1D
WsV2svvvEzvj2iQHA5MpDDf54ZhCpzXjQ5dFguH3AGmFNk88NxTwT78K8ZpS
ECxwecJ+g2gbSg92DaltheKKOUtel8SOwuh5UsqJhgtDcD8lsmIXqJG1zHmL
fi/32cjLz1UHelWSmnt4M7HbaqEOL/WM+QCLtraMeY3LHkjM5NuwKk7TFYQ6
PD4sLfMjm3lm1J0XBEIDKMyt7esYBJNJMdtdTBC/NKSnLQXp/oPkJ5glhQU3
RJYS5FBqZ0aC3izMc3s6lqzLRZ5WU7uPtSmEKNVrxXsA9jRXNk/LRQsNkNg/
qORz/Sf4Tb+JP1/AEjoEl2Q7zQFwlL52m01MvZY3x297gtbLAEA/q4Rvuce2
Vk92r0bDp04Mf3AcEUQfB3uGDOl6+y6L3f8rFOf9pwee18HhDcXmbzCSXDIU
2NNeid5R2EtONT3c5CRxK8YcKe+eGYngPNNGpyR43GY9J1OytZ1cySqe+NMW
p8Wc4YcSDxJsPPnJvii3G+p5ill3JxYB5qDNHIFCRTvYNGqSV3uOCHnEl0DS
d3JEz4B3pGlHdK4tWvGGD+ajbbOSEOiOT4XUD/HBm+x5I8jIR4O0RILt/Nco
BhIHIeHJkkvQ0bpVbNrJtRjU6936UurrrfcDLVdxJQakMStyU80nwwvzXfPk
hd8fGLMh1ieF2x63FarV54QttCAMsQZRf4Yd4zda4JgsxSXt3swNp+8VYAMR
ETXUjMZS5auxI/Wr/q36BgBEG7FoFyb0/srWzKttqFjepk7ASYSk2DTP9AjQ
Ykb4dvIBuQJ68tdWw15POxaURDUBFbe8pgItENsdkU9M7JsEWk4nZdo7r1Ch
q4a+QpHo1j0WffqT06771C+l+rKyFHHbyHT51mswveiloocwargrojeg0kw3
eCI7rs9Pxiv8j+7CkUhWYiTPNSbH+YX46Oc4NoJbVtlGxd6fcIFdXCV85ACL
sKQMgkbW6v4skQ0uLZQEZGQaVY3Nrhe0+pkTSdbP5yDDD3BWBSg5pIGGbcJw
iQIsxP9BU2FEb86/sSoD/7uGKEag8HAuyTOVlYKSbICIz1r7gMqrH6FNbpfA
tBIZS1Il/dR2DiYyLnC5BySPS1spM57okS4CUy82VFF0b9gknz04Z8gH8vvO
Oe5U3oYv1t1TK711UkGP9wQLUwA6S5Mnmfcg0dY2ZKC2vjYQsPcF/n3Smjzg
eh4RjTQaFo+jWprtYF5yfwpWL7GK74oodgf+Y4N5XzrmJWbvBCUxQyA7nn+A
igfKqsgjM0geRYECuuZW/BmN3KWhfgPTl3Wc309b+gay52x8E3yjHP3BmYvH
WWX5kTes746XmX9s7zFjatWDPs5qJkWDfWPF7EDs55UCax+94H6dl3Abw6Ku
JCiCWYVIoZ0BRU7y2+LSSCTP9b5zH+IK5Ar+fwG/aoKqcuuDGfJDMkTlPPD2
wVcT4qnWUxIDw6XGAJqz96Fl3KGKihU+bgl/8vbrb+xw5ayFiFtsTl2WoN67
57/dAajt8HNkEupjxQN3Plf0sfzQFDgvXhEaAkd+Xh7Sjs2zQ8YY6w7LP/eB
bddrWWsIFIpIdZnoquH4vfvKKL5SXCrHdBeSdL6q8Gcwmjp0zZgQA8Gj3DmV
e/eURruFg97eQacHatKD1lkCE1CDtcE0O87mBeaGmjKeQxSXnGFiPeNHLGN6
9EtkY/HzMalusIkdBT/0UwCIcJJJ1cfkIqA9qlBPDk9LqYvs68HI2tDRqCk0
jIHjWWMyxxQaam6aO/EmOJdxOLXQ33dJzM8YmYWmvlNpeHJpPHC0cIwTgtpl
2w9Ewzl5Lf5uCOkprrWH28A9VRQVtXRwK9ud/wr/gbEUwJRjely38Onh5m6n
YAvF+l9MFxWkaHFYfhkS1NbIMSvSXJtZfkMNbndxuDGt/hfMy9Wd6Li1SPCK
9ERiZTYGpao5FPIagHWlhN0peiUuQNjjuvnmZ+GJ0XLjWP5NaurTncg1qOwi
dNHQYHlnzTc7/Fs0uM/ebuIKzDobT07C5z96PIVXgsMMvAODcsB90YptkEr0
mkfrQgqoMgNHCL+5dgxeooo2APgZvi6spGoJCgjkMpnq4pkdCiaDla9Kz0/0
1ddOB6BYwoX5boVzuch8zPno/UGW++gHu5boyjr64QOMXAoW4RVr2C3XLKpr
71P0h4tpSnn7FBwnIq4LISdjXbh4igcYcUhH8c67o8Q/M+mmFSvC9WVXcSJk
Oo9Pc4DNmAu7lkJ2Q+jnGQDuXZuuhHxYx56rTRstJ+PZShnfBgQbCnP8PPxT
R2j9XrJ62fK/f8ZaouPme5wA9PVA2i6AJB5gGxLvjKnjpWhrZbSRPve5Hz97
HQAyK7aUCdyw3D81k4bigo7Rn2y35q3NBixnCovGIwlXt8NgOBGvUBcAfj9n
XS92Dh67s2w2lZtwKaPm48idPTZtH4TgXa+ClyQ/IH+pRt1HFwT519fDRjcT
M94LB32dWG4sjkkBPbxbo7U6XZAfH7EB+yL6Dxqvivb63IGLx84NIGkE00o8
vxp2VzdOHTw/NT5HFgEyVcZv2aDYKyXQSKI/KJxLZQ4SWcJvqhhm+PCO9WF8
RDirrEDLsAXXAh1h03SKVF4PxDvK2BQ5RdgttvJcOeesDCclF39rR6JBmC47
US/IZUEi9qvM9TKMvJxoLrMSjpwM/C5FPkHVTFxWBIvZDRKMiITeDFkC4+QJ
rkB3XffjAsIVnUszNRHib2mhP8bXgXx6DeM/CFzOEUM3B9jp2fFzE+aFXNxZ
13ZaV1PISkiwWJ5Ay/P3mN2VmOGbfGRFX2RvjejzTzjpvTg36ErrpR5znAcF
y+jZjV/yTm5/TeSFlLIsM8Cfvq0zvG4r5RdeO0/sIVn87ml8iFJ4E6M8nkj7
Xje7FNfqTxNSBL4Wjx8TXIbteY++54T/q0g1TJU0BwQb+F6KZXgAmFLqDsNL
QZ9wlkbZEmHBfoJHKjtIbQNtigK6+tAaBQUBRLyjQqaJSDecyFUa5VYijVOK
4s5Habc8ifoPSYHcislXyKrIYlbKR48GW1nNp3llaUV7mo+ayIi9hPH26UPR
yAdrZbHxkyP0uW4C3nQJIvaCCJte2rBx3+orUXAPJrO/6vOH0/FixPmDnFvd
HPYHz6topKaN9rMy7K929sDAJu/QX+Kpj99kEKnt2ebEdqK6lv3UlV+4kZzU
jybR+gJdnZx97hD2H4rDsbD0/jdn+BY71CCsjugoPjuHaA0gssEDwSE0GWcp
nESuc5QES8wbtgxrenaARnaJXIjZ0xkMydGZH1GgdfeLiSdyEl5l9Pc8y9R7
H7uL8phnD7oI5yFCVo6rzyisD83CGL6Gr7Uu5y/EjSe7CEbH4wYjgzzMKMx6
t3nytsHF8R2XBvipqVhXHBDEDk4yk8CFf6SOV37akpCvzpggOaQxevoxrlj5
Dj/ukkuUJzC43eqX2RcVWnHZg2QHlm+7ExWkwBd19qwGeg4rpT4oTxGoj56c
QI1VHNCe5ipobfcdGH4fG+EixMhGsUX4+T3STP4hYF+k6gcrzNs4Gq4dyXBx
uQ2tMncORQ+plQ8m4LbeapfEavxHU3/yMcilnR8ONC4L1K3AkNSq1ptdQRAs
xaE7zSEb64gpKLCC1zWk3RC/bnXpYgycMDllsUovcErJFk+iR15dM7w8e8vH
8FRA8Wu22xqu918OlRXl0tUHgJovXG6KeQLkVahu2PZHrgVfUBwG4KYSC2g9
uXPLAKX7keq4lhs7Hd0qF0skS2+ceKIXc6fxPr018fhvat+HpGjrAFW/x265
B/v+xcHmzFeMG6s/NhAOWMG923mTK307gD6pCYAEqSFnSYODu/dclirrvhkZ
R8ZTPgiGJHwByzk1gzIFN8roZXazMtfnXyrHcfsfdxTYMfMFxAwp3WS7zWC9
GQNllGpODcCpy8p5hZ7QTCUCA7W5Tub+y4BViCZ4TAhZSq+CN1BIhj1x3RK5
R8lshj9nKHsgDTK6bVKYuejtgER9fKc8Q2H2ozuseAQrCwU8JikNfUcY46vB
slbq4LXw+huunsyjtAF2/q44WYaSlw2OWAcpp4iMFMBqkA5ggKJO8TSfddFg
mOD7/zO46qks0QhWFNuXwwIYcMixkBWwz2YApQCD2fo0Oen+HgDRNBHx1FbK
kyw0VUhxhSi9BTYgAE4pY8mgeYvoSvOj1zoVFZ6KfHh9hRwuODIyyu+w7VnU
s99pgpooSox6yCjXzWVasNydPawg0r1kzJ4lmOsytU2eGkddQmqghfmVhLT9
Hg1HzkkVYm0tbj1MYz5LoRxf5Z+HdDd4flgmtEVOgF/54nOxR7tf47FMHx+j
uM4BoxFtul6SW00o7l9jhrVzjYI41GHWlnMgvg/EVHPbXIgY3PrYMr+Iu/l6
6xd+hW0INcL1ll1NG+QwsIojCm3bYhaAASJhXlJ0NB9ysVvSI8EZ5QUzzUz3
270YXM2WfINZEeV6yXzDoWuvzArO+nCxD5cHcbD05Umwl0eXf9QLmJWzKbi7
1YErU13zFMzslDaOQEuCE6nVpD8PMXYv42hgjv96xm0z6ytzJGwFH119FFQl
v2OmVRxgPdJoEfl6LxHGsPjfkm37teAI0Ywe73/k9fQ/FXW10P9+MU0p0a40
XB26m5AQrzPIloVxyhp5GiS7W4S8+GqFYDMKlq5JoTwbbbbsZannn78Syly5
Ir3OecB8WVZJJzOxwBT1rk09gHLIH+LFgIllakYpePTP6sEkgcABXDoci25j
LlYwUj8/jNyy39PBJtrFMR9xQFAz9BNv4D9GV1j5wFHcFY5bP8DRYfBQSfI9
05FBlX+IPdlCEhN1gZ1ApqUf5wzP6TLou1kt87iCKLEPyQ+7kJLnKENNaFTl
vv22PAjIPTjfT0bZn73A28KZ4QJwuur9SrvEV3NBe9btKlVly8Y0M8nCOJBY
05lYbgue8GVnnMA4qrmvvtslc0u4jTdUgsLzoIIcNUUItQz1QoTKeG+N+hVf
+FZEH9vdnm/Hew6bNhBPD4Fx7M74lkIcmmeWlLhpjHuRVi0Q3pctfXQkwKUk
rCuT81ieE3W13CXJvL12zTnXqybAz2pJIzpNwi7I/rXcYY7cgZfSLnqvjjZH
PtzLY0ZSLai6Kes3zu5CYPH3JRYq0nwC4xe5CQSI99j28miDdUUYEPSbGBLo
najtwSVuqfUUGsCcXE3xMHmol3ut0aOwx6cYwFHnEd/xtboL/vrGN3MolADS
kZYVcsKlN9g3oOWddXVYN/M9Xhsqn5qdZJQe8gCgAz3CizhRkn4bf2NBNGPn
iYg/U03h1FZvexql1gylk3TrtvbEyyCbCmlPS3uLeD2OHmHRF9v7DHdpkE3r
VU1OqIqyPheZUI3gwZw3YsEtql1lAfhm4+U2Ktc275SXgCpVMEP1TDPDG6Z6
lj6Zjlw6RJb4hEvv1DgRZene7dvcm8NypnSZ4dcZIIUlV0Cb7wifEh4pjN+u
cvlGWdMhinTTIfoskL4rv3ZokWKnQgW51k6/88KweO4IhDCti5+XRimIHRLh
DzOoXdG4LDIL7EQSAKKNrdbe6rmFl+Vl8yvSHKQmjdDTm9XIFO+qxtd2cJ46
tr8a4YFAlRV+/wYPRshrLxRtpFvnajDx7VbYClsgzR3tox1qHKOLTtAN317f
E2trVAbu2A3oFr70dCYOiid23pyo1555liX0iT+4gW7Gd/oyF4o+gxfYTLAX
zUGUjvEpbXm8DQdmMwbMvWaSiJVCGxuubyUKRqPEq7wGEt3rkSMzp1LA+m7v
/g9kdDlJGkyXOvqupRrk/06b82UbePCx1W1BtfvkKZDubpVsVAppQ4nQqyuI
ke13ln8IFsueBgjUFbdXjXyGYM/ZDd1E1wAJfj7Bkx99KnezJogBSzTkI0Ry
ap1wfHUYHEhqI3r9HikNGm6oqLcZKCrU+hesZQgEJ6hZclgTxR3wbFSBwEIk
Nht5zXNrf2ujJHhggW5f7GIJgMvzA4yHr9ahGL+nYVblAHThfvZgmx8nB1nv
nb+Q5SClOwcJEoXjvvJTKO0zAZZx9qKM1y/ha/9saKeSYBlE0WKaeQFeW00N
j9B1W2Mqiod0W+nx3RiIYaj3aMWl6q5bzQ4g242TB9/LSowmQhgPs+MhjNyl
LtQisSuxGV/JG4+Vl1th74tvZCbUq081SZ16onwhSNEa4J3Q2+NYNocv30Kk
lPJWjfW7b9XQ+/Rz0z5saThzcPNgQs8bjOM08yEl0zfaPyVZbmjL9FXlAJjL
Lf/f6Rk2p98v4d9WSXoik1te+7bH4QTDOvJpuhw0MRwWT/y87Mb67Um24e4E
3+7TQPRoYGqAfkon6btVnM2o1ohhKmv/cdLn+lbY/vjOGrzxoFMGvj2gF3Rc
fw0wawo2rDHEVHEwAi/X+7lAvZMSccPzz01V5VSOMqvYL4olBeHMaDx4ke3c
NZ1+8M313L+awvLvUkSXMW4V0spIKR3phoxvV0JgAmQuBs6mbAOVkT6BtVBQ
fU4zGGIx7DBgamLaFXNXNjMUVNRelMMx8mW1KJfusvvN86ZKgW6cA0v5JVIZ
wa3xtglA9MA3nwT3kE42UbvAYQGcOA9gQWvFjL0sQ/eUK2kCsAySmei0uc8a
pH9xtlopG2vcGcvqDoi15V858PiY1Lxd6Y/PvHuUmLpDmpbCocP4nejw+MV9
oE+wI/MqB57i1QE7y1tvbxSMWKnOAHuBAutL61k9uXED2JTZwJ/KEtgNNs6t
LuTuvRLJQTqWUgxcEJ015wf+mkKHdpGky4j7Li9pQHaHc5FkaPtY0kx9rBDr
PazXpodYOzXtcX7JEUgVSFjhmuOKwCDyi38j2PGDjSwbUOrTt0g5Dpk7sbNJ
53fiHC/tgA4C90+nknyMJGLw6dl6OVrh7ah0aYkWlh8gTOGl1vjGucG6bZ20
hBenFpHiAgw/yalvsDywUSoGXfPvrR2AiQAN20f6GtFTF5FgusJ2zfD6fIuW
JL8VrIwSU35ppdyy4g/eS4s2SQgYtB/6Ou60FFfgKAEQjNsUAAktKFcKJPp5
h8c5mdPKPGQE7P4KaM9jDpe7+j1dpT2+O6Uv+JjxmJDiCTZIgbJCTubr+fzh
HrekTVi1mhvCeH2vN8X7+VlFf4eDtZ9Zfdt77ycktsFM+X0Dvi41iYqWphxu
zjPYPL3y+YR8Ksu7p5HshGeJfk7CqQHEuFX/KMqMRl9B9RNrHL1i4n4xwnLG
1dPTi1/x6LtS1rO/bfvymVf6KNZGXKt05sJukV9q7I0RDGK6H3YxbKIDgdgc
la+RZz6i/PS+KRR/t2InK05fDa/JOuRMX1DMEJ9/yDHUrWl1ssmkMK+JEVeM
OHcXH79d6E6czKQZu/SPyIGtUhyMGDtYztgTXGGGCMpgZuWa+9w1wh7Nqo8p
l3eoHtZfiMHXyQljYp8VG7V/0kJpuGgave2HVRdU5Hjt+9cabKqHY49lilPy
K3cmjxA9E/2ke88c01L4J1ADIdFPURi5fJ16U8jWvYioKDQTs+PbdPoLN45g
s7aAh0wunCaSV+5oS6V46DFlrsbaxBzRReKBKmOjOum0PZmGx6Fv3pDFmF5n
Bjx2HFGtnqvWtgnCoTEWiMFgvW8G9l+YedKON8Vr9sZZN+7cOpK7ohdkWRJc
7ZGJTuwXJJrlxyoDa13tqIwPqwaRv8k9dk5MkzFVP/TwchaXmkqVVzqDDU3u
zapQ8FCPjLEbDQ0324msQx92aMHQFuJ1t1LRuQimKvNvRXZXuQ0MH5DQ8/sr
5m9+TGUU/kRoQUEC6XfxzA5UHuD7pR+6zXsRgd4dwynkDyjEDVQa0rpm3GAi
Zk5mxxt7Qja56+tOsnvp7qMwg9ag1C84zSQWD37T/MHIsQ5EPFp1Nhdkg4/v
U4MN2CsUuXqrJOVTY5gyY2uppA6FBzJIDc6dZ4G3WjFdFulkm/42rfeiFtDR
buXub8ajaB/PhpIOsmu2VZuaH3kRfvHmAa0V/20kaj1KZXGO4B28e3zvX0Uh
N/X7zBG8xzQB/qGYiMlJ2ry9RZqb91cnS8MC7OPOpA7XyfF8wZVfODQNdCsF
atnWnUCRkiYge20TdaLbPEl0vysA6z/BlhaU6K2EdyS+Tj2XlNN0ZoTivHrY
oxRIwIOVU1jojY3xnAO/oak9CzXit6DHTM97jvW5tmvHaCGYiiFx3vSRQqeK
454DI2NrU07E4fHEpDxHf8PmInVOYPFh/cC/nS9aVixg1OGFJJcmN+LQ0cOC
JHAvanxD38cLHej6w64w9AwBmkKl7PF2Jr1A6rUCYSfkWyYdw4PIIjTPE7j/
Wftk9LJdLyyB1gf4prlBZMPkXz3n4gATEBdldgQWoTGz3JadpdGg0Otdnfr+
acDQ3NtWsw6urSI0hX5qUuFynzIjVPvkcCqLWGVDvbtIK+aO9FXzeAqi0sQr
EShzABQRDTDu91jnPprS0yuNFfjRr+j9HSXr4sOMlrw157LUKV/Ikqhr5eJQ
rJDtWX1uGgQ/w6Ndc4QLWtVVzxOc9ovZ8Hf8uPyKNsZFEEZnXzDW2ow7JOCC
oW9enCanaUHNOEOb5xtxg680iWLe/11GhadffGoNOqMGionZrKMCifB+l+pI
wMa9w+vK3fpjZGIQ17Y7LeWCSlna/56Eer+Sg8M1FRBAv84/WBvkFvaw2RZ0
ZGtpt/eQr3VOkQlyxaZRbqAV7SoSMVfpcZtcTtY7EjdvEC7Y1vY1M26zy7dA
0oA1izzI2D69G3gZ7k7k+h2VOEyzTQ4JU5BPzguIhjSpNi9Kazghg1jAoM6Y
DMfBWLxnhB1pM6RwBKzp6APIxEzq3zZSurF8cDeqFCqqTvI0vQ+My9iG797V
v/4qKwJLngSMcUmhemRtLbiDC2auDo6ehVLcic2/BAAtfx3J8m3c9cYg5D+7
NBg8Zrd540JexVZxMipZNAK9f6esfBOrN1nu78ZoxjB8krE08TI6Bz1NbiQX
zWt4JQ4SeB13SD7DM82PntICJE+tn9937uuwGk/EWnDb7ssKHzG3E43kJl8R
OzIK0hGbBgSIZ0nkRflbUipQU3E1AAYQBc3ebI7ke+80oMCGRJe0SY2ws9ZO
QWwoxcLPM0yrIzK8dzzGktnNihtUlcHahA6vSQF+RJSgvOtmI1o9LZglUU7R
MlJw83WZZ6VZtfsuKmG9dXeoGGuPm8qBkT6ZJfqKptldeKUMjvBYbcwQGw5T
CQ7TB8kItzQQCmZeW04MiH057KWLNpQvBMkPdltNmwotlT2dt6BQaZS1Qwgs
Q2ExEuFXHzEtUqifSHyGNPMiBSrMTp6zkFbPpIyZUB06P828V4IfVm569o3R
N2LEEuKc/Liq7ixeFm4N0avkA1Q8tehWz+ScEsiPdsUsbdAnpnVibVNtfRnN
0VyRWZAQpqlY5vcWN0/xz1Jh+P+X8p9M2hC7Jk5FWuZPg5DwwbfZVMS7Ev8V
ofWR+b+PozTXAnPb4wOrq5mMUQkQPE2jisSeY/Cp+DUI0yA6brxEMLlN8F4z
bjB/YCChItRsq0LH4u0CS1HwDAC6wnrJX1ZZTfqa5MDCXiilgLNlXS+TxF22
N6c7LnI5t0gnXnZfr13j6YdXS7cFJKsbAbfKEubHdJksHPcUVl35AQHWa/PU
/A7GbxJSrEBXXegsvbPp1fHq7rSy8k1KuIzki8A8LzoqiUJt0ZgeukUIqZUV
F6mTISHC9yWPCRjJ3LJCCKrGN/Z+fDjnNp0WXzYnsjnBwNi+JPQIsPvpj7Dw
p0zSKWJ+bYkCxr7ZZayIg1xNQMAMm9R7lSRD+roQ5EJKK0Wy6fe8WYEAdCri
dlXMsQZM5RMz+0NdugWImvEDzCcDZDY1c70sEowbdfJ8j/MFMkUVhToCfg0I
hmR4ZfAfgxzVu2MObQZRyiIDoSTJG0orcukH3AGvotB6zW8DiA9YWD5S1H2j
bl7LvQs/7mIEU0745QYytdo7h5RchVnN+KaSmQ/YYe32ulnEbiwWcJ0Qyhd2
5Nl/igiAtzjNm+WITncLul28Q+Cz2giYn7HVwEcJk2J9lM4hRX3CPsonT5j7
50gsVqZcaX/flAjGnph+6ZIwit6n9nkyARQAgrzJgni4mbbP4JMg4GAjQ9FQ
HNzdrdBxdipULe6jkmYKAVRA+cTe6LsJkbshIVdAIkCTYTfaPEVMv/kE4MGf
RgGXLSyZ/ZwZS0lE7p+RPmQDNEypFETE63tgcmUveelFeoPRKG+eQmLE5KDI
qOWnyYVo1tKM9m4wueVvm45bU6qhlKqPQtA7n4bcLsH1CYqiCyG3mxatUSNR
VUlZ0nhTwgKlw4euBziduzSMgP9NZ9U90MiUhIVl/fMsRUzWWxhIpPP75zRt
BJ/KC3RE/+zA2Ze4JGfF/C/uYk3R0RuxzyBn0b+8TxVZJKoDBAZe5x82lpwi
+g2zQ7Z3573LXFuLjrW5nKVvCmBrHgeDixdHO0Z+r6eYMhEf+3J0Sjw5hKbY
gth1TuT6W5oZc2JexMspc9keN+mOFXzD/hdHVamioJvqMfWpaG/OgqKvqAgw
RY9StPzwoP9PBKx5+znb+C2XZQFGUSZ2LanR3/eMEj3SmmCXtpsVxG80zCI8
dL0Mf2tQ2Yy8H6v18HIl922+b6/LiwZcF+9ZUPtOpQIWlHStCUbKEfKVluxB
InuBb0JHZ5eO4u0keieVYpXE9/6Rl1JYlTQm0GJcqfB8QBn2nWH82lZyfIzj
lyIswlY5DlV1fZS/If2BOC/NJV8dNIde7KhckZZHVYe+9PMO17LuPPZk3drq
UIMl3THEZ1IgLm2mxYaysVH4j9KsKUorRZaarAAyQ+Y60SEoDRzWqA7BnVI+
N4NbBRjEG8CvEdk9PMUGQfMNmk5YptAU0yddJXWY1sqv+UysrCK19mat18Xn
Vht9K/mwjHg2VKIigODhm3H2DqzllokApo3gzAYMwv/jRP9+l1DDnQcMVVAZ
Sq418kSZJmavYPQg4iklExR8TK/8bGXRktiYtzDdCZkCLtep0s57+IqDVaOR
Ze1OzQWIGu+kVOTandY0922uu17U42IRkNnMU0psv5/CXz6+PVYXDWBqyp8Z
3Yyr4l9GCkKQ2HNh0b4XJfFf8FKQT2QfIhaNsqyawZ2aVDl1CUBn8dA+W7J9
xm/7NXglKQ4Il38vufCI5so6fC+9y18z0zbtgCP9WtGY+qgQQfPR4g72v8L6
Je16UVX4IVIyxftyQ0ORQMQ5TzQhfZNbaSt7EN1L1K+OVAKMCOIOcU0pM38+
84uVQT5CieQnqIzFdupSxCdxqqACxpEXz0tnJvgz5P9NHZCwdMry0KNQyjCn
dMtwaj3EypsXwQDks6q3INWC8f7dNwp4dZmBnxILgm3nOE2oJZThBtHvX9vq
zVHo+EiB0MdHDjIqWQCk8uZ8iZ8Jx2mymuHgFL9AwpLy4pOFQqL2pYlNUYFl
bDCG6d867TDjgSh9oUhnMavaitb63lVLMBGK3SM/FSto19f2/BBZpQpbG1W6
vF4frU2z4YwdRl37XACcPD0sfLNAjkbf/x1cRJ1f3n3UAEmfldnOPYepM3lE
XKghP96K7yMPkxj8u0kZpf2dK0rv5ziOrHTDE4RTUIIDwKvxlp9K27yTnzbP
hGsToYoiBFHSNFHOTImtziTKVO9roYuo6XJ5wt2WwYzZDtJEZGk/7tBMvJvK
tvpDbGfVWYQly1ItR3rMKWdTl0xHDIBZlLRsAyfEQCww30tbUxzBOwLBTLv5
q05Ik6ZKBi+vjm903pM+uyCFqB7/LuhFBe+D0E8FC0zgff3kB3c9uJVzCEQ8
wGrL8qYb5WL5eXG/GWtc2IdRRFPTTlV+X0NAcBjqChTxDj/L+xBuKqbLJynW
UtSUGL/tRO3i3EYs9eWrQFSLyhAmCao+hXBo2tkHpqsALs4jmlQHf+z7YGsw
7jaqmnUmL4jdOmLt5TQlgwDllBxwndrQPvjBlmtxhR9lp6mTG2SCh9Oz3s1o
l0fUCtyj+OV7PEtxJSrwy+rD9Jg5R7s8Oj59eM3O4mYwaA0T3Y8O4VwmmfDS
Wqoq9z7ktXzp+LbOxZhq00NxueyOI/FCA8m+3rasUx5328QHw0ehKKQinYDI
ln21Xi1wNhkZccHa7z5SGu0aUwJ47R6HEDk0H+gHID65uafGiu3vB8KY3+d+
Ft9JtJJ3FYtlqjmCJJtFT9IbHc2q1aiZuwYBZCi3JgDZPc0ObM2jEvYKSevX
/uD1aS0EkzWZSPlbaeFwQAQOqhnLqNKe84ef8hocC+EpE3Detbop8njg7AL7
DDSsH1YWsN5o4syW37ElO+1R+dKLENaAaZ6cd/vzffBifK2iVDLpoALWDLxO
PtqPDnGZkF5Qbsb7zSlvvmyL4EZc0Z2iuXSrhgcatUulwUJT8Y3UhN8oP8fn
gX3LEyo7ylRoAOzUPfZToVmLa8XADmSgtUwEZyP9ER0WS41VUTl6+23G9TqJ
01mKCzqM1avvspD1YNlf8hTvqvGPFNhe0ULW+qvxUCZaAvdJzQKgXnZMs13A
OcPb9U5/hAwGFr3aSdsDdbQEvn5BXAAHggBx3DKwuMqAPDmdPkBxZY5P5MT5
QajqInQ6dU7xHWb8vK/0wlQzyh0PyJuEgo3EeA4IQGCuFiMjE+zaRaLH3N2o
+k/Ow6Ljl8ZU9n8erDgj3dI54CS7BGUVppW3vnwsgTQxaBjOwgHz1rmNXF14
NjL9mCIfJZHISaklyLzxl1wOGdypS56lCGh7KcEUkYr4fVpwxrrzkXAIdr4e
4yojBR+R1xcaCccYp8yaD8Qhee4YB8O/zXoSxT2H+lb3Gi8CNJJ2D+lq3TT4
3V28fZHhK94trsq0cQ+fItHpESZQCiistdH/WClwulNk4zswquGBwMtnLRRG
ADpl6HPCuSLET7KK9W6CDYc71T+KTy9zcS7su/dzdv5PltsGPMzNVsaY8p0T
JiXYq0HNUdXlPxQEMGhb0eZvUTn8eSDYuB+gF+BQvTxOw67XNavh32GC+L07
Gixw49FfsX+Bunz+4Q3z1Clx+3fddUr68L39OaO9uWKaLrEl5P9B1sfZSriv
O/UOKGEDF5zMutcaNxo+hq/ixdcQJ+vWcIsIbmoexw0dV2sEOmzkr5gtegQF
bdtN1QVJfeioj7AHF2igGAONfpFhSHkynHO/SjSrw54FvsUUU+kkFEyLaYRr
o3v3ONbPzIQQz0Ndg17PGj8KN/jPSBHHOIeon+LtBdg1zEEKZtaAvp/RVukh
rpGa+o7UHbYqkh7Zl/Kvak3rk6Wpy5hr7Rz96BXjjIYkJH/Q6Ib+UOuMbdCJ
pk0J9KbR2EF3v72uZtA5deeJBF4sVlefVPicNJYlhfzypisX32p0f+GwA5yi
NaOWucayYkEDEnQU2vl9tCRGlR8LgFryY2ZXGuq4uRfnIrSMYBFrGrNmQ+6e
aQzfFOYVsT945tqHu90zBFKb0q31T/0uevRxKlutliy40ptMA/jXDyOct0lx
8GvbA2rxmGcJ6aK0/YNDeME8PTSDWnsdlYR0wHeooefj2P1vtydK8TnxZ8WG
efzBBVwOCQxWLIO+aXVXvb/7+blaP5qzT0HweOpWOk2naXZ8EtzZeLEhaTgv
J7xFCZVBCPvLoJrGA1Ik1RFKQpGs7FFheNiHHpXdc15xQ6+upugkxkINQmBu
gavPerLwbfwape9GcCJrym8h+v680bdAX+L/tToLG81xDCbeh/f4SL5XMKgk
sEG2cs3KSi+aobXV/2DpOt8Zie3Zufw2fAx4SfyBfosxiwmyQPCTATG4+S5b
zDeLaoJ7fr0bU0+14GBI9zfgrrxEykV9H1+TuwjDW+fxiJ1b6Xq29d62voul
2pNxGSrDHUiF4PSCL7lxDXp38jNh5joqCwBCTBP9yIuH+c4gZq8nI3KpGl2y
/bZ3Dxg/BQJdswmTNqimMlu+P8RcfyA6erh9mOwAJfdRPKR793uqfpdfsjCs
Ir09nWk749c3Ui9w8tnTKuyQ4VN1UyoON/CHReNZ4ByBZVVYmDjDUaBcFhNj
VxDt+xQjetEHiRL6lcGaQnsfwqHwJz4/LZirr7OtNJIrUQYUzubvhCeOMYHo
fke+PWJgLPg9oqda7pN5e1y79PUHtgZ9kNHeDuzN5wDs712MxmRlC+FfIV++
Cprzk3UehyrTKvt2wmeZNIrGS02EJsa2Wk+D9uch5AzctpzpNafYZSTs1G0w
kBI95Z+gU5CVgvZzbZC9QLZ+5xO2FBxrPGjSf9OF8XPqmEwRn1ccMKQmgnqq
Zlzvi4mhlH2cEOxfXUcoeBHRuWp/+ujqIosSLY1oTCgkeO527P8R+Fbdt8NQ
PVOqsJNxDSNyR7uC0+5gyccS3pIWAauCykKgmpOCHtwaZi92wJxjyKF19Uqa
onSEIkaYqcGruPd23SkpgPpSL5TSYdmxnThxo3faaBTs49+/opQJsQwUlGgg
FEZLdjpT3u79m26G2X8WTRDmPlTc+4OSBetVIJRolWmrzg3QPnEPdvC3kcqM
FqA7EEx/DPJxlB1Bxl7gdko3wx0bOpupjHQ5eEwmqhwtOSyA7b4xCG9kCzOy
qm4xsbCD43udpD/oZrHJbq9GJMMjXD/BVhCihOAO2hMmkv8eidufPzuK8LI5
tLcLUKpFGuwyCOSZBmUQH1TD5iPx4BmqrGMBgvrqWS3EwrQsEfjNGPy/OQ1t
J6JFjVyVbk5ZKQi5x0Hgu8/nQJUmwCMreilUI2qGCrOFldnseBZ2/cfy40UZ
bdQ+1ZHpuxki11PpSW/wxLg0nOaPryu7nuBChTpXrVy14yk0NfsKVpEr6lfI
LkwZz5aEjn+LMRNtJ6jfrTUXrECvV089OfDpDuHbkC0N6uGgDKQjCEQ4iUL6
KsnJ6P5sq7JPXOwDkPE5S8LgbDvnMJEjLQeVUrJRwO+9BzAuuFxYiP0mdqa/
+hgLHGLD3lNwvS+9IyeMUxGVuWTlijAInNXlKJflLjnpIGDdaCsO0v0nOnBV
7U5abtopXR1cojwh+c3NeRwQsWQZs4Tz744NPiBpbbrp3A7yEE+vaI/3UzMY
dYKtAKb3SOI2cztbb9vf/+Pi2waBfj7J4P/jRE9jecLqVcaNja6ANHAhcK8W
CLdlJy4o7HbCWqgLieFeEhy+CTHrQ1bmjA0GE9UM6SSXx1mjQJCF7AK4wAwW
BKJMSh/zD+J/LXAmnPvCnQZChWailIoEbXxHzX5XU+AftqVirPY63cNTZNJp
QhKgZWopKqWT6AxszqIGFQuPGw8ZVf78UEBPGrLZ8p+0LtXwiRqjHBfH7Knk
RjUK/t+PBp+quIu/tvYMx8pf2lCyqm/nIOtrUTCmmfg12rn+Kn8CCrkKklL3
d7EDMnnyTu4k0MHjk8HEBBaS+rWk7Qvhzg12E0CmKvjRsH9UGYJtlVmujJdt
xnnGSpek68MCCinVVR21ObnjyX3TvBz9+ItQO209haXCIl//5PnHjMf+kvqf
JWNnT336phtykPmDE2JQoObjg76uFIFwoV923Qe3Gfg0YecBCIlQPUmpjU4B
KOS/4J8gr1EiRSjY7SiijiYQQAuoXtW1ZutZ8Imk3HCNcto3w7dcTfk2d/HC
ASROpP6++Gr9iDM/5WU9LCz011m4ovxYgOSiHCFY4t+4WfV0eui+aNqY5M84
yRiN0GotV67EbM4OJ/yJfiICRIIi3sSDSss5SUyi83DanRKa9XERqwE0I8Cw
hioBG1548QtPvVJwQLhcF/7cJUh//LCDoU3K8M6B9/Vx0xWgBzmpSvDU+8Wp
okT8KIjeL9HSBVFd3/3v4JDBvzUtgRtIFs1dqPQegyIEcgVyrPRsW/++2fde
rDcgjvA4D3+YkNl8AAa+RX6yEWjCy0Ukpo0t+7cGg2eVUE9AfHet2p8hml6E
+rllim6d51FV5JwYbUInIia87qfWSPMFH808brl+NjTjJvxkm7ef7Dfh7R9T
70yrs1pvO5GWuletduzZDjcH+Xfk5WxfCnlrEMR70W8DIJpDzUSVy6cE3AfO
qjGK2BExuRqUDY622ES1ozD8KUYCB1F6t1TKaa2mThUYFwhIZq0tUtAHyy9/
cFFx5F+aILyk6H1NpCn0qKWwsMfq2J73BFX0UmXB3pTHYP0REQIGy3UJX2wE
xWmCyzP/fFO5VV82O5Mk5n/JUqZkUW5rACMzsQMR6GzJXzmusdUjU3LpeX/T
Hri7G8byMuqyiJo1MibbEkrZsE+MeSIbXVGx9dU2MZJGU+YmbCDvjaq2xmj3
EKIymmN4sytbJzE1eSVwZnDyBZcJmwTSPLmy/4k+Tp3n3skKRZ3jIj1PGtWW
vZPeowZg59KMz4wRZcHej/LYBdmEtknBAEQDFljaiC3wSTqA/Z8AOzd0TylZ
PqGDAtYJesxqJ6LO6di9vyiGWLoKtwz8xQa0FPsyGPMi1HKXEIDRok9spcTG
WmxGGtpocQlMVQTm6letT3PPioa/Q7b9hlg9zZr9dpysIBngy60ptUsCv4Zy
0Gr+MEGxOicQjWSuVPIaH7627Q3q9idDGpGsauLDb5r7d6q0FE37N4F4iDKl
MvUYEt2tTo1+ZiITWs+9AmjORIs3my7u2fyW/ufvAjHmPz8h7mDOb38o61dF
iK8GpI/hzjRaX3Ms4HPhDydmjmEUGHIxT/rQEYfgebtDyVECEWGnxHxxgRMx
AbCCt+ekWiwxSQKy5cFsiRkH5hvQ8HNu8aN4cHyashvILD1n6Fu5f1g94VVX
nSswihhcIFm1rMVckIrvD3vDR3xWGJX903jigZhmh1MFZSj2lLUTRweMrWiS
CGeQdPdGInAYQeGHEuYmWCboo7yKA263tqEJDD3SrA4udjtFfnXzg0wJcr/K
R11Bf9G8oZNSZdNcsRUU+tcIVB08SfVPsU48mb50zxsq4SFay0ON/7nuWR0f
65JlLgqgU/eTwZwTyUrycukeZxg8lIqCP0+AEggLP0eLLzFAv+NBWt6+d+Cd
zNSLk1LbP7QYFxq66CnmlWZJtph13xrI7Sr/NYZn+XhoASwqWKcUD5ixpoeZ
32kxA5aWdOAeSQgk/ryI3JFKOFIInN/uIEY9A2kXmDU+t8nA5UaR6Cb8jcAh
is+1vCvlNs8nJMNUN1zbRXDkvpsogUWYB9KdJMmdqhqilkixnOvG8Q2Pt9ll
EfLvR+TiaQxwn48DXJ5dYVzFrhde4NT6fObjJZ3J/gRI2WtlkwqjhZ289trX
d4fdtY/W3wqrTeNuFlO5OCCi9YN8yMiYn0A7OZ1jwsfeKBtFCs2fPNX8a3CR
+HGl/M4UTVvFBwuk82EU9p3TD8EcYyeO++waRQT9qYfktq5GWdwzuZywMmJS
3X6pvjtdJc4ZuAdVk+5reMrar5jAqoSsjbWSnTWr5YCAa7xv1rWqkXxjeb24
b3YqIL5rKOIr5oTAbJd5Nsk7Yzp1nYbmMiLggL/BlE2RZ9SvHqoFXjIqN7ll
k+fLbcSMvVke833uPEd5+SBWqZoqxCoQu8iU9qR1laGsQNJW0P/aGbmlGjj0
lklIZqbTQaHLRJMmFj9JlWGkBXLj/GsWL5vuEEI0/aMaLfJoHIwawIu3BEiQ
rCgG69jvTlHB0VMbUcD93xTTQRZnmfsV56I2JFaEVqKGASuii9kZDf6AaEIs
BSjmzTRvcrmcjaEc+446s/PdmIRUPLbCy6M1AO5DC2GFW6l90WP4OVf2NcyT
TV678Fp2U4zZpfKRMZHR1irMUv9KhhhXIbmyeBKUN7xL8LmVn2c4QdA59fGV
zAN/l6R7Am7IF5I3BZtrcDQI04TFkkCBvW5qZsxHYAZ7/qKdJrOryuy3FrtU
JtwjXEkgvfRQrCKIrE5PkWVTWBRrN/oqxuGhUw9RTYaBTFMGDtAzOOwvHH5z
JWC87dsmcP7yC5xkzqmJTMiK3X8e6qvZ6Ga5B5yqmOGxVBX3o0yu0/O0XptU
E1TnABPCwQz+zrQR+zi9kNqsqX8/hkJ6TadmGEg9L3S0Ufq3MK/4kuBGFxXt
+ej9gLDl+TRda2SxhaWVtR/9UPhL0SCjGYPaIX7OKA/HlgeSocPS+mqg2mqW
jLcpk4YzVi8HeHdwudE2omL+dtgEvJWr1dUsUhfWPyJz7eIJO6zcm23XbQmV
QV8KxdcW3SMpPvMTHpUul0qHDt9Ncnoud6MO6KjwBhJqKhKtyxXi6WmG3MEB
fw+ax/5vGcyOqqvjLYacqE2gAoWAHhnkf1EX/an6LpExTw2A32DJkjfr68y/
cR76YtiJrXwhHf0/slTCUD7MPDwnr/QvOgfgEBk586nRI0KejmCuEG5mPEh9
s+NtFYW5XjEdNb6jN5jy5BIzSZlsaOuTlGC/fNAMWyEGureODAN0rbKEd+/F
+1pmrTu28K3VIS7MGwsYxDbpXbouchr6ScFffFjm2Q/dSp8HiuP83WrDDYr9
wIn5Na3SpW0379+Z+DzVZmUl/EoGnXr4KyhN3QI/rbPZ9OY0F/uypCu2Y/2k
MOTMPnicIqHaI+7Lg5qnCHSmZBgwNkhLocZWPWKYpzXnzfspReib79YjYE8N
vpNmzt7VYgf1Y2aa0E9DjvbuJbOxmDsp30slmeL7yb0vaMQ0sNht5bb64vzY
ItZIXzMVQQMuMkDTO8O2rC2PQ8jam3Na7iaghrQjYsSDr62HVPv6ZF7qAL+M
YRGHu9kMx4/jn+BR3GucZPE+2++S5TzHTBcTh5MEjciA3nFnJFCTYIxsbXO8
l6xmgih06G0kKlXyLd1bMHqpq+c5AyDOfggVXmaL8WN0hGkvu3W2uv3RcqRs
fop1A9TcjLjPD6um4yqRLIRggCdCdi61ocwhF23Bjtb6URrvki+kSA07Ib/V
6ks88sa3i1yey/WzWkk3YxoT/nnLhgNmFn3RPomzpI8AWG6Z/w4l3hRCaZrO
OgytG/QHtPNHJfDWA7TYJXZgaWAVELdmh5u8yXA1HSf1VRectj2LKJn6PRx7
KexkrsZguDY8CxSfZjmlKAosVYFjanuP7Trkwsdq8XUYGlIimpPz4o2Kgt/w
pK+VePescZK5rxkAcWikuN32xWmQK4PxPT1BrOBaxuXo5CMhyTZl/1vHaI5z
cP6xwfMvb+CwDRfn40Sxc4/0Q/0jKg3AcYTZ0SXqpRacvOrmrnwBHnGf0TzC
iZedtl22btKEHGb1j+Ue721xCIYPtMEuX+s27li4SWu+zyylAzGGz5IoWKB3
2N13Rm89pKvFEKWCHPtKuZOMul3ICrBOKKEae7BES6c4suNDLQJ00xcZxwsS
Z9c2ojL6FQrl7yb4DSb2kOHmxQuE2bDk2qyV7wxYqaxuY+CQqVmrMyWp+87+
NTuQVZdnnJrEyUDGkBTxOCqKTVUOBAetrT8deKWSYLQCzojl7dVg6uvILNwb
DRjpjayut1qNxGfBvJfWp/PyM4bHybclhdMNToFlNGPqp+fhE5J12f1iSQBq
bDA0JzWxAQWoyhj7Ar/9WLAstW3gE2GjDuim2PyWEpDpd1GqwysznzOxx8/0
PNoYrCRdiZmWko3X3opfkUS+izrQWaS3T2gKCWazYWhbJtos2XPa+BawVPWi
TN0P/UwpgLs9F0eNVLVElZTtdTa6BK9VzFkCZ1yz69BErShHUqLFpjcj1ACT
5rLeEQnqfUok8LsZwxfoUyxotRLFu3RhN6udmmXxqEvoC+kheQfPfzpEkI9z
Pwo14IJsoFSP/kIKpShzSYxxvrm2BzhzA/K6UMZvjkGYpE/BBUM9u5MM1vzB
otY9+NFH4U+OUickNvt80V0ndwwEe0LChpHUySXdsjkrEDDq8dMQoSkgeXHw
rQ797h79Vg9mD22mnWUadbktAOGXkrR7UaOxbvRlmyx7bH+4UIvJPFpp0LLF
iuf7DEc1NM0guR2lEb2mozN+sNK8JVdmqxefXkoLX9AopBETnLQ/t6vC0Sqt
g5k2SxNKdihhMOchTFIaH6EITsHEV6C1yAGJ/sm9Y4HzYfhkm4Z0EXNVax28
dnGqpxSYA8E1mao0ade0fgbElsbyl0iD2VVoc6Kh7zkvQmjNmOoKkmqXOBQB
QYTYK3WarfAWxGa1qvgjWJpqMNk31s2t3S7TyWrlURO1BaGf3gnh81JtjzU3
2HLSYU0nMizateglh33+el4IB/svBMBPFh4eM2gUlYbZr87DkpnfrsRv9kxE
ssQNCJ0UjHb6d1ixGzOt9KcsJ10xHb2q6xh3CLF8eCqluSgf8ObA6a/eajoQ
6VUTxI/EKZrJgft4svk9fFQL897f8B0/9TFT/MNsAltyvHyg9gkbk2ScvWM7
jlIoE4RZ1Th4aiuSW94x2rvLkk5gnGKWWZlRDnSnv+jcF4pm1HRBqowm6G9V
TW/igU6vLqa/iF/LCGcT4m5LEZzE0CorY8S+zrUCSvW6xDD8NF41RrwViRgk
6f1slWs5aPaqoVnU6FhcuZRb9iJ31PveGKRggxKz+gA+7ZK8UxqF1BF9lsbm
bd3ikCxUWUPiVxNgCztZUAwl6rGM2ozEklSjDKB7IJ00Ft8ORG8fg/YvT7T2
TGfG/7EmgKKEzMYaEH4VUuz9G8uxyOU3Mbq3YABBWTwDX8iVi+ZtiZuV4VCT
xfSJtctEDptN8hKACzFQT+Q1sWp6w/pf/HFPPfNrBlE054W7BmbibZGCEjhm
OWzLAq0/5fXYTG4Ylzjk1yBKA88B5+kvwX7JKGlsAprhZJecAA1kBNHxt+xB
OReB5hUyzC1mrS+7bDF+yRPkMospCVxWxUPjNQV7k7s8eWzOuOWujgAKpcu1
Q/xLW32VtDJu69Ct+2/aqOKk/bLmuV1KGBZIZ7cMdnp8nOCSmMGyyafvaXlD
Ztrbl9fvMH6PWy0aXPresqgYRKjbYVaQjdKDwqV54qxXqjVSKPD0dqQV8ef6
xMQcW43eZkAiecLuVc3l00fdO4/Em5niPWufGi8bb9siHUoCiMMpzV3AQ7wA
QJ/aOFy7PPP3eUQVkKdBpVDJXQozc8byQPbvLFC5JFSEo9phBubfeQuOjo1N
HElLWP+A6q8kJ+7XgkCUcBxHFnmrCbChG2mt3KOhn6YClHEZlbiCxwaQRSte
SS4YI+huujBCU8yi7hEuEhRVcOe+IM3giv5NqMP2r8/OM7D2Neq77jk0OXpj
mhDjtAnQscTPzvSn+vR+YCeL0neFRHfyFhAXyGtk79Sgn1UjvVXoadkW87Hj
xGonV7mHfCnr8TXGcoohvoI8duf60XtL1JuNOf8DEoZoowetywq70H42Npui
HPTXEQIETRthVtNyDdt47guyiIcQdp5nF2tyWx4mug/uKS4qBGufQ+r93J0K
v9ifkbl+fla+NvngrhVCIjcD0RAY9ojBdCrnC/kbmFxrC5u/S7q+OvNBs0vS
hQivUtUP/UbBug+fXTLpwXEVZzeRPj3PCsWXepE4SIckmQPXAOIjk4S3LhE3
rfiNXhwHs0sG2Cd1M0iHSv8rO3eSfDKGUgRP1K+a6QowDDKq8UNXltWmGeAg
vm1V3v0Nt0yohK9ni+Cs6URns8BIQEaTk2yOlhHDW8rrOUBKLGIQedy4AE4s
m7eXUJLZM6y8ZKX8P7Vnk80C1QPKFnVa8hy70G/UgudrBkeOID5a5PvnNcXO
8E1POCUr4Sql9uwHqu7KOSPz/4t1mtgsgMDU0q2s9BVpyBYJCuIJifYlIM90
/1d7I2DYK5HzcAWbQobvCURIL8+0XNkuGjvAhHDa65bnhewlRo7O+alk3LhV
GUBTrQjjIVeYSlEENzPu31ydNBdW09iS5YB1H+22ukrpz4jSVNF2uykwThcq
FZrjcVkpMD1ADYEr+3KTizmCxju0hrhKhXeKnZiMCjPw0k07TkZuHG2oo0b7
oMWzkriWt07aIr+ljaWYkpXuSM/SmxtUQF0Dnf/H8KjMJmsU+eqR/fm+Iln+
Mz7p4b7cfDMdMTRYyUqbUI7yqrWQSwBGindUjz3OepekC1XQPFD3VAa2ov4t
SiU8W2I26vQzIGDLB9RDrkS/nq9dEUwGjgUvkjfIzKQ7AQ5GIDxdVtKFBO/9
3hDjXzX5slihJoSCWFMnMYUyNG2AUmpqjAAkJ889nHCIpwfjQes5iriiI11R
2I3FUa95lMnw4jFc+A3BuLMGMMbc2ZTlG3NMmFVrVjuCXpd8wTBPzdljp2QD
oCTNaLHmX2KKyxhCaBcq1wtVIrqV8blN8xiR1btLyssJP9xBq2OG195hFeLL
MjOre7dRO+ROq1H5A861z0NtV2VyCESAWypH22oXj5d23uQz/8HdOgYMh+Uz
ZOwlylZqer/iMgdmTRO1wA/rxPFXzMBka3ErASyDGPO1LHscF7NXIYuEyNvZ
3XiBDtReSOA2pdlrL7NggpRrfYRPXRUfvlQR+HTSa8h7Clo396Bnrkct4FCL
jL/4vuk36m+pCW/wu24Lb01L6720l5L3KNXXeUeiJMEDrU0QvRREjMQH/ON1
7dT5/TVcsdMtGLypwu6+fVE1B7mvyI6i0YT7aI3t3LQfWegUzNdHfl4ntsUG
OCWFBVS6VWaLIDwnIs/8PrOJalXId0LV+xxHRzAzWvR/dA04REtHfmTq6RfP
wycB5LiEOGi0JppoNDM2IpQ9Iae/s5/Kbr1ILDPbOrSJ6xTFTtri+b89tGS0
BaRUHizr7y8L/9j8fwFAtAA3psXLK1FMqh4o7GTSVHxWhXWyR48O1tNak/MU
HAKzQMT/J1ObiR0f/HWmE9nvv+XXG5WBvPBntkkPFE69e4Z7b/ixv1SUwlzC
HcUazmkuWqDV+7YIESv6rckaRkDcyq3NawnXIXtPgjRod6E1SnNTdA9mC4nz
tYVjpW64F8LHilJtLJBmtYfX2FMwHvRxM+y4CUmoWo4VDt8hVkqP8N4olLVN
OgE1ggvoNx5HeTjoZtOWCxO8AUxVR+yCy7mbECFcMV3YCTJZbVHQuHI30XqI
s43PQK6KNxVceu/R+d+Z0a0iPQw4S0r1BBFCM41a/zHQorDkByt+8g85OcWW
bUzViWG5+zEnjnEA3AuPQaxAgsvvFsFOAYasox1TPqplSyhS7LeP9f8p9kJi
kQq7mzzvYVhGHj23TiFgTkKHQxI4ZnghSPrEgkV6nlQqI3M1mCVKXpGTVy96
tStQNMpwBreE75pyJas26PjL/USHOxG45A0TYVFX1gQgPhPdeZ+rH8QJ9ymg
VjT1acK93zdc0mxTS1Q1y/aADal5obu+VLK1iwhVrjx9m4Qpg7sf0RkGm8TF
mbxI7822Bp/aTS8ZzKRt9MJXRmc2QfDC7DMiE/yhrmdFCwvM1jyBEN+i7RUM
PJ9CwTxrbDdLcdJe/R2zSnDhrneepJZBSt0f+wIgigeQcrA1a8ukOG9Cr04q
aXLcrmr6bi1geZDrxvEYC2Nc5meL52apUbjU2pP49dRTTFy7H90HmrahvZwN
xjvPZoKr7AHS60dJRyKaJJT51hLjvjMy+1cxFHnGco9d5c/PF0JqaPmKc2fa
xDez5b3B+o0xDtfdrauTiMxLecdnZ/RKZ7GORvjU2MfYGnvqGhr1a9Ymb4uX
kakY7lTzGE54bzMpj5cqohE2p9YCS9wIXYf5Y5ZEk49a+I+8FdC/rDkgM1k6
QXLsOQQDp3LtPjgc9nV0S1I2FLT7SYq1UmH6nShX8+OsBZxynHg2g9twYXWh
B5K77XGsKUoz99NAjO3RVBexBdVx5+GkWorltWvLK8MvX9vcmffv9ZptVtxj
A5EkcSsq54lXfrGeVKuWQ3M4jg8OYO96Beam9jCU2v7786X7KO/Az5jhDlhA
as1/nHnJDHdOzAblcmuhiBn+lF/b94/1Kpy6Hle22h9N2M00UJjk7Kp8duCo
grq91D6VJmzh0UQKyvOufMJNSkf1UZdBud6VYpn2S4Qu029jwN21tBhuKh94
saq6/KQUWM+ATc2maor2KpRUK9UPfnq/PGN/wFdyuQXIlyJNZW4dV/yd4i7p
ZDTWRayjLIZccgZAeCHU1r/DLZo1IjOOdDCJGedbBc6SKrZYNBpuoQuWBf9E
FcDYZ42sgzN/KEFMu64Q4LQgb83ffrEFKHB2HG5WKJ8cLbcIWWiCn977Pf9v
FLSSB8Uk2PSQ0bKSVCpnDiGqOiq7FsbSrUk8YDB8hsfAIkP1sH0N6C17cd2b
kn2xpcutazcUbjFfD8uHBBqAQ5VSppRx0ZnX0j22256L2C5WYm0aaJASFYcC
TERFlVc36wb0vRO1WBdZW9OycsxxDVdmbuJr2uAmHTqwusEhBzIpUPu2UnrS
4TIhWuOeXrBMTD1y3gFZNe8enNwwQjHX28MA1n0IWA3J/tlX2xpoKY2lwzpH
4qQMK+87osiNA3kBC/dYpLZ10jHWlFB2OkOwoLvAYWo6xMY2dcEgjsttNABd
zSijSiN52hZ7VmKAROWZ63yrZ+oy+C1VGxd4YxOSSa2zr7XyXqnIP2tNi9ck
umWNgeh4CEYFtNiqq4CUJmY4ERZBiJCC++byh1tGLdPJynwscVe2S7yRvGVM
Utx56ONmmdaelinMIvezpxWas0Elqxu08SNVnJCc9sbnh4mgmOwJH8NvLDNc
KLQ1ySWfkbwJMMs1PnxBf5+K9RRdGp028Vdjr0FurDjhlMHOIkH87UkJBnZc
aeXIoOTDTb4Lp9VIA5Ja4shg4UHdoNrSs8iwVuqyTJnY+vUJRyx52SeqpRLn
J3sSPqzN3QAsT2u9ttQrGvYEJqjezr+ddk7a9da9EzNijldsPddjPrjdhgCA
AwJUJz0RHzR9ZIS56iJM0MKzav6OjVYCSmRwaB46pf696FEoLXf12iFKPssW
NSOGKLbY9wLTUMN11jQm7qrbkp5LOfvohp+HBskRqwCz1fDYWAj/epPweUGb
rqzz7nqh04D/lVkDFomcP0eOvesoF/bwFIDJ002tSqD3YvLNA22IeqtlAi7+
+SL/F1YtILwbqrJ8TJnjdyCSCLS1/nXYgmRhByBupL2M9BIlRW95bo6aPlSL
11f4ItqMqA8uHbx1U/qO3WvJXNB+Gl36rnFzJWRJEXtiRKl1a2UHGdOZxxG7
Hud3I/Q0NgZfsXPGn4WPZABtNKAsyMlYQlurvNvexrrZtaqCNkq/RXAP3B4T
Jd6dIU9uTfYDjFo9yEgsL5/MVTEKfE7fllltQVQkQEDqyWQjUGYzFIcqqpZi
O0CayomGjhwRCkqPKVhL3+LzZcIB94fIhYWWzWfzA4Sc20V9DRQvBBRZ7Lc1
4CwPqMrAZrjt6mb87m5hBcMpSq57pZx1QyFfiqm+cZn09uQigQvw+7SJUHw6
IupzUX6i9TGdj3n+MgRbL0c2JmuQmpriBJYgACogPP1/QSPpCcQrXrz4Vrnj
IwneuQHdxqjgn/q5lTa/pLNJQBp5HyPDgIezk/7cLPLmpNXDFZ7rLA40AG/N
C/3fbqlW1wjXrqJLZmeq9HwiKPl800qQBRExtRbYF2JHhhXXwpHxtrfafUZC
p3C7KlCkh/CMa8MhYpileU4CVV9L8ieQNLKyCTtKgmnhn1cSAUQCquXZxdr4
RydvKOs0tGJSYUNH6PuKxO+d2sDeYKOvBa7LgDvG1lJf5AAZrcw3DxQMDNxi
bAUGfSZvU+BFPElXEXwJsgQ3upoTNQzqCG3D4EBgYp2wkP9oEY2eYMWpiQG4
BBBuGaPQpk7l5IFAJHe4cVt3QOfFrh1bHRS6z9ehl685SMX9EbNOJy1UaIQv
KWVnrko8rhFRH7CYqEZ5e9oSFVPtpL6JkvPY6DzcbuhEO/Droo703fpNcs7j
GhxhW789kknoWFWJoGEb/vLLC4eA4FupmB/7VlXmOKSwK7AN9754OcfPGpgj
zV+uklQVfgum8HeYVYC+9BcoXmtigdHEmmIG0Lv5NVge9RmPIoX7BBRD2EGP
ow/WsvO+wpJ3KIWQxE9dRPhjuuL/4puhHzWaGuKFLiOmnzbju/HdkVcykbmu
c3BzsvKutYWq5m0BZFOnmplDs/VSqVDIwXiLYyc8wyTE/PzPITZ7G8Ignun7
zxJrcyLGlb//b41duISHRco/R7BY3tDnnycLcGYyIxCrFvcKWu3URgO4/FM2
G1gOTBDoHTB0zxL9EXmw7XmEiOfNlqysFUQQtiBV6fsfvm6KBNWxTI0JyWAX
Sk22jub42yMFIWgG4OwShRh5hae6sd3V7xC85SG6yFNa6p69svGljYtVGI0m
47m5NniPJJDegjc+hSM8ry8Lv+9Vc9kTBWtURfRUxvkdKoFCcGXh0F9pVVXT
+dYHg04gkityaMA8mIElkxUT8mZ1YKQHpcZdhkyeZbPvOA5xEXLPE9HR3It0
0ShC+oMajEENpCoz/5edyVMAjnNDy3kfk4XjRNNhtTRzd4Sdk0IiXkLTTRE5
OUya1gQvHPHjlGRU2JTn6hllrLLMgFmJjx6rL3Uw21/dkOGPa8X4o+I4RSx+
fIHvKhfenrUzcomd4TwMiibIUD+m2apPZ2rnGlJ1vGLQvzVLDiKHU7ACoO5l
4v8pQ1qYim3EhwaqbL4cLeLAlu7smAFfL/vNSpdgYZeSfxhZ7JWYY0+xPfVY
BTs9ETFtEUq43Xk1xz1LzM7vwlfStLK2HPABTTYt/TRH000ezVvYJU1y23rK
cElf8aPYdEze15YY0kg7UPKvO6mjcApoBx59JwUmPq6Ji/5jlmriU1R2Q9qL
zks3bCW3yhnkKODd35lI+Y/PqIDLwcjfkdMCoXBp1yeoWBO4BUIkaN5tLlwk
STueOS0OgH2uen2nsuXFJDfXdKhdL/aHg7XtYjYecRCEG8OwjQ+Z9cn/Xd/9
8oXSNISJPSoCTvLizUY7q+spaNo8sNpXfZ3jxZmSmqkPWgWDBGowXCF1eaek
BGUIffFPSX5GDyiFwIDr36K0rhimG4q2B0OlCcpRbjia0sUd2KTtfvYLhkG3
7bhtmoKklX7z3iZl1V68itMjVwxDR9enhFFQ6CVTm2OxALRrbl76+jm8CJDe
P9DyLIekd8gW5SaZ/ZacVzl3SWyiIR11anF3nxwtkXkjcnT93YaGcQrHGuZ/
XZTMju7/mBm0cduE82OUzkkWNaMQj1ps1ZubzRv29i4hmdHxE9/62X6UPnv5
81nORv0IF9QgwNs3vZNf0J+mMqMGcWJytJv5qM3wb8R8Qugom9gz2G/mlVLI
y955+4vyvFqa0hJK7tLsi8aZJwsgjVgJwb1e6i5qGCes4KWMn24XBHAb1Ksz
g/7SNRuqn3LShTcoYVHzmQpvH+IYopAz0GjjRw9wc9EwptpuC7vsT+DoXzKo
bw7i5XCSARjnIwb8/j/rQCSyfBwMQeBGVf0VJUkCNy8QTaExsxF68nZHNP2k
kNx+F4pmdlFLXYZWj2rfGWhA5RAxqvFPued6/79PLtgEOsgF+GqdnVfUMkw9
nnr8+D2dfYQrRvDdgGSQHdluYW3MvNrsZdq/JiqgEfSEbgqvkS7bz6iPQhL+
yP85CE4+njuAQeDmgKE0VE3k3CpmUWqPjFMUDrVCGU+2Bvu2YUwkM2a80z0w
l4EUH7yZpuZAGIzfMWj4Wy+7TNjvvMpykG05JTfMu+OIqLCv2lBWGo6I2uAQ
uw+BFIyHZBdfZ11mRcG21l2Zeshck1Ltls3msmAS9XiIFNradvC3jLDTKAfs
a3UJ77UtPhScNj/55NHwq4bjtpf+bCJ2nUVq1VPOJUhxuxtI/s431lDZm7VA
hJMUzLrolCYrL9iYe0dZIChCxZRf4CSZKnGYkeAQXXkwTr+h5ifyJEEEHn7C
BKl5Y8eaI3UqrWLZHaokaYbMy0/HPQHI+H5DVep1mRNm/snLKPtdAggAur9O
UM/4ejWVR9JA2BZofZ+mGtK6S3xxX6phcLQGXMXyuDcKQyDqEic0Irscejd5
uaGPeFZpij3fxxysrhyB7VeogOPtnm3TmNr01VO6HbH37fWMsRwAhMXrDvQs
zjO2/c6wi7NmVt1c39E8pueWl98hs7Gr7FFq9XWSCM07G8ySy3q4nRZ2L4PQ
pmjDS/Ki1nNRNgud1AyaV7fKwKc3L1d+/MMznLR1aFqHF+1WtFNqVaW3sVE3
UWmHaSErRITrl2GiR89mhVVhh1n1CfVDLJ9KXzrW5K87zb/ufJE+BG8eGr5Z
2rclfLDAHS36WCxE1m1PaHxfetas+LsFdBCnSdgjwjDN828u5/GPB4Hu8lxN
fFjCcPqPPLI+3wlyg5an0u1xiqitKBzGqnpuV/x+B2srkcT1EHZh9Vdx4bgZ
nY6AImX+i13021sSXKtKlJxoks23J7iKYyA0h49S6Y5QHS4CqZsx1L/+g5Q/
NHZewwW4lCHVKmM/5V6V8YiBgUsQJzfajLjMwHhQSkg4bZlr8yoqlcYN/ndK
ODsDG00VvRHr5Y93mrcdFsV74JZxTQh5soazvOnObt5+CmMAl8vfCvszQJnp
HdBVl4boM2IG0mY5NhGLJYB1rYnOyhOnSHq1qNof+itPvbhu1/poj6/2RPKa
j+CQgHI8yKXXNjK+YZYeyfF4hGHfXPBUEZCbzwYXT1uzU1Q8eXslxPfgW353
a6kIqNgYlpUIZqOLkFJmV2XQmIkeim2+o4uj8sg+ZoeodkcJXlFwf+xzEIaX
gCt80uRW+9R1TL+cBQeUKvhuIu/2tnmyDXIMfc9Jc4pCcTHmSKTC77oJtqs9
OJn7JOsWfelzPwr7zk2rC6zV9QF/T/8RcoWwtAv3EhSZ6A5EZwyFvftsVm5/
00IQciaUZpFnimgnfzKIVtSe1sQiwdFpgBH2L1zm3csDzK8Me9uU9FlpF/DM
WFn6FR5J2lb/Lq+2i9dN79KqG4trXEjsxIqxivDUMe0uSzFAXGhoSfdIxzae
oq2E9orRn7oWY5bVOFYXtdfjJRpy+0trjAZmzBRfJ7hrE8upD+rNwi42pt6K
9Gam4nzjC4WEtOFHrVSZZOH1oP94hVFGuIua5rZETRRcQnPVeiH3cHR6Ttyj
PqNMW89F0Dt+8UzsxPCitEIoRfDJXCubSQYCkFqOZxcwe117S2t+pzra7r/N
Fc7InZlWMnolmvEGpZcKlIc8E7OqLF1teKv3LZA6D3ZkfloshaWsxNsMDPiX
WvhrP8iQC0nQ5PkogwE6DOTK+CY+xfTVznLFXCW57/NJeVo15uNE3EO4T+KH
13YcGwycUgXvp6UOsGBGSp4I5lzPZtgyiKuM6LPR5v/b032zbVzQDDXQT023
E9IIiVAauqYYz2o0EF+hsFI1vA77vN/Ry1p5v6+lFehMZOMNApGIJ6foLxO+
Lf1cp5646a1hrgep5iVyMuKh8lu+0fwMKBNcGV4wvtecw8BY+bfq9T+4mVFu
eno1OKt2IhBy/TRKgO13WHQIKOYIm7ppjFh5/RSZLhc3M1LItysAufpM72vc
ZuznZS/EOmC0YJADZ7mZvBviJsvdRPwmHw/vwiz6r15brKHKI5mTBGfTgKYo
lHLKo3rFecSl1xkhYOmJ5ZQpVOXNLcg4yiUqtFyUH4XKY7RFYed1tYoW4r7d
uiojJsf4SFnQ4UUQTK3C9bDGnXFHCgj8k8T4NhTl3tdFLjU6gNV8qzxfSl7M
G3YPN7nXFUyLxMm9b+EY4mekcckU+IWp0+yJ15DZ0/kzGChe6/f8tPmAsXEp
pFuFJOMmP8Mw50+zvV2Lth30OesByp/4KxWYXNIGYtAnBc/ttgZ0lBPhXpq0
YUP1QuQoatYSGQ6cuu20RtuqyurN4PS91qBUXuFS/Dvf2vfn0ITrqLoPzxFA
i9YNj0+B2l5TS4qLw2JQJttL61CKqL6hLAvy2SpoMsgPD7lmipTs8hSl5/eM
FY9e0INhuNr/V9Uowarh5plDHjMPt7bguh8K4YsbokS3fMaxJR94YBeAEIp0
uqeFQCkUfgw6AFDGpq2BBjmLfjxKdjayaOaEp46jSE9I48atbPlfkUNr78A5
4czH7jxUBomIUoI7Xonax+cnjgQWWS/6a10DDWK/6Qgp6+fLbw62mKSmBMx1
e4KrZtXFCHaFzACJ3ZlqER2keRYsDPVn+B3nLLo0o+iTv3R5TYRxPQ/iabXP
TUEAJLyn4A302ntB7/4NBu8rZ4PvlRYOMb++y925umPCS4p9MtGmpuEsctvT
jdzg7bF6OYq4/9Ed0a7vC4O/z4FyN5vem7QcLgz6+olsymvlnSkHBXCielaR
OANchicoXs3WaJiwlbkhJvjrelBJs+8aWWAd4Xhii5p9r8Fv9PSK/R+jUpYh
EjDhOOAMTD4ddiei5MBap3A1P55x8S4RmNkD94lYvYlXC7yULGGrLydw9MiU
XW3kndeEwALygfvuZL2vppER7UA9yHL+BNe1DDoAY2AGjge6vVgUtd2dnYSO
044kF+Wagr7DvJupD9Ne4Jrb8WJb0gdgz2WTyiSJRDKrVtaKEw//daYrkJ/D
5IN5jxedS7DkO1rwMhbc2K6bx8G/HoZXslC0fVO2hRBRxG7MNZLCSmbqTMEX
Vd/mlSUQlTdEyNJfGdS2H1PNFd/dnHDbe6mBeSVZMKz/SrGK3A+Qzv41dURo
almiJqTI4VcmKA+sNdpTQgk4mbPrYnohCLqYffRlnk1mF/At83raGjycXhgh
0LrVC77jp1suhUTsRtNDs8+J/B1WJAgaL07Dozj2JoxrA99YSmqH+jdGASVz
6HCU3HCrrPNWMSQLymgMei6IeJ/6ZZREDvW/BUEPDmF2mbasS8nEtwDzIgRu
jaZN4+ynwlFBQmxry6Uf77tN10q9ZoP10Hzk0pUjxNqeymImdcqPpBrnQ91K
/8g1rvhu2EiCUO1+CyX5quqonVSxGc0YcMqhLGnO80jt4T5ORKdmnyZSKr3C
1ctfk72iTKrPJaLoSh7yK+hpxdb9FLnqLkuVbn+HVUieZtkQ4HGTRTgOncAy
DlDd7sP+a/CwbmtKkKRJsqeSx0cB9iLAY4dWqC4hNPbglI4mLcar62SOWWuq
EUO9RnZXzaLHzKjfTItqe9L7MMNT6nTCtVSuW+FwT8QdZTRlZnGDliad5oDs
cj70EB1p89ATL42q5kU36BxLloED0GH9Lzw7/DuAY4L7jSmdXHQr1ZedyO7n
fUp2pxDDdKWrrFaX7pislEHwQGOaMCzkNescyDs3V/zZqkSWgIqG5uFuexpo
8uawnNB1nX0E6cekppgtObq60VhnBl27JHJEKeZyOlp21EHhf7VMgSOYv6lE
rXqEu4+unDl9GU+YkydbmzjFO1W99auokbUixXnZnDdqdfxPEvKQmMXqlJhT
zqKR3lcxqgg7JkBrZa2EFXF8asA2pIWCbrKokDL4sdiz0zH7CFBBz/edGmm8
RqE++gr4OVe6X2sW5JZFsjGNwWzRHl0ly9IE8V5heXWgEseQND5uVwWWELMc
uyQ/k0kkKKxYiNB9XlxRJ4OcxwmGUqLBFx1WXODQhPMjMgEZTwETKuIGEoRB
46rsrWc/YLeUqkcHgl0RkqKkXg99A7WOExarWZ2c1Ktu22HW9Cv4avSlScSN
w5nA1f1d/sdvInsTy54ldsC4Pj0i2RGZVL+/iR4Xe4YNT4snn5lKtcKferjW
opCyUw6EB9sauqL/iYZhFpAdd2vgnWKXUdHs8u1g+Mwepp80rBxL3hHYB0nK
OaqVGGeN60ncX/sUnp1jZBUV68QnWgBbwlkfnNENTMRxZgXP6A5S1mlMmryd
UGbUgtPaxNvZ6XdjUFFSRCYTvOpHA1rXy/IjneilXJx36HQkkFt8mEB3E93n
659H7jx+IA6mrWjIgoIs2wV/nvoaFZlhAZcLTGUx+rUNyx0+wvEfkSAZCYr+
uNOYbhe2X4ccxom/VXHti3OVKa1d8gkT/25o4eFxbeLQ7cRD5qhx3/o0fBYy
45FaqZtnvcubrbQCTSGydvFwdgL9pN42weAQVSzLWyO7MiX5j17v4UWscAu/
EbCoVrlI1VmC95J/OnBQeBH50/byPz654Qg/IPdQuYtoe002CdCnQ2HwU8He
3SUg1YMpv69zAVmwFAUTPNU0Vi+M8+UCU24d5CzcxLs1n/IMU1jOt5QAuRrJ
zukQ93DjsfgJx6LSd+LaKGmYYOEthWU+N97BMjuisrbq/bNs/mUsBOL3xwPY
F0aKSjxTMla/iEvpNNXo41Dec3XI66xubd1PUrBQHr/xS4paeAamNMGlzvVe
GZ52MnKykEKPQ5eZTq/26apqH7ljHoOL9syeDwHUE05T1n+nDyGWK09uhHnE
hhIJTXLeTka6fzAZcQLFMYVWByDWvDEuFnEMfar/U5pJEXpoRUj5kFd6rNUY
AdoXAgOsAaQdQZxAZO9WP72fvHYBdkPcAvbtAHIGpL5An/zUUc9A6k5ibvJa
ZJTLGCpn6oyPDr0T6b4hlVdDnxiwXpQs3rw/bb1UTI4nWi/TqrMaRYA0TvOb
qCIFUDQOshViKhO8nHD/oXKEA09wNtpr5mshzQwTALBne9TnjPZFEBEj/ZWc
UOwpRj7Zj71/ltGPwpcS19U8Tl0Lx7K5T0ABmjoTfeOEVHz4SoZezhSyo4oW
wPEsgwOBmLUcobdTR1T5xL/E2CJHvtQo2uq32n1skg7WYFzPx3v8LEyBkIAJ
FMrx+KT9/czjkC9EkR4bvwlPM5jtgMHKgXF3TkYUFgSQHUqNDb4q20L7iAfk
VLRhHXErxhVcJ8+Q0YGd/pdNmc15uTKeWdUOzIPA3PdlNaC+CU3Tldgtt6lS
HIdUHVXzy/CEzQwevWPlW+6FI17DNC4poNHCDQ6uxqrhwZBgX/HzBeJmeFBs
8I9zZ84djxtozriktX94lIJE+JKV0902Yn7+XFxZNo4yiYuX1rTvFAfljc8c
1nfDaR/Go9zg7J0ZiyeqRKIYbFEvWdOLVnC94YJDzsk/rSzma/fsOs4wCvaB
T66db+TbXLxAvzvjGMlCflPIH8gJc4p5650BpH+M2ZmI72vTFh+CbCGpy1U1
YGrgb3MhL8ESTu32PjS1kPdvH7lbVC6nSOFKjmPw5Vwv9VIvc/62e4FZXmCK
xXtLv8jl1V2Ji5OWEhC5rlEs62R/xU7xPIyw85Kn5NBCAG8LGHXV904/K28E
QD9BY2p06JfwN7Z2mEXFMt0Cgvc0+En36XDZCjmEwHjQPpayXKTBYmf4ZIf/
JC6EJbUP4uMQCBFffcO+ndmhtsjkivc3eYAS1Z2d7KSzKgQQK0jWBtKunKZ0
6ZEJIyE1mhrLiQSl2Ol1AQfcKfo8ZZZxO8ps6YNCRTumOuNNyaazC6ETc3Qe
js4ABZTwyYh1h+Qnv7FjwWBuZtnD5U22ICh+xdz5XFxgmn902lN4pGlPJCVr
TPMUBpyV0QK15VKP3cskf0h0ItAGOFl1UhXVSCuyxy0f9GHiemfDt9J8hbT/
QN8iyba0n2P/UDSYyMUtc2V3kjvRMvdcmMRzXp9BhKVBheffarsVKqC8Nnzb
t2uLxbstmgdtBbasrlMMw/iwWwmu7Gewqv0CpqYzEPJ4Ot0Nf+CJFzLk1Xu3
8t+UTV5MN7HmI2W/lYhABvpN2TcS3K8lPlUIYjAjPOu51xTm6VhDx2fr1T+4
tjKYa9m7iP9nQUiD3/Rcfrc8qdnbaiKDQ0yfd9vj5xTgFRR3cMYv/mKBUkzK
rSD9J+mRvkFEdR474ErLvjFzuqt4oNaAH0qv/UkgWAzD0DjUfPqm5SqUcf8J
kIu0u/9Qd/dpo9RD0NYsF17lEr4+4EMMx8lYrZbWfpjBmSTF6czrhVJeexuG
UNRXjuc/pFlo0sNDNRVrqEiFPVpwhezXMr67Yxawra5GoVlVfVvApcnQ5lW/
nJhIWBcocGFQ6FHJ2by9jIsq2vUGa9sD4+R0i2Mw+ADOCK1RiRTqNY84A9HL
qETUXRc70sEd4l1E2fVJdpuj1ppnlstAxZn1LYd/L00xaMreFNlO4vElkTWw
0UmKsAbAvzydjt4Of2ajPxpbL+B4SsfkBgK09wbOE0wXL4jvTkpqRiUlvz1J
5D/bzXu3xO+ZcUjqWdW9O9J69Jk/x1+L1Lvl3EO7NVkh9q+yFtYe1cRdzu7j
ekZ6lHc0zjKB0s+TeCoVhYEp2j2trvjiWqotKd0cbXLM+IkcQ+eO3Q5U/qio
EdMLJ8Og+plemTOAdVQmEDM99ShFojDShPT+1bPUlcOB1zjRRINVL0/kSdj5
Lv2icVNeoViIHy/J7SLEywKr9JKNBofoGQx4cPA3IFU6jFJhVoqkHYocTOII
do8ApTjQ+8abJSJ04fKB/eJNKgyjq1R3Q70h29aqEtSzsQOtZ/uBpR5m7QLx
Pnbah0oOofs/Xjo0DB4VGUDxjgpYcyjxgd5woEuNrx6YvjIUYeGkmj9OSG+i
bFQD/c1Ea8SCDHbppwvHm++sC8d91iKGK5UA49xIrq7RaGzbbm20rPXc74Wf
6AUEk4TaWsOU2cmKy2Izma1CbiVrKyVurh+DQUgPsgATCifrlb0xFseCEXfY
/R+wXxe1xi0eLlQxbrZ0kSfwZlt5TBlR2d5RwZcKiB4tCG3F3Dgkzqxjn7B6
BMECqhis6mKAB9e4F5iPwoDtP+d1q6NYvGIZe0/bLXEFhZx5fZiBphnmOAGg
+lD+V+n1oefT9kdTD0qW4/EF88OLUZpIW0yOSVVUQgK6gyaTlnHkfUlaTRae
SnfTeqP/HUf2zkZGFgP4mGqF/dExn6R2ILYfXFG5G0GJ70m9xy1vUpmNdDxi
D3eDfJVzRyvvVl8S2rrCT0LhDuvQfmwHRneQ80+jahF6TYLOB7kU2i5tkCK4
ghpMzZqOH6B6gw5eNf+ziUYeFys0+Lsnrz5s6tvVnezHQ+lVnuqK0mYI3w13
tbMzGyv2pIuwhe0bjj3AwhZKxhC9HuiXB0P9yxJcNEUrwPyB2o0phQnq2+/6
vpp6LWDgAJAY4Gb6nyW/iZBc1UwQObn0wlWLGH775mAv1BlkDYmdojcWBcbb
0QEmo5Iw5psNDDnASC2VTZNR6vMR25EGrr7g8Q42SoYMpFSVmIW+x2UdHpv9
QBrGAW0gxGBJWjj01To1dF/jjcKNdc9cBBQWxBhN4DACeo+QRvqcNcjkMvyq
Lc5vRNQ8OeV3d3rOYRODHZhokVrVb5G0Vr/SYeEq2FhELduD/aSr7GZXll06
OtO+V5zApzkgYt29gDmtvC1V8LueneCRrKqbuJf9fHa94Ap2JRbhjgjvcG+z
oU0Yf+izCTHzwhF+l6+KyGaFrbJOsU+AIV2w7nfDrbZDdXOk73+jzvQEkkAj
Yx4NMPxNsNDOtvc7VGgoHphEJrxMC3awHQACraHIByYKcHeSJhgpOXBBsPih
8qsJxv1mEZDQywn0ffWzWivnw5Pn66PyHAb5X1fFgQien4ZSwSV2bBbXAOEq
QxkHapLdmcWi1V05FqOuD48jqZK2bsF9pIiV3+lHRimZQEvRDbQfnenNcDV+
1eqaLRKfhI4E6b0vwfpq9qEsUcLN241GF0Ka5IpMx2ewLPAcyNAr4ccSFJ8q
S7fif+M5/6bUkOxyH1jsk72nn+jrKDOFPtLXGswFIh/NZm6GMQC468Qt42xv
08UYX6FVeP9zKTOHGoSic0qnd3KHhob84cX3ndGKMa2Igj3LUsZMQGwVJEd/
CYsR+gCZ/husE8bqBi6ba6eoNn2Uo6Qm7VKrVyXGHcnle/iwaWXODl4PaIHc
Tx2icSCOltBIpgNPFq3rbi8FukHtw9WQK6U8kYiv/birVzDbylpyJkroccP9
Ni3CB629Pdz6MZEXTMy8ROqbRkNRHxwAxGOEG8kr9t9vYHqREhY4HtIhQQhN
SEQxHcjDpck9rL0fgTVVFdoEw9HiRuNq4l8VqKWrXW46+B1+XWfyKEmxzTln
BBLJhAiKD+Hu7heYHrPeGN5ZWKFr1KK9CECfmXpmmMS2qG27uRU+PpMOJQQu
umKFWiGuvxDD8A2xUts6A7nbanmroDjZba76hU7bU2P63W+oNCyRmn288Skx
zqJcI/8qKqGBjeHjUmAd2HWSf/sVpPS3J6ARvOHpkPm46/NT15mUlFOZihW5
VjATTv5p2uffqWslq5pmXLbVp8QfBGQsZ1LEbsMCy7Xu2FG3Cld6hLUSOS1O
qmRtVWi6iUP54R8d9meUTaN9Cd9rg6Pdf2XiImZJo3ngF4Ae1AR33Z2yAMLp
LlGYj2yWaL91cEnFWS9oLz0crLqQiDQV9o6NzCUArTV7GOIAIQwvA/zbSaGu
vsemavpvvsdNPC+AJp3JiT3E9GhUq31u+sExHgc7cdoy2EKgQJCFM4B72RHL
fNBWIenOSdao+tQ9RMTtWkoBrhHAkXC0zYKz9RNRTudHgGRbtss7qd4H/Ed/
hI5bJsVJ0h8RjLatJTfqDqoTPQ5tbZdowgIOvSF8eAhoG2ojZnN/t+g0rqD+
rEtw0D98yC2GUhE/c9F/kENqnPwAjKYNNb69WhrlCTWoerJrIhqNdgaqh/BO
1kTNC2cTvQSa96qipt7kxmTgS8H04mjkuXnHDfIYij/qU5XtTXddqb1V2YYN
57TnfgutI/DMaCwrnrtcnVnlfGLAkWcuO5GIFb1f6JRNwEfi2r361JFzV/kV
EKW7gS5um8xb1uF66Fb/n4Elzc35MHZw9wTvRKAAP+G9cnjXCEhKDzmBMj4F
E8CZu7CORyOZnDRH8qs+OosAEeJlpwTwMtTPTkJGf+VDITrqCd10+q2Sb8bT
zHA1kq6y/CAMlkOT56ppteaLFlm/ircJ6+et5MdfiYojTHXRlnIjFCvO/m3A
JHPJ3/nTGclR4tndd8fgQR2QI2f4QY6YOiBAQBxSwTsiJ9XMRPIOuyvWRIn+
YV7l7Zgonhn5b5F6HyNhQOw0/S7RjFlR5AmUpNwGceNBw6q1cQo3lIJ5l/Xj
gnogvbgs8Hxx5t4VccFg4UkGS48Cu5e4sFJ8KhLaf4iySy/olGoOZhRaZCZs
rR0GERSbkw8CY69O8f3nnCgME5v5v/ubGrPJZlbdcxeK0gekyHt0qsNHERLJ
ZuvKvGpEcbBo3G6WHskysNYDc578foL3KSOAUU/K+QBiUAEXWtVWUp13p53s
sukAIasAn53AQfQj2iq9ZYqm+wM/XlV416cvR2VZedCef9pVJca+JuQv6nTY
vjWF5zMDs/WPx+qZP1+qWhe1fJUn6LnkkTnDCrJk1A4ODGcYnRAKUHU+dvL9
s7rrwuON2ZB37+TccdKFbhavTLMBQHTpVFX8VbJHXYX3nymzWTdhZ5ZXLzCH
KZqzbbQslozdgwUfBAAbidLbCMTwFHlXONEc494IyrmeS6apNYOxRrQevKHE
xfovqGacnCDGBGRQ5JxBviMhuBm/JqlcUw86NkjmpQmzekcJdpe0tYU6Ixif
+PD9bVLUXwVjmt4cPUDYJy1SCoN/PFHWfwXelYisiDu3tN4My1yeDmlFZJfT
tQKnl3zbB1T42zrZtxUtlOjqWTCh2lGLHslfQdzIlmagyRT0HklYUmRAvPGT
2KQjrwlaemIbueLvRajzTtwT7INHqjwSjG/vY2/TxTZoBm0DhLb3eGOhdcyJ
YPaQVRmPTq6zCdLbb6AdpAJyK2Q64XkaSqQoxg5PjY1F5XwynK6GR+bwmbeZ
x89UJzvaeDyy0CGg/MKN2lU6mJ7wDRyh0XWcKRHei9yXMDRJqqTbQkRFR+E7
NekZ/tiYjCJ98Ii3hz6lPTJLSs+9tj8uWbeWCh3chkZMOgvuH8Wv29jurcEi
SKG/qg/pvtBD20qg0qDZFfJic6srRl/bhPFhTO3WeeuhVZVAc0Xj6YpgKLTd
HsFvYD69tSNiKWrCon6F7CdyeM8wvwp/hg6IooX58Up8uwsggH8yQ0zLaOsx
LCwoaAoPxBNLmOBUGa01wHfLZeeqMHkKJzz0ZgF7d7rzUG7NMGzEENm9leKe
aVe1Eg2ll9aVwIBdHp0frYgh3CDma4fYAoLTmU+FO8Ge/plC+YHMpU0Z2wt/
UMDi5SpzSR7fr7Z33vJH9Vl1U4J8NPA+hEHao62TftgMqEC/Pg8NwlfxM4qJ
6qi7KW/FOLvo+40k/xdDLdRCItghEI7KU869bv3LtyW8chdqkm1ew8wJP4Bg
ARwewF3uEuBNmAtrm49NVRSk5C8jUgFGZTif4GXbe+yDZ0nle94cWbTjtNCk
Z/Va2j7uLwwQ1nWIWv5VB33Wp7hPPwIK/B2qTuT7n2PG/0O0DEdj3Ghfz60r
cYSGLBALDcyRPnkKA0cL1B+Xptimm+tD6B6FDcY28qiKD+HLtENsnqqn8ghd
2PG/AK5QVD5ix+OZ999DUCEUJo673EW9c5KKWx81QwvJHhF11kLFTHkFrC7n
p/NeORnLQonbVVamFCMNT1ztVnc5gdyQxyCYv/PdL6FCrLHmsgjStP9A02IK
9DzlptDbdqJBFClZEt9ryOBLNQvlTsTmZrtrqM+3+YiCU5Zt9XR23IJxcMCL
LJS66vBY+ikW1518EoATw29Fmwtx3zdsvGKe9QP9TrNvoejcG1arjFozfPdD
THYLBemnt0OqHU1LYqy980MeBybPdJSLTYtAh0LvR1ibIqUEDB6IAZUWpfwe
nB+6uzUzIucFmu0SjuiVJNUm/Uz5Hd/iEzIffDUr0QE6bYrhorToH9XFa2Tx
Cg62s1OaW38KcjObohfkkLhI8s+vdRThSz0zZI/x3Q58jCIyA5tb882NIoI8
9BShUKNvPW6qVkkWtbA7RKVOY1jGPW8ZZuwsGujjFWTQ4/EtUpRYLKJ/e8WY
qqYRfTOBNMj2HB4A7rFYTMuh9z3mE6tsnmzToiRGnKY5wgv1XlvKPZcJS6bR
SZoKiqLbslPkVHvkDyANO2weZP42njrg/Vi8RTGeQ8xlnkLblXSFa5SacRlc
PxplcRYZak5hdlf1kD9SXuGiabv9L2DUusM8gp/rLGhJk79WeKTM/X9KsrmB
ZRV92Ze68t1TOPjPz0IIuc4vu/nFbh9e6V0oPNuLQ2s3XVvYL1+xuPD64kwv
M/DotR1/2CsZFJcir/pTF7sv3gmrfREMqx0YOjZbJa4fUQs1lbCtPt+7XY4u
n6XNDMjjwS35MGlOZRvstxL+/jc9+pFhKzVSolHR4f+8z/YP0algM/WG4KDq
G2Rlas6pMRUVeXLeJy/Gl3/ycps0ryPw/kDtSwJC9nwVimLi9/Ag4umSvgNO
wLe5C6X8mQ+Xr22AtMZ8sBKbkxkOsL09r++RnH2UxZi0gf6b/0C8KaIeZUBi
Nv11nwCLYv3D79VAX9zCSUsmWSHKciBcpVz51qmFjL9xYJ8mX/PxhjoREiKv
IXgmjoCKMw5rVF/7xORVo4LB5kA3oXgrm5Rgmg+CUrd6i1YYIlwoEbpdGwu+
m7rFBlAA1raKzpNEaT5YaUwfB4cIIvTlQg8TzUYZRXY9rHbvrSspElgO4BOe
dQv/BwaXX2xOAB1MP8T6EpoThG/c/TZE518hg/9uBtxrTc3oeEEmjlHaHKCN
0smtFuFTfk9bu8olQkY6on9q2PF/xSyiuYNE8z8Zjqee6FD5RsU3Q3q4C0Y6
TDngsKsWjQldefqAurjOhY1IigLFIyhy6/YBO+OKv+wLwfK2Kfae5lrnclfH
rMs+EC7ucuJmtLtbwUlst6+N/iV7xVpO6qqQh6tE1THS4C/iAli54y9MYb1J
/ZyxYoc/WXXnUUtl4Uw9Bz3Eptjy+sjnDQOEODKkdDN/OOxNUhQ1Lb1iI+p2
XpGG1lSdPuOIa2wRC6TT2zn3Qax4n8hD4wSDSw1HJCL+1F9muFy4tAFeTTDL
9Mw417WUKRrecI1sIXHZTtL38jiWQB5D/p3enL44SjqUTHqUqt8yFCN+u4cY
KBwF4kQke/sSbMPnsjZFsJ8Cuz7Po3WQRo0JW6o9kyp0WI7LuzSr2wlSWDXa
kvYKs/dHrgPReAN/xPwCSe2tCSDjFmyhfR2ESVGQkmPTd4QMMsE1JJL55Le9
bLNU2zS4trdfmyn7cwAyGbzaxMZReEwJ4OSXBQoNUU0k4vFcT9FgJhhTTzy0
5nnASXN+rmGj4zic0qBCb6tjagS+OJeuHuxZ0JQHart4RHmADzASiMTaGzyj
EwleKynfqqf5klHFTOTuip5bfT5FXKIuUNWEq1JURTKCROrxDtGTVfg0RE6w
3ca6ZuvYx9DTkijtdWa55Tficpvnd34PXt/hdg9SVIxcDxY44Hdm2ZMfl4p2
7vHcRP8dliDfLxXPkJ5Op5u5qRtDzZ9tiplFeP13xASLgtkqgNZ36SJXNrHc
sB27pE3O/lce4ZhNJxusnbsX1m+hZNSR81DiWeL9oRwSLtFhAtQuuhQ73sUh
ERRZ7iTX2oHXz7s9q9BlNBwwlxQEFyrIqLq1TjDM2sj0a+0uxOweFnG60f/X
F8Zblvaz7VRDf88IIUYeFsrmcWlxVdhvU9I3IPGX9jk6lfMUjn8BCEMIQ0LX
72dyQ3bFM70LplkomMxeegHe01LEGYimTCn0uyJHz+NJ4CiLlaaRac/gi2vG
11V0NkfNaDg0MRrwVQMxfPu/SM+PrUXH4w78CoM0DKtP40yUD74t1x3fM8f+
YsiNxXn2v0iNSw8x94wu1nKs3PgzjJngm8dyXve4cGT4DrbFygw0hc8wU3sT
zYs0/Hd+i9YqF4yoqj/zm7/dCllgYDO7ypx1C07W65I42aFBTZIwCXshnQLX
VHLxx/nKWP45cyV8DdK1+zeZpFQ3j80YyGCTDIfzuqbNU2rP8BXbhMW/2G5U
eDPdc+Rm6cy9mkML6IEzDLBaSLLSNp4Ds66HpZG0e2jUk+LC3nDog5ZmXkzn
kfq58qADhKs3gbD8btse/rbnr/0mMKyHeO865ggcBfXuw0QNeag4hRXocPz4
dyM69Rgg5QpAJ1dw1wuAF+9ESd7e6u8/9mPaxROAU5dM+1VHv4Zxv0pu9fal
daFCj5SOApB10La5Q4ZjK3H5+bcPAHnUUdMX5c6Jd2we2dvjLMAbK437y0Ra
cBvB9maPqdfa+3awinDJpdqDokRcdrhN59o8/uUnqg9pWxRUs41Q/cyIvzql
Yjb3AP62jFawNyRMqdBOGQsY8sEoUYQ64x5/kxtZ/V9hVDP3h1Wm46qI1zeW
AKzuxYLHQ+SV01yVrIilwCNUjI3/JH+9AWL9qLduNiJGlMb32Gxz0qZ47sAI
Ec1s4q2z3+jNHntxD0lqiXYDB2O5x5KOsAgcz54xTGT6N870jyIGZ7wQ3MRQ
r1wifMpA+9L51CiOQA8nXCdjU/P1hdYSN1d1KfjL9Ro2/cNcfsNOyo9vgO19
7aTFZXkiZEVZu26uS+wlVdBUZXgoRFmY09CWbJHYNGowoRLuuTtL6nMMr4Dn
sTjjbO66OOxBeCM/BeayBNhmgxpGuTMLC2skDZlmlCx7FPtWSdT1UFUYD8xi
t0EbN1AvXegZIDyCNog5Fu6MO1L91wHTI0N7hGw6ZGUkk2LEE3G+1ucYxfTj
nutYaH0XgSp+EkLNHhG8Rd4GTZ0Rg3ZFxWGpUdp4Z9kHL55LTIE5xeAkzNV2
c+jyNFoDKOSPvztxXmbPI+lbTJdoJDYBW7VcboYw7ukAWb7k79eqz9vCVlb0
i3sGah/LeuvhIJ/Ppiqt5IGCGmxRVnv/BaZMvuSEh7TdcD8KtgDbG/sqmvQ5
EAv/LQQLzmBYi16xMCas6jDuSoKU/koImwp5qF3v6ZyFpHpAoUwb1FYeJGeS
9hnfd3J42GA49CH8DVv1mpJRo+ZoTnlLPY7INXOhmX7VNNHh+PcvVxeagfAl
3rs86Mw5Yc87XVN+wjndJxnvn0jOxo8+X3CUiSBueI2GWxoTRXDIu+Gn8G7j
z9AAMXIlr8C0zuD7pSEoEnrMQL+JuQ6DyktCDJx8TH2wjj/O25LrUAaW3i/R
6wUe58yPT6A1qUtnhRkrDWoO40WXYCu1opQ028wh66TRXJuYUzGnTQFMKXI5
lKKi9oemWOSRgJcmWnCFWRdjOa9hZQnLHpzuCpaQCWO923PGhq7v9utA5Y8a
jrrebl6EJeinzQHKhLtmWAK2dBEcPymIHYDNf/3hNNRPuHp485d5cimsHMql
2Dt8DDqNNOiDZgULz6aw593SjBaemRPpXWD/qRfEi4EFgKgikj5gZcEtTHhI
YCDi0/UG6MgcMhoZuCQ5RnoTdNcqYzOu/dEbibcIlW0fs9kXrRRVfXtB2Mpt
A5AMkg1d6ilaZ28I8/gq6/c4aiPLXJ6d1wQ5r9FIRcJkG1DOzBCnheHzALzN
K+dIkrWYCfNFUKbM4zJ1XbbESl08gWQ+npVGJD9oWjNDPLojoe/jRFtSkrW7
ihdt5o+Q/9Ak9xLYiA5v4OTwcv8pMAYBByUOK5XjgCALHhhATJPgf4yK5gz+
lR3NK8Z+u5ueuKYNS4blgAc1IJ+CgIyLe7ptxk6Hw9qcvgDP9ZX9v1AqBHzz
r3Cgbdotd95fQaAk3CqGx8zEmsr5McMKlBA1ndfAaFoei1xmJ6d85JjbIidA
bNQPoPw0Ax389MdqUs9Dhma/86Tw3WJi9nZdgP8EpWQRvkWadhyp+zsLIhGs
StkJYQGfazGsHpwojfo454CbLuwBcJQkQ4ejW98EufjnNfyE//yyMpbcdPjF
3IW/gYlFuxENNZjle3OzZQuRA7Z/cZtkkPLGdRp3i6dAyST3p3QmdTuuc3cG
ZT5XmZ6NyP3xzQHatYpaknesCqzKr+UKlKtNRTYh2w/EJp/jxzusUSeyJW2N
V26q+SrlRpW5yuMRGMre3fYBnFaMpBVC4C/I6y4MEw0WWeO4SCL+c31DTqd3
Ygn9P2tj6UgoKOmOcoZToZsdqSbxxcSUefozNgtOG4UX0R3Cq1PhpB2yK475
OEdpVn5xvRRLfiEDfj+/jZZx0d7aD61d6foxicIX3yxwc7zte/pS1aJBrceb
fj2mlznFLoFr/HnqMqyG6UQmb4lA5ESZdUqn396HCL5yDTU+aVuukYzgmTps
ixJoKMWRhLp8XFaRba+6FYOar2jBzqCqZVqMNsmm/LyfFUZzL8n3ViVcZB8c
XZvZzN4j228kLhJ8XdOKmb8ZAbIQir7yLiAK79vsZuu5GOtuQSbplHWINf7y
ci3dJ+/1Mnn5GpyA1X69bqlQuyz3lVc2r0tE/B0xVx1IMhJNnGhD/rd8TzzG
4F6AHL5cGUYInXxJQV2NZMWZr/osUKvRJd1JayB1F9wD+eUWzScP3WwGXQDW
JFIs1PGG9sGitPejTBosQAgaw2XaVL/Kxx42mYmv8FwqDlLoebuKKnUxsCaj
g2i1X97YUrE5pNDWqXvKEaFJOWdXnx42/XafyJAgGsXuPOWIFu7ZtGZTJm4G
lTwO/PjX/xzMLUGNkf5sscWZbueaPXNHnerftWeA9zY+AmJX2XerH75dSJMi
PGIQ/4uhd5J8TBrm07+yV9dFztG1u0HDC/xWIYid/wk3QMmgGKP54JG4vSbO
GISXeHjrgBC6XhlZ4TDI5K19JP///XpuOyCurjKIN9kE08uvC6GxSel6SMIb
Zm7lZL5aeKXBI66y0oOz7JFb2QKSpCJ8sXOFByFGjkjFwugeulw9milHORce
InsysUjsrf7oBYhhB8/k7IDZuMocsgdVBHhI50HQu5upXUx/CIA1jtO+e7PC
dIKivuHM5Nav2JF7rWumBtQH6vlG6Ktzz7dG9I0hPc3RQIVGOXL8aluRqc+8
uQT2WjGm9ulz7RcTg/3TDAMVjfcIqX+DSALo6giqMZGRqTFjJdI6cPrCqVF0
uHL29cwaE6eR6EgrFvPFsxvWW7AmRy64p8L6jqQfGTp9d9Bei3+fCn5w7JD6
EDA6l6UHsLauYO8PSv4gIMqEMrSkA63J23SSx/APfgxQXkY/JsotC3XQTT6q
ZIW/7yCT7qgSgs54Mh/oQy4SEMW5sz3nZG/VbDZ21Wzp8XADOE7yWopiBhtL
s/ObqghrTQ7yO+LW2wwIB9eyAyoaDC/OYB+nxKMRHxjB+ueWW4KQnZU5ZEZU
dzF4VGOS9A/uRruUoyhvI+y4m9dEghofXamoWjBWSTCV0/vHiAQmY6ifeJuH
7iz6sRL25qWwNMciLXCK+36wZLogtcvrbN+vzfxnyVR8jIulBKxrR8fN8aFo
9yRXpzR14+k+T+8BVZllHFQU27SJInT/NOvCAQh43OSdlfD521cBL/hsUuoP
DWWWC4B77Y/JUAJOy/+4659fHbAuuHBer5AF57XBY/xpExD9CB1h852HzZfy
NdfK33QW/sazsadViu9oJrM9wlNP7XMZxtlybFJsbE6fZqVzChDdgJzhyYtD
APyRr/AjUpE2m/7VYTuJp1PyMLq4Mxjnr0zxxJf4MVRtxl4/06fLeG1uHU6V
tvfY56XWoEp6fb0OJv1JVCoPLu77ZwvFwCzfqxEpN0ldXDsZfcT8dnoKg3zs
4t+iN5FnfbGS1MjhjO8U1iWSPmXGb8HS068Kq5Fmwyg9cVTuKh9cNfSUjTgV
P4ZlFq3Zjw8QejxaHZqRl9hodiODuGiPJ8H6n2hD/NvRNJ+dX98ic/urlk6v
NVKlZxYUeHhShPCC67QFRWJ/CBoeq2yYoG1AB7Fyx64TNmxJgHxbwgepFOlt
Irep2VGBxJm2kX3z1fG2+9KzrFrV1MTvNKKxZyI3O6HqJbeDOaXQuVcpfgmh
gBdr/t2kTgE4xCPbj8OkPl9msrLrlw/M3Gv1PXwmol5FqzDtGPaACXObbsFw
H3aLBoITGy+l7MkHMZk3WESAaY4mPVPs6My+zRypCaskcdQVeSHDdEaUlna3
gYrZPOiKuXgBfo8JTb1Q2NA3BFfwxwtS2VGmjDxlHCvadsvc0iBRTS+R8avj
dPybG2iabHGb5WUgN2q6hRokHNAzNk3wYIFlI5cCgxLlGWTVySoDO3+MXMlI
Xjwzt4KUusBvpNVq0OLgFqC07g20+IG87m1J1ThelhywIo7WgnOi5apSvFG7
Ae/8Ci6yZi6er9VVTD/A8Lhu0sp6MUnR1CUj7EvxTh/dMv3sRNEgWt+mePBJ
pVKvCT3COXJiW9ujSVLUkOXkp0bLKwnbVkyqBojK7A7yuMKRZsjxABc1P5+E
iR0JrprosWNHiAVTxO/+kOyr7ZbdOKo7iLELlVI1N74WQVKjKdD5wIYC12lj
GawRiMec4Mhwvakj2bLDkckWPLAM7TvsMZPMQXKK6PNjwFyI5WkHPg68w+gj
+Djaf72I22a3vZKG8YpdE8jTJz19Z/gU/xnEqwGhYAW6hkyozLCHfeuPYi6z
6knxIWcsfTdbGBvKRINwJ+xBYRO2q58NMp317hE8RUgvC3gKJ46YLB/3lfpL
cdFLa8TudOPEgFk0fV6mHmStpm8hFZP0D/kV9AkTCnj7B4JQBiYUUj/8ij9B
L2DFMwvPbscTKxwMCkhWt6fLDT5mISy9g7q9aOBNx/YQZAKJTEs3YzLDGQTj
Z+dKXUAly1b/9jwqEwu8vVVaudKhe+luqNXH5RaoP4AnWdx/9kiy+spoPUJA
z/OWVp7aaozJVt+ZZSpZSWFkINC/8KMie0/a2LMujFrmrbyRHJbg2Hw3gI0p
41dzJ4Ud9Uveh9NF0eB4KDyb/1tkGGuHOSzj7aW55RfdEG4XMD6+GzDYtIE9
UyHpqpVALz7jtYJrqLaGINzZoPmbL0aHH9VBvmoqT3DvuhuSiCpORe2iOF6x
LZJTn5H6X2iSDjzxLUdv0bD/LxzLYJ4Bh01DJzFHkrXHATaSf4XDWyevPMSX
YDnUGtnoxBPtG/lHUVToNOPYNqjBO1Z5DauHqJZ9X/kkyGpTTk63nCzmvnGw
Q3TwfIUuvKqqW3umTzFxtU91Tv45vZY0T/MjtJTJRkj19GCH5uhesssslrJS
wY2ZZAlkmr2rSB0G1uVSxuq4oWqyYJAn2YRLWus8qPmSdksnvpw9xDTjmfdV
qmmp8ZsoB6wYaPKKiZXuBZo/CYbyxlf8+2KNiWYaVkauFUA4m2WR9rELxoyy
mvED6deCBLlTh7/WOnATF9w2f0LQXVAKdgwZzggcrfPh/VXVbk4otuvkOn2Z
z0Luen3Pt+86ohOPe0jeNo08i+hon5C+OhLwqodwJ9gxFfYUBdqb2V7Vko+R
PUnjd+JuWCe/5srOLjW/FCmgYJSl4YBzuZ3TfybYHHBOYA689cd7Ee4pASXO
NUL1k8kOA3C35/Ge94gx1Gm3b1Dja0YclOK3iPlhXsZs83PsaFqIOCzz4dBz
tCPG4JoOgrhtp3KQR0F3gHjFl0zG+fL5IeCju4GM6+rzt1Px1lzp1sUxC1AV
f+1vLKoQlKAOhrUk7CBYd14qIJ4JJBTynpkfBgGoUXDKbm6yVMFHk+ap0Aes
+AtkD6vPlgKJa77D0wfvdmBgQ+TRRXBu2P3+Rqw6S8XlPlxA6Ug+gMHjRAzo
RejRU/1indFZh1g1EcUjw1yfVjZfQ+vCtB8IrEF6agSZC0+LaGyxDdl9jsZQ
HsUqvKpQFqsuimJb9de1oufpWCzUPXBa+R0VY90fb2pIW/G6s47dJBmXDFsj
htQhOnnQnqzm+bebDIYXUnV/ZtRRxPZhbnqwYY8CL8PWoTAqH31Xmgnyo9XU
DSOvrSTG78+0JX3/YRa9ADdxVoDyx4LFsM9rvuIBuYk6HT1uZgARUjaDV1uD
IDo0RpCCMRltE4O+t9nw8EYx1+SyWJpJcCXv/qSjN/PXNBfTlTLrKKCicQc3
CZr6aN5DP6GTvDd09L9GsLaYv7np7f2VOKlIkys7myWBHvo/+z8zrs7+4Bkc
EnAslqtIolJ7wmDadNsVbOj7etszVGQ3xDBtzd/0jTq6+GZ1eJFcrRgVJt1A
/ZAIrIf7RqAKBiE63jVxmKs+KQWEYFUHn6GvMZg5lRlUpShmT9HCOTWSVayX
aAYR+Bfr5wXe/j82eq5Ve5HP+xtx32gsuEUVbiwNdFnq+Jn6xLnMPlKcldBJ
ijtlEv0SyBkKxRvRVEMv4LUHb/vINYn9OtIxI9KkAzQsZFrRPGA+EMRRLpDW
85p3/nlkoxJAyQz/lcSMTUy/wN4zzzyHurF3ll70mo8SzyfjbEuEISMTjCLq
6iksI+nLnyd4o33YQiUukunxzOYjFNhKuDSfmgLVoe/q36pMpUNw647dalVt
Cdvzf7eU/n06P7MV49y+Yfzqoms1DxW/5yagKX1UkFv6iTRi7Q/k+zHkZ3zP
Gio0zwBZoHdbZv25HnMhvO5+oGjZo6KHMnwp+Je07YxVULN21TbJuzEyGaVh
EWy+0/OBAEUGsprwBO0rA1kUSbSlapSLDqML+ANa4hsW45hosjYWsoeXKIEz
C2xqJHPdefrSg2u4FTFENk7rSCwkufpV3WZjo4q+/kUtY/6x7oM5XQ9qnwrK
BZ/1NSIAIjcoXUpi8Es9fKL78kjvkuhM8PW2XoPg9GCXe6MFDA8HRgSCjlGt
d6R+kOO9cvJDnbZ7PMFhpC8GxZQoJjBljbez5u5FL7Gw9ipdz+aPfbZbFoYm
qelb/bBtygG2CUJxrJ6r38OXaitjbyo+jqZWk2zMObs8kRqDMulCxM85fP2q
bskCjvCZUiVIBRkdlPFIXQdOCUcTUbPO4XbPiOoEq3O8Gb8BlWxidxH0kaEz
T+fCgFa2/cQ/7CIgQcd36VNmqcQMMjo/Pa+jlfPinn6RiMZ0njTdytrf8dsb
cQ6XLtLNGwFLzQwIF7Yi0dc9G2IEO6IAI0ObLorVpQkp+gmmoQeL7P9Gj0nw
QmB8Wr0qAf84E7RU1FGqdTSac6Ms2UYWIrBGenOl9HP3toS47nbCKfGJK+oT
AFhbw3Nih/t68TguHjXVC406GeSyVdKGwFmgSBtW5zoU0zeCA2QpDQ1pjF3l
PQvxkgTape4JoRYuGTCcqh46hKKFOlketbFw5/6O8YgKe14vi/loXlPs39Th
GLHNH/xpfZMbCnDMMffy91WtDZCxwCQxu/Z2MKCKNIr/fgVwmwxhGQd8KgYu
MZZXDfhM5GyfOB6gErYPsxETNuom7vvpCdWawjX2B3dcaaXF197jwG9PnWR1
QnPRLKf2c2Dl5MsH7oAOyq86E5CrJXIQyksgrsRj5E9u63w5YuLB0qbqKAJT
4w4xIoF2z5SKaYqPVb/fgnJj2zgYcB7Y4k0MJH/nYfqMbpRlaaBmev5Yhl+Q
+GVIax8QTgWVQ8s6QwnvaW0yV245AFl1dfarUnO6YI5rUOhgMvytPKju070h
5I4Rv+IZl/XgWrkqBz7Niw+VZBLjbnWLn3zhXJ6APv0V8M5Z7IeBtT+5NPD1
gu11LPt3wqfYG3BbjRapEoEoVhACb7JqTgNRQsdtM+0krtzdLcN5qYIF+cbe
usFKjlSg9VWfLGrLe9leVoWHcW6LT5Zr0Qamnohu0GzLKpje1r6MQVnboYp5
ucclMyiTlFxxsaj/Q4b59Hl/4ePncLIIvpEQDSh4D3mFJdNSzEf68cIsVrJO
c9nAKsU3g4eiCqje6bsyhY5SxxJufeWVMUvKzYNlGBKpTFMFG5Ok/opFijjo
keQlchs60U+4PwDOz/kp9iRHoIIQXm87w6SQgXXBejy80AtQFHp0A/thz7qk
4un26B0sy9F4ujBCHYTTUgWhKRXkKEkHUZeE63q79c0KU55kDk2Eyhapst+j
763FJ7RclSK3n+NX93A1TKAdwNpNACUk4q/EcUnQQ6UX8utYqepGjoZGzC/+
DP1V0fHEIVxo6x2/HuPr8GYEv6utoaeNPHESC8594z0a0OsfLLLY7pmz9ko8
fY//lLgKxn64/4JSd/IWHd3JqgqD/yC+kyRQOY6upwDx9960NhC1KZD389N9
juqthESzhPmv6adX1/jzPJR8+Y0F3qYaY/t4S4pISZDq/aNiah7fDFw0plX8
j3+1EzqP6wvUoZhi+LSUyq1YKiFMDqKzS+6eFnRbG7rH3Hg5ww5lcq4h9cdP
mnFjaYM/ft9xG7X/8OJEWH05W0WIbrKYSRCltiZtfo8ypp0hBOzdsZTybxO1
Dl41+d0Vsuqb5k0qT0WcDt2WQm/qDwb9Zcf/vEwLG2kLOaCCtvPJ5R1eORqH
T7UHCC2qguwveEDRzdXI0KJRzio0EDUMPHMtFjSshPtmQcrL0sxUSu1R338x
65lfAjbxQz+EV4loNOJ9EEHZoyyUhxXlZ7/6OQj1o3NikMw3/XUgrMgAA82G
hFCU71JD3DqHuEBK1CCi76EqRRWQClFEh1LBcdQkRurTeyuqiNdXwS5j0lHI
AQ4JA1yrpLSYQQ+IEFBobQMdZadtN0e5w77mboE85TEQ0P2ttk0y3cmJl4eF
yzFLag3stnoIiJdJVM1p95dF7N4uiGOprxH7oMpbtA0pzEdoQeoo0Oejczjz
CYhP3vRVLkdp2EbXmujeICRB+JzrYukxZH+OKfWyfWrI5UEItY+nRomFyJde
fJwNoTxlK/CHhiIO9s45GOkoyyHQC40J2EFyuMEV8p06kpVDXwwiwGqlWlER
eZ99G8C8I/ssl+MNdGEs5Wq4icd3l9+3RLDfRFLspzopP50noaFMijuEYU/k
eEQCYDFA5dQLNL6nRwiWvaWqcf6TdmiAEUH9iFLYoVtaAzVxoiCY5guW3SBF
b47Es3+sorierjnIbO5iR3f+9NvwNG/i0PC6FNjRf+82HSGPLbvuEIbyHgmO
94Gd6NdzTwP7Y5+zV5Xk4i48FbGTHpSs8kpU3j3SZ3g+eC/qRwBkL+nx8XDN
qkhHhzUqc3zKaHD1nh91wFJlg41ObamU5EKIppVDK4NbwmdTxVZSDhMAg9z0
yA9VSj0yvJ5clbzsqkAZ7osJwgLpBQy+a4BgvGykyxQU83fzMss6HuM1nTm0
bY8Fpmy9C7BRjgi1Kdc1/Ry6R7BeJchKndF4KiO57pEs85Dp+qLTuctUPyOe
i0WQ2kreST+uXefTCdyHCSI84hmSX9Wq76DhnHj5WrjpvvBTMrAYOGksG4oG
nLTXIUj5T84Kd85fqXqMTTXXEEEu/4RTXhQWlN1WX5u8WDFMKhZiJ0vnJrcs
rw2fcOajVGh1RuNia0HHN6/p4wwr85i6NUgGyi8o1pqMvza7kOIi0VRViiht
erYGbpl8AVJole0/rnBbp89JOWM++hv0qmNFHyfnglU+YQwXto7bNkAX6ajH
r/jtOo20AqBvyHugiJVSUr8dlWrVc2nAfGLe28NZAPJTjlEWVWc6EaWk4BGx
kOdCh1YXb44K+lc5kVTTpfHqZhYm3I+86oyzjX53p5MHYx+wVitVHnMeu5jw
qJmT5V4Iw0XNpNbiJbLOlBZoAzOI0J6NfC2w5tPIINUAYM3Yb3XMtK3RNXJc
J6slD1786yvfLVezmhD+X3lNb6wYaU3SuSXkJDM3Hl3bqZvS/zhnmXBPMYdy
eatBkxiaJa1/BZYns3lVMdCzCsQZG4tAqnoc0ZWasiAEj2QVwdvGG4lKN+oO
KnVgh/pF5leMEHt/y1a4fDIgSeMGk5XiPGCMDTNBQLehCX+Gyps0ntq6uCaq
d3+TeKx9nO6X1oIwCsQiKY9agXmKKelyIAGUSdIBRVf///z6zjD83vmCjul8
HZEPTuf2b8zGUNcsPl2T/rlotBoUUUo8+eQ/CIwfyVe+MuxUjJbGj4Gm5+AW
+yeB9lpSByZrY4H08gecXl2y0DzXgFYR4DeXX7lBSrz2joG35PgZa9Mt7NXe
y7vNQ6dpFerr4darBPdo4PK6cl4ABaqCRycrSvfrO7lMK6CSxZkaSHLzdYBk
MxWTgDEmjhZ6ezTz9uCx4SrPQ6QjhevgOQcgjFzk6wVBpzfkik9L7iZem12i
JqHTi2mGC/j8PwthM+5+HwjMjKjr+sQ0dt8XcrEfOljtW0thgJhRWuO1NyXM
glVzD+DVIXFIFBwCGFnGfLBrLwyvl3jyafJ/krGfL4Qa6mB1VaNsywB1Mrou
kNkoTGKbyUjcIC5Js7uk1p/8kYvPG9BB1cMMN7DKF4u8bBgtqBgHW58o6MOP
piWKAdBVq1aHT/wh++mZ1G9b+EYqt/ROwzOTOXdLe6HcHVirPaZPvXrCGn6/
51ayCvLA1uDfuZeBaPDlPQBL5rMaJ/2A4VOSOwUZZdORiSzG9QlGSrJt0sP0
0MEPWdoQM9hPLUU1zDFMniY+WZlx/nt3jrS8CFWTtSYxptAPm9EQ199mbccY
76UxlqXsDS/rRdMXjeJP5wJ1nIHoM82v1KpVu0AbLjR3gVhNygWaYFFf0Qfm
iXJquefTZA9LfiLSZmaICWKNpsaa43JM74pc7aJlM0xZUh5yqOqj2+pPCu/X
PZ567/b6MQIdPHhlQ6e3awuvnqPXE36lHb7+6Ka9GRX6hwdrzQ+ZTdj5sJIf
81RCOxfBiq4dVxQjbEa1Nz+JEtGZuNFKKsKuQArH3pweajHL1U7GwVNRzjuN
o3wQbzzhEDcZjvRoKM+zXEfYdknRWX0GEUaqB+KJ7yFnwWCLgrlyMDSmpq7L
anQW4U6Ll8Sq9cIP06mpLT/0PE70FV+LO6jlbap3dW0/1xkLjHjowZ86srte
tr6QJUNinI5O8eW9lU9LqKg0IOVN0/jSZaqqe7jbOnBzOL43a8mMDho1zUs1
6EIQhAOsWWXUNkbs3eVmiEaTPjeFzpXiIPTdL3CCaEYPQ9AIXHlXS8BbGmfQ
YSUxkA7pkSgKkQOC7whnGT4dWX89XF50hSQNsKgI3FvyKqCiwR01jQ0uofcB
7HyxLN9ucBTvUgbOmBMldOWIR9ECyWJe8InL32k4ek/srKJXR/nkX88/ivhi
WJjmURUk7PHe7UX/mtruoswcGYc1y+6ICRMrvoxH+f4LbJxeDntRxwYKClGR
H8KDjCE1/oXo/c/nb53Fgf+ukoQkZhHsF4ktkjNANjO76NDw3Ha1yueIm99X
XrZX8Qw/NWNsvFQw0lce9zsNOoliLOhFtsagyE5okqDUEtblTZqkIRIbNmL4
O+GIuyPN5TwXnzKbmJSqzcjHKdIliHXyQa8HA4qiNjZkKOIDuAw+7budUwLw
EPMleuO8d7hgntHdUuCNW/rscfr4SzuuPj8yK4CMlN8kDO7J14i/hZEfABeM
dJascQzA3U66SNL2dlfqXFgZ/z+M/5k/fZOiRSogq358CVGefZPySXqETlkD
5OxLEcft/hZ6mJirt9/MeTR3ZV4Bheks+I0A0P1HsFS0afqdd7b26ixCyqUz
K3+hkDTMEbaQAQaq+lOHdVQ6prX3BT14JZlZbtRsVnpRgnrTLnvxgWJufvjz
3I12MmjQLh1TZen61dRw9Y19zpQy2EOOIjVIUbCKZ4dk6Lv7Bx9SmSlBE/+N
bRqMmCjs/+5pxf7kajEbquiKUKAYNoo0gNuE2ylzAJf/IMRk8hmnHZ1jJYHB
+Aw05qx7RcE9DshJvs2V3D3lI7qaLUG7lFmse4gQWEmHihHoNYJwpEjfSQPN
6Pl/ZESkIqDK43tQAOCqc8IMpW6fl3dILOuwaBloXBl8g8bCr9gic5Jyu1g3
jn3z1OT4ZY/hmMWYzwdUXAF9LbqKaa8jJ9sEZOzGLnxnnxBMLTCWVJY3653i
ixyiTGhDxmFRfoTzruswWU0huQgQYVKgtqZoA4tZOLOlsKYKeUJBC6WHdRSD
7b/iJiNfLGR+6r6IHuyTARDz2d4M+9nY0Bk7qhVqM3L2I9S+wefBm/sttIIA
RaurCxHEepPSWGibXf0WG3GtJJhszr0zAGVniNxrgkUonPlQNB9okXd/rMR/
IpaFtBya3ct0Ae6dmqTiG7Aoh6rF2urJ8RAYs0hJoH9REAhyOBmu8k2q5dgQ
l7NmxrM2wqN1/5pulpQgOQVwMssoTrXkgot7mPVSm/2GAlLPzJ3FGta0OGlj
bOP345qJT3T4hXUzPEfUyTLQAqewbx8wMl6TiFX0LJqwcT25SG4+QnIjJFg7
izNAptn4DZS9+IN35c2xKfVi6q08SqoPFLVcBjghTI9iHSyNqz8kDS00H4uz
uNyAHKHnB0Fq2u4nAvlK3IBtAFjzGdoFFQ+CPoMVaSr7+BOyQIWknTj/f0Vu
bEDmWN7L4wrdoo+vaH/H6eTqBKd0dOTXJpy0a9UsyiA6w4Jy6qmPgw3uf0O/
H656oZ0sTU1+LBHWyKJ5AbfzbEb6UZb6UBVFfpF7WTkdzDfLPLe/4kMosKCQ
v54kh93vxUHIsWYk95pRrHnmc0zfp423yrMwx4AAhqr6C04U2dIYS8nfeXNy
hp1MjY+LDPdAa2kJHrkxqc3HfS6FwUfjXIgFtz0beRfn0rL3jl9sWfPfuF7j
MDxIafJ0ZanOzE2isAhZWpp8Y6TGYkN03a57TQQymiCVQ+qU2dGlLduPlmEk
+y3qfj1+g8lw6XkNGT7W7NQCdRjFsS1CJZeDMQcdP0G7Ri1dqbhDmU2zQwG1
p3XA62DA4WgioN/0U/S+luatLvCx14IsWDcJIKeQHa6VE64YSL5ABQMxEudR
n3QNPAgkN/zMM8Xo7BOeTeusoJf4B8nxAanVthDcPgSO+aPQ56VoXoL5E7Fe
VEndQYjNc9QRTyG6j7YMsAjrgim0mjLuRjIGHpI88ulGPUze9YnLe9ex5eH0
fYMzS5uJn2PHkL3AyBeSYatb52KwA1Z0swzgUUEdhaG+P+tXZsHYjET1vz0E
S1mveMyE4phey+IsaSWydNXl7uy1Wse7ui8hKSrdr5q/XVw2rSs0Yn2wUykL
ZylAQyEeSb1m5jZ3EV06EztzrAOKesVbP2O5NETQzWDlycBTzmBn+8nTpckb
sGeQNig3dgZpVU3dwClsUOvLR7J9YcghfqU3Xvw3gV9+P7poYK/nx+yfw5iT
Ea7dQKE28SwKHDpvQ0qwYE3KeFR6rLt+K0MiYyIIiu9dIhpQQRBZEV3qyshK
yyWPRgbzTimgVxU4ef90FqKud1HtfF+qNju0Wymaiukrfa06qUre6n2/tBkf
Nwqo1iO7IoA3HP2LG1i/ziEGtKj6A32WxghbLSDxW4+b//xoY60l11CijbRy
pHpqdCvdM8qoEm0q7puWSnIjbJI1Nxkhy/JI5r5FmmxqYvgit8dSTq08JtKZ
xYx0ZmhJCW2BDFrzJpYqN6xuHijsuLuXvG/TgdM6YHmHi+gf7SF4uoO3bJUq
nmNLx+a+lYDe8Y8p79zantTbslalplPz6PDR7GtbpCRbm7VWzX2Hm61Skjf2
L8c7Y3tW+hA8YYbIXFaDMjHcGZHgMVeBijIy3DFWhCHqeqen+sZ3BrIDSzw7
9xViYNulS15fxTd6fxu9DMnjNvljg/X0lFVHkZTSBukD0eJVK9lW5TIndzBb
pYxjSYHu+kgQ33WFB3Niabp41Rtn+fjC5AmJBSgbiHx3AYVYBY8DVoX4ULXV
FCcgRZJKqeY6crw2gg1k8WgZidqhNYaKlX+IYQeOqcCojstwNRGEAytscEMU
N3+6yelpgyrSMxE9eFDQSYYcgrhJK6NXvzdF0MvKMEd7hxUbHbY8B7bvPUm1
wCsOGW6ODJe+R/L1X3FS0mgIsHZDgE+6U3C1FJiqzrwxziVIAX3vZ/h+nbZ6
UHihmpI/2AxiSEHvfN24GrLfzScdrjDhlonml9qE8rNMvBo/Rpcnn153ighW
KA58LuAvUm0rHvJFlAXGDo+HsTXguIh3uOkM3+Dp1am9bGLTHkDMDUfZMZdv
QjLWir9/YwzdESJIFgH0phePwPuOQR2hPAlBW30kaAxmMKM8hIrUYIxX2V/Z
XyuJuLglRd8cx4Mi2UuraLnKe32d+PXRRQBQr2I5rxqhFfuJMYm6FPj9K/pH
3ONubKIn7T+2O+fjdAmfWvjoeEA7PCx8oM83ZoWflhjY6Xk+KIc+7/BNwkmj
dK2STcJoBnv9d4s47E+ceJ++rgkHVtisU8ZiXudyawE2fAlff6Ltuw3udcHo
5+uXdAfZ/7DNHmD4BB4JIYSigYkCYqX9cu2t8vPpHqEksQdOPdoiQ2jjT9qG
voAnDHUwGI8ja84uPXTzk21F8ZVL6SnAs+sr9Z3MCEJAEpnxWGGfu6TNHRzM
Y6cOen2dOPUqFZo2P2WWJW9quJdHXqX8SCUV8Zhaz2AeH0Lg3TAjZVwIhC0X
Mdl6y6Wdu0363eEODwutYO4nSaCWUwmoadrI/QM/KusyyZ7c8VDBd44b9LKA
H3sL7OgFdrDMPWz/2CQ6se87UaRrHX8zN4W/zIMRR1DA8qMB0BTSTS0A7B9U
Q1EJ6cgFe1bNvhMsE12D4ht+YuKTWUtFYIleCZgmO1RNWPdxq8chnHGzYS15
buRulM1Nf+0WD9qTME7r3C9DYJuO7NtQsqY9m0H4rH1vEGVsXK+8lGZ/ugEj
9VoNmV3MgzgIbQrhJ4vg09NQdyRqdmLHtVAs71RDYu3Howszs85rqtADEN8Q
VNFOJpiKcTNIDicVr68YqD5zk7EziEAiLMuzfXRWIS39gVQYLDJQ+vMbj89R
pP5ffgOXDHsgxqrZPv9fVEA/mrHUrFOusp1tTIXp6gHZWPKWy2yDI+WQ7Wim
i/nTup5D6gvD7ukqcPnbm7R8ZMT4CQe28b21Zc1s47j5gYCY+7P60KOGBELP
X9mibrq5xtqYS0eTvIJ9Frgnj5TL/DHFHmrbyRrx8HGIumxMcfBzR1jxsscw
l5aekJCskaf8bjYWwxMfOAnpM5UoGg/9SrnsKPJ09qf2WYXTP1NDIc1e/UxA
7BJ1HQrAkOsUupiUyoUxAuuQgmPgQe/TcoAtzNejWNXQLPkt4ciG5UyPT3SE
iK7Sx1JbAloj3mckrf3BDD/qfp4Usf6+16O9YeQbqYGkq+N/BOSFc660RsKo
89tgd6evyjU/DEjbSHdXHyUK9SJ6XyeBMmVPEJ0VX8EhLmf7Ee7HJbVQAfjA
+iCTtwcyevdAa/Upn8jShlSAqAMtbISXsp0Xhb4aJETgb052YEU6u9r2Ju2l
7+w85m39X2z7d1YE40Z9OE0v8n8NO/G9X7pYMcIjSsJI8A640pROYU7qzJax
la8d4s4L8ey44fS56CotNtC7wIkvW7raQ7o1yK0HBWX1wZePFFUxWfabUh8Z
dCHxEqhbhiRihgGcUsY0zBtd3OzOLcWMTHaQW2/JaE8Ap5OS0Z7E3TNaVoQ7
y6XbRfrIZYEY11ke3KjZUVjhNE1GTy/Q+yXuIIWBeqU47hDqztVOTwYy6lv7
p3pfIYurYmi3ySCpY8yVWkoEpUfLvpMIlynFoNvat6qyf9Cm3Y5QqVZ51gcG
zDrnMVeQIZp6cF8H6tMOuBj25XHM2vX9h3eekk4zQyhJ5CbhbIwG3JsnQyFC
qlaTTaaq1SROFqVerfLBvAz/4HzDNdiAF0JeWt5fH1GLGS6uKRCPY8kflkFo
Oc4nPMiZcx5CypV9AJEF/Pn0gDGY4bfEnLE6RWib9VesBd00U9HsO72HSgPT
qSCepYxRkt0FP4EpwNJgW9R0k2u450s00RAcEx5IDyMyqmM+2fEebie703bk
rR8iAjojly6fW9VOhFwJZglVKHVyT69qOLDpyFaOm9yKeAYA7dfCrlEOUMbg
HFRNlNEa7L69DG5TRse1DrUrHepQY87D9jvXf9aTQdVeyeGGcElh/5VcMeI7
SZ4xFfqePlS4XiApPOdSr2cDcdrUY3jfxaKB6hwfeWzzp6KTXiDBUSHFhHbw
FoEhG3xu7qp9NcFTKoJc1BexASiqJHyt1IVAogUK2VmDBpFsVuFlX9F64stg
m3mkw4fZmwrkhGb3ASQf7+kfyP2fMhgYA3ckIlxwt6zL9NXVav4epNxzqd2r
zPHft33k1/MIV+tdakmXn8MT0cUiQu5PNiMy3n9hay1Y9vj2i2kzlIrr51IM
F8qFZETXJcyvr7tQO1yOc8dj7nPlhE1PlwSu8NclH3aPzWdWpD1fxSHmQCVB
WSZQtE/thimJNleubA9Rbq/zlZiCd/0MhlJrehA273TLOgny83EZ/EWtqJ4r
VjFq+d5Shs9g3FEvTuxFcQYYGfoaCKw108R89fPrg496snOCpnrosuVykxOA
BrouxnA+HzwYxCcX90sitkMP2nqFCYefrCXDY2PeJCET2sgQhJxgDfYro80Z
OcpdBOpp/xK03AcjE99fBefzjRBuGa+hBhgaXI0ivlWXULhxchvfUATflw+M
a+3/77CDXn4/3LVZUvJeHgUq7GiQ6jV0lpJniuRJ0hfIpLp5qZCafr7ZRkCE
lDijWj0lcRZLG0FKd2y/tS2Iy9kAFxgHD1Eg9SSap4BDzIjESfwdvRBtuPbY
h+0zaSmka0uNQfv2BQ/HG5mdXiRClDn9XhcvP1AaSSeol06Z4S0hcX3LOzCc
/ie0WqKFniCiM6opdnBbPzinekMa1T3oc9VL6shiWEek20C3sZo1RbYhCLY1
5mbjxeCdB5TwnpiCjml7LkTi3P+7drbwiNLcz/9lzD6jIBRbCVeWruDV5hnD
VbLuO0gWWkgogYHtUOi5Qh389DjBFczMFzBzqWwlBBb7+lxs5YuJGTPAHvQ7
r0sLSgGxS7PIDSqjgeuAN7DWZ6ss0FEjzjSWDXVk/giWkJdwIv8Hf/leOtqs
41SNyI8Bpfl//q64k8EYphWyMO+Deh2yBMqXwgLlvzIEccvSWXdHJ188aygo
rG3s83DqTlUNZUPqN6Tiq1z5yQXeyQJeKGq8njom+HRvp3ot2gnluxpP8xzJ
oo9Id/YkqalvXADirMmtjEgikOJh+dRhK6rfQ7qocK4SERUgaNTjIP+VrmLE
z/hhja6wKy+dtJ5ozV8xjOEG+jR2PuIEKwkHSYm6KVaGbmo70iytsU4zaiKZ
KRINPxl8NWnxZybt1bFdBOCQ5pv7zkm9YDAVMig3WodlUKmOyQs0T5sqlLY7
7zAn1TEIriV1+IHcSB3M7GpmmEoayWVmq28ZsUO9YVuZqUS3Zces6v1FQmGx
uUyuY2FSIHAUknq7dleA+vrOJ0hw5f/tDPs+lAJBj5yVD3oBr6wkBCoGQyLP
BvL63kBkiri1yCwIfQKm1QhcrvF/dupb397Bq7vj7JS/w5OgVPk3VVDxQ0MW
98+WWZ22q5ncEquf0dJ+6LETHGCySX6q2/f7jpP6iDhgsHvnvXdIB+4Gr3ge
i2aciGUD4/a/pehNyPRAvgP3pRebRFp8Agiv6Ee50Uq6TJho8PMOD5AO+YoO
4ln+7KP70SoE2NkXLoysrtuxXxoBaHUkFqLmk8yqd20kUEvti1RWsPRApCpU
ihH4gfQQ8cW1P4jSw6g4poeqxPeUeStn5KjGPeFKH9UU8DNjHmCcWo8OS0i9
lFNFfELzFYjw7AJe0u4dwF/dQFQLZOfsrf23+Si5OhTZqUij+w6/3TMj4qaO
fTMS4D5Q7Tzv4Wie4AR8viAbvK21SmBX64Q9hu/+l/JOdXcRJowNsksiufJ3
tPnAAJj6Ag51nYeMwiZg9maOjwO6XksEk8uDYL/Sppn+EHYbKPr4THavlb7P
hFY0Qfqkb8mFZjtbsLitmzYIcuRAueqduImtvTBZQFGuKkerUkNXuR/frc0Q
jFFrJsXxnjAVeX1F46M7vWa+vvW+zuCIXddoPP6bAy+0LpnLHNaUunDG2/uW
KLjrQwg5jN7grefKhBcBLG3ETiDnis8+n92xdjf7UIFo8a+4U8n0j8wHUKXc
CUfZ2lzJL20g/eMSPDbt7sQwmX3FnvlJUzZLJD7WT7tpA4hTHNwPeOCBN77D
Ho3JisSe8u5sz7fGU7Z86AQaokJtEb4E15xzye5mvbkZN4YByvEXhFo5Ubpc
QvB8dzJG/t2W4L/fN3h4r6/VdvTBK40G0o7E62TwXM/Koc3d7Z0UqB4T5nAO
vXTCtdDkg1sqc/5e+yNpeDx9q0sA0nC8FAmEExYt6ToDUl/QUDoN4r/7eKHF
opiGvoJ1uRIBjgvAwHiCI6Sia4RTiupk/egXKkEW01hTiO0HEeIo0Sx9Zvqh
8xLUgE+FYZCpDYaXjctuH6TAPJwzJhJ2CALCl7BGXCQlcFlwqN8K3y+38v4x
JN/4vaHtm/XUo2BPUsHHjkiY+oKqdTi2Bj36K8FfOuUz//3VHXeBxz5SQHjM
b97ltSh08U57p10RuPIhsHA/S7aJ994AqDPB/HRtrdjs8xuTpc03aSI1IUaI
27ILYGlv9I/7oN/ApgYyfuN5Pn1xzeHreUn5+ZDSa04YlYawSQ2iaTeCP0EU
wyVKiVs9ooEtkagFFoysAZ8O9bdm/8DU669MvA5GCyYKwgPxazubCczzu+M0
m8DM5+kmqpPLLslchIj5t2Ik/3nTXrpGn5CXc2yTuVLcNR8RQmWxc6Lwxvx8
/hZB9lMr9+ZRI4CSfs2sB5P0D+mcTKIL8kpaUQqa8KoFM3sNYdmc53MxBm9x
k4iNWziRo+bQoErF2bn47uz0dRy8kSJHMXLziyJ+pwEj9NlWxqLLo4uXhM5K
n4t05917AoV3ZNeoE7TYVd8BRB7lEEcnEqkPm3vxNbzqlh4LN7eSWiUOJQHl
dWEMpQL8IQl+QsHxPNIjNgvCpFl+ZT0p8qhr20BbpFvYrJtxOl+eQVti+kpB
jZYYaKQbPxNHaJtwyGeDaGrNx+0auHRyTyO6DsaV3oWZeh1Az8LAAH4MzD8q
n4V2qEAxVLxjjWEVaXBMWHsxpDgthkKqxy+Fa1cii0mpcUM7l6hF6fJ0/t9W
wwJIj64hNbomjwz1ayg1lXSv0MMVEjgr9dLafbKoHzyL7TjjarJd0btcUkXi
pw35EXenaslEVFpJya5n7KPfSSghoe59xKRzW3TYkWFwfmAvgCdFw9/CjawQ
1VRDpw3wxezLPHxqmNMs8cvhKcwXdinn39Ter3utqJJYfKpORLWW1mxpX1qQ
um7FWDcBPchXhXhALv1wWXUXcyHcR7UfF7fUaPDflL9u8K+Q12BeaVYAcJZq
FQmlWGVxDw4ALexGxAiB0QwP3iQgJy6y/ox/Q4EA0CQDxObN3Nh27tNAHYO5
6Bj0bbzXHIqFb/ILJORe67YNIigShM5lkTelGHwHCl6oEkBV2QyRvghgZoOB
7JTHQDlk/frLqSCykaHHKUtR3XTK+Y6pdrsdwyoU4aoc+Oxhn3VAnjbxHDDM
gKmK+WKdvRVeBbEAyP4ZpSC3jUQr8h377OfKbZSpsk3kVcXMKP8pJbxREQe3
BMeVmy0EMV/JCbKy3e1LjJw4b+y2el5AckZPjy7KPl+Z8i0uUm8TpR15fR8I
BM81jlxowf3IjpF4+/O8NSR36q54jh15lV8FB5S8FnF8mp+KhM9dBbtCHnPy
o1L5+HVLWHNUhITlpJeYg78q1Yza9zuYlYBxKjao2HmxusqpBbFEjiuD6pCB
9MDlxgYtqWSEOTyxA8M0gXWveEZ3qMz/SClFF0WZwMyu6l69v8EoeX+HnwHV
VOPw4+vJjaM4m4IJ2ZLNH6Y+e44xbdzTVOezGDtgkiEvcrMeQdrBKAm8oa3A
orBrTQo5mr3bbV/5zFpZxmB2UUNCkH3uMCNSk8BndYxNGJsSD1uAxwGm5FbK
ogyzLzEf2bVFITpNKIYfLwjgwXE9904KkJ9w

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "AHFS8uhOzEEv0qANUjCa5shxFe8bemKFNhQTqRGtC4pjovR6jkEwCgEM+HVx2+RETJ81jdGctIsI8rtsCu4TOBbfINYgMfPtAhYoq0pIwXzpBYW/Jwh89yYqmQ/8qwf+UZ/RCUPZ9uTW2DZjLM/8DQwcPSaWPn4uluTziVOYaXqZBjqnFFKudtGOgi9fUYcdgmgi1Cr8qg3AFyDXZaw0JPfMHv+sI1tXM9FJgZxRxGML5AbLTGN/IFFTwiD7jWhtuRDpFuy+jVAMmzHxmf4Z1zAH9roueo0Q70esLvAB+Ipw8MMzvlZmvi+UyDijAU2F/28fwyF8nilQUheqcKn0pLmvzpqBrI7XpiY1ykOLphCu8nATULoNeaIX4RHNkTD4syxkEA4vSVr8CJ4hlpZSFGYyzT0PF51dkuqBuQx87j3/8ynMGn7yTBvR7eEAV5eyUpFG6IcSEHZspMmuhTB9Iwo91nza8pUZzK1xJ4eDLQz/ByeAJ9FU6LniJBQqXADlEHosxL6Mn49ysGQIK46vFtRlqPKJa0GmrkpbnU2SUa1+zld1chsIQVM8WfrpBI/bzquZB06xDbGPLlL94V4mvCvG2icQGeh72COWR6K7iNs4KLWPdaCWWP2a4k5ukbVr7PwCpXuOQ1P1OrjLqHaXcOG8HkydlSgAbIbnnrkOvP2sHJG4QOf/ORiRm6/d7pdY6yEOAKt8TVYZeqBqeRb8CoO8ZEW81J/l5fhSSgLk9nUXvErPBdfVrCd19/OfC/sfbImoauwLoE0c8LmoQV2tN9NfQsdGYS8Frk8z87Emqww7p0UG18D8AEf1KlGd6IuSzTIYkfCXb8cTTKr3dVFrND+bkc72tj+JHyhmKQgU09onVhfKpaNx+T3XCrDFzeXwTamT7RAJS0TDN/6rV7It5ntgElaD9r7CKnZ7Ek5QuDHlLad/kILK1MzhWJnxrcHDqIZc/RQ6V2p5u8FWuExjrsEFm+aGiy9nGPGHTvlb4SAsQ7p13coaEO6f3h5AKkq4"
`endif